// Name: Black Parrot Front-end (FE) Only
//
// Description: Front-end of a 64-bit RISC-V Core with Cache Coherence Directory.
//
// Top Module: bp_fe_top
//
// GitHub: https://github.com/black-parrot/pre-alpha-release
//    commit: ceb22c57f269726a5fd99b722521cf7df9d3907c
//

module instr_scan_eaddr_width_p64_instr_width_p32
(
  instr_i,
  scan_o
);

  input [31:0] instr_i;
  output [68:0] scan_o;
  wire [68:0] scan_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,
  N23,N24,N25,N26,N27,N28,N29,N30;
  assign scan_o[66] = 1'b0;
  assign scan_o[67] = 1'b0;
  assign N7 = instr_i[0] & instr_i[1];
  assign scan_o[68] = ~N7;
  assign N9 = ~instr_i[6];
  assign N10 = ~instr_i[5];
  assign N11 = ~instr_i[3];
  assign N12 = ~instr_i[2];
  assign N13 = ~instr_i[1];
  assign N14 = ~instr_i[0];
  assign N15 = N10 | N9;
  assign N16 = instr_i[4] | N15;
  assign N17 = N11 | N16;
  assign N18 = N12 | N17;
  assign N19 = N13 | N18;
  assign N20 = N14 | N19;
  assign N21 = ~N20;
  assign N22 = instr_i[3] | N16;
  assign N23 = N12 | N22;
  assign N24 = N13 | N23;
  assign N25 = N14 | N24;
  assign N26 = ~N25;
  assign N27 = instr_i[2] | N22;
  assign N28 = N13 | N27;
  assign N29 = N14 | N28;
  assign N30 = ~N29;
  assign scan_o[65:64] = (N0)? { 1'b0, 1'b0 } : 
                         (N1)? { 1'b0, 1'b1 } : 
                         (N4)? { 1'b1, N20 } : 1'b0;
  assign N0 = N30;
  assign N1 = N26;
  assign scan_o[63:0] = (N0)? { instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[7:7], instr_i[30:25], instr_i[11:8], 1'b0 } : 
                        (N1)? { instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:20] } : 
                        (N2)? { instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[19:12], instr_i[20:20], instr_i[30:21], 1'b0 } : 
                        (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2 = N21;
  assign N3 = N26 | N30;
  assign N4 = ~N3;
  assign N5 = N21 | N3;
  assign N6 = ~N5;

endmodule



module bp_fe_bht_bht_indx_width_p5
(
  clk_i,
  en_i,
  reset_i,
  idx_r_i,
  idx_w_i,
  r_v_i,
  w_v_i,
  correct_i,
  predict_o
);

  input [4:0] idx_r_i;
  input [4:0] idx_w_i;
  input clk_i;
  input en_i;
  input reset_i;
  input r_v_i;
  input w_v_i;
  input correct_i;
  output predict_o;
  wire predict_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,
  N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,
  N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,
  N404,N405,N406,N407,N408,N409,N410,N411,N412,N413;
  reg [63:0] mem;
  assign predict_o = (N52)? mem[1] : 
                     (N54)? mem[3] : 
                     (N56)? mem[5] : 
                     (N58)? mem[7] : 
                     (N60)? mem[9] : 
                     (N62)? mem[11] : 
                     (N64)? mem[13] : 
                     (N66)? mem[15] : 
                     (N68)? mem[17] : 
                     (N70)? mem[19] : 
                     (N72)? mem[21] : 
                     (N74)? mem[23] : 
                     (N76)? mem[25] : 
                     (N78)? mem[27] : 
                     (N80)? mem[29] : 
                     (N82)? mem[31] : 
                     (N53)? mem[33] : 
                     (N55)? mem[35] : 
                     (N57)? mem[37] : 
                     (N59)? mem[39] : 
                     (N61)? mem[41] : 
                     (N63)? mem[43] : 
                     (N65)? mem[45] : 
                     (N67)? mem[47] : 
                     (N69)? mem[49] : 
                     (N71)? mem[51] : 
                     (N73)? mem[53] : 
                     (N75)? mem[55] : 
                     (N77)? mem[57] : 
                     (N79)? mem[59] : 
                     (N81)? mem[61] : 
                     (N83)? mem[63] : 1'b0;
  assign N87 = (N147)? mem[1] : 
               (N148)? mem[3] : 
               (N149)? mem[5] : 
               (N150)? mem[7] : 
               (N151)? mem[9] : 
               (N152)? mem[11] : 
               (N153)? mem[13] : 
               (N154)? mem[15] : 
               (N155)? mem[17] : 
               (N156)? mem[19] : 
               (N157)? mem[21] : 
               (N158)? mem[23] : 
               (N159)? mem[25] : 
               (N160)? mem[27] : 
               (N161)? mem[29] : 
               (N162)? mem[31] : 
               (N123)? mem[33] : 
               (N125)? mem[35] : 
               (N127)? mem[37] : 
               (N129)? mem[39] : 
               (N131)? mem[41] : 
               (N133)? mem[43] : 
               (N135)? mem[45] : 
               (N137)? mem[47] : 
               (N272)? mem[49] : 
               (N274)? mem[51] : 
               (N276)? mem[53] : 
               (N278)? mem[55] : 
               (N280)? mem[57] : 
               (N282)? mem[59] : 
               (N284)? mem[61] : 
               (N286)? mem[63] : 1'b0;
  assign N88 = (N147)? mem[0] : 
               (N148)? mem[2] : 
               (N149)? mem[4] : 
               (N150)? mem[6] : 
               (N151)? mem[8] : 
               (N152)? mem[10] : 
               (N153)? mem[12] : 
               (N154)? mem[14] : 
               (N155)? mem[16] : 
               (N156)? mem[18] : 
               (N157)? mem[20] : 
               (N158)? mem[22] : 
               (N159)? mem[24] : 
               (N160)? mem[26] : 
               (N161)? mem[28] : 
               (N162)? mem[30] : 
               (N123)? mem[32] : 
               (N125)? mem[34] : 
               (N127)? mem[36] : 
               (N129)? mem[38] : 
               (N131)? mem[40] : 
               (N133)? mem[42] : 
               (N135)? mem[44] : 
               (N137)? mem[46] : 
               (N272)? mem[48] : 
               (N274)? mem[50] : 
               (N276)? mem[52] : 
               (N278)? mem[54] : 
               (N280)? mem[56] : 
               (N282)? mem[58] : 
               (N284)? mem[60] : 
               (N286)? mem[62] : 1'b0;
  assign N92 = N89 & N90;
  assign N93 = N92 & N91;
  assign N94 = correct_i | N87;
  assign N95 = N94 | N91;
  assign N97 = correct_i | N90;
  assign N98 = N97 | N88;
  assign N100 = N97 | N91;
  assign N102 = N89 | N87;
  assign N103 = N102 | N88;
  assign N105 = N102 | N91;
  assign N107 = N89 | N90;
  assign N108 = N107 | N88;
  assign N110 = correct_i & N87;
  assign N111 = N110 & N88;
  assign N146 = (N122)? mem[1] : 
                (N124)? mem[3] : 
                (N126)? mem[5] : 
                (N128)? mem[7] : 
                (N130)? mem[9] : 
                (N132)? mem[11] : 
                (N134)? mem[13] : 
                (N136)? mem[15] : 
                (N138)? mem[17] : 
                (N139)? mem[19] : 
                (N140)? mem[21] : 
                (N141)? mem[23] : 
                (N142)? mem[25] : 
                (N143)? mem[27] : 
                (N144)? mem[29] : 
                (N145)? mem[31] : 
                (N123)? mem[33] : 
                (N125)? mem[35] : 
                (N127)? mem[37] : 
                (N129)? mem[39] : 
                (N131)? mem[41] : 
                (N133)? mem[43] : 
                (N135)? mem[45] : 
                (N137)? mem[47] : 
                (N272)? mem[49] : 
                (N274)? mem[51] : 
                (N276)? mem[53] : 
                (N278)? mem[55] : 
                (N280)? mem[57] : 
                (N282)? mem[59] : 
                (N284)? mem[61] : 
                (N286)? mem[63] : 1'b0;
  assign N163 = (N147)? mem[0] : 
                (N148)? mem[2] : 
                (N149)? mem[4] : 
                (N150)? mem[6] : 
                (N151)? mem[8] : 
                (N152)? mem[10] : 
                (N153)? mem[12] : 
                (N154)? mem[14] : 
                (N155)? mem[16] : 
                (N156)? mem[18] : 
                (N157)? mem[20] : 
                (N158)? mem[22] : 
                (N159)? mem[24] : 
                (N160)? mem[26] : 
                (N161)? mem[28] : 
                (N162)? mem[30] : 
                (N123)? mem[32] : 
                (N125)? mem[34] : 
                (N127)? mem[36] : 
                (N129)? mem[38] : 
                (N131)? mem[40] : 
                (N133)? mem[42] : 
                (N135)? mem[44] : 
                (N137)? mem[46] : 
                (N272)? mem[48] : 
                (N274)? mem[50] : 
                (N276)? mem[52] : 
                (N278)? mem[54] : 
                (N280)? mem[56] : 
                (N282)? mem[58] : 
                (N284)? mem[60] : 
                (N286)? mem[62] : 1'b0;
  assign N205 = (N197)? mem[1] : 
                (N198)? mem[3] : 
                (N199)? mem[5] : 
                (N200)? mem[7] : 
                (N201)? mem[9] : 
                (N202)? mem[11] : 
                (N203)? mem[13] : 
                (N204)? mem[15] : 
                (N155)? mem[17] : 
                (N156)? mem[19] : 
                (N157)? mem[21] : 
                (N158)? mem[23] : 
                (N159)? mem[25] : 
                (N160)? mem[27] : 
                (N161)? mem[29] : 
                (N162)? mem[31] : 
                (N256)? mem[33] : 
                (N258)? mem[35] : 
                (N260)? mem[37] : 
                (N262)? mem[39] : 
                (N264)? mem[41] : 
                (N266)? mem[43] : 
                (N268)? mem[45] : 
                (N270)? mem[47] : 
                (N272)? mem[49] : 
                (N274)? mem[51] : 
                (N276)? mem[53] : 
                (N278)? mem[55] : 
                (N280)? mem[57] : 
                (N282)? mem[59] : 
                (N284)? mem[61] : 
                (N286)? mem[63] : 1'b0;
  assign N214 = (N206)? mem[0] : 
                (N207)? mem[2] : 
                (N208)? mem[4] : 
                (N209)? mem[6] : 
                (N210)? mem[8] : 
                (N211)? mem[10] : 
                (N212)? mem[12] : 
                (N213)? mem[14] : 
                (N138)? mem[16] : 
                (N139)? mem[18] : 
                (N140)? mem[20] : 
                (N141)? mem[22] : 
                (N142)? mem[24] : 
                (N143)? mem[26] : 
                (N144)? mem[28] : 
                (N145)? mem[30] : 
                (N256)? mem[32] : 
                (N258)? mem[34] : 
                (N260)? mem[36] : 
                (N262)? mem[38] : 
                (N264)? mem[40] : 
                (N266)? mem[42] : 
                (N268)? mem[44] : 
                (N270)? mem[46] : 
                (N272)? mem[48] : 
                (N274)? mem[50] : 
                (N276)? mem[52] : 
                (N278)? mem[54] : 
                (N280)? mem[56] : 
                (N282)? mem[58] : 
                (N284)? mem[60] : 
                (N286)? mem[62] : 1'b0;
  assign N216 = (N206)? mem[1] : 
                (N207)? mem[3] : 
                (N208)? mem[5] : 
                (N209)? mem[7] : 
                (N210)? mem[9] : 
                (N211)? mem[11] : 
                (N212)? mem[13] : 
                (N213)? mem[15] : 
                (N138)? mem[17] : 
                (N139)? mem[19] : 
                (N140)? mem[21] : 
                (N141)? mem[23] : 
                (N142)? mem[25] : 
                (N143)? mem[27] : 
                (N144)? mem[29] : 
                (N145)? mem[31] : 
                (N256)? mem[33] : 
                (N258)? mem[35] : 
                (N260)? mem[37] : 
                (N262)? mem[39] : 
                (N264)? mem[41] : 
                (N266)? mem[43] : 
                (N268)? mem[45] : 
                (N270)? mem[47] : 
                (N272)? mem[49] : 
                (N274)? mem[51] : 
                (N276)? mem[53] : 
                (N278)? mem[55] : 
                (N280)? mem[57] : 
                (N282)? mem[59] : 
                (N284)? mem[61] : 
                (N286)? mem[63] : 1'b0;
  assign N217 = (N206)? mem[0] : 
                (N207)? mem[2] : 
                (N208)? mem[4] : 
                (N209)? mem[6] : 
                (N210)? mem[8] : 
                (N211)? mem[10] : 
                (N212)? mem[12] : 
                (N213)? mem[14] : 
                (N138)? mem[16] : 
                (N139)? mem[18] : 
                (N140)? mem[20] : 
                (N141)? mem[22] : 
                (N142)? mem[24] : 
                (N143)? mem[26] : 
                (N144)? mem[28] : 
                (N145)? mem[30] : 
                (N256)? mem[32] : 
                (N258)? mem[34] : 
                (N260)? mem[36] : 
                (N262)? mem[38] : 
                (N264)? mem[40] : 
                (N266)? mem[42] : 
                (N268)? mem[44] : 
                (N270)? mem[46] : 
                (N272)? mem[48] : 
                (N274)? mem[50] : 
                (N276)? mem[52] : 
                (N278)? mem[54] : 
                (N280)? mem[56] : 
                (N282)? mem[58] : 
                (N284)? mem[60] : 
                (N286)? mem[62] : 1'b0;
  assign N219 = (N206)? mem[1] : 
                (N207)? mem[3] : 
                (N208)? mem[5] : 
                (N209)? mem[7] : 
                (N210)? mem[9] : 
                (N211)? mem[11] : 
                (N212)? mem[13] : 
                (N213)? mem[15] : 
                (N138)? mem[17] : 
                (N139)? mem[19] : 
                (N140)? mem[21] : 
                (N141)? mem[23] : 
                (N142)? mem[25] : 
                (N143)? mem[27] : 
                (N144)? mem[29] : 
                (N145)? mem[31] : 
                (N256)? mem[33] : 
                (N258)? mem[35] : 
                (N260)? mem[37] : 
                (N262)? mem[39] : 
                (N264)? mem[41] : 
                (N266)? mem[43] : 
                (N268)? mem[45] : 
                (N270)? mem[47] : 
                (N272)? mem[49] : 
                (N274)? mem[51] : 
                (N276)? mem[53] : 
                (N278)? mem[55] : 
                (N280)? mem[57] : 
                (N282)? mem[59] : 
                (N284)? mem[61] : 
                (N286)? mem[63] : 1'b0;
  assign N220 = (N206)? mem[0] : 
                (N207)? mem[2] : 
                (N208)? mem[4] : 
                (N209)? mem[6] : 
                (N210)? mem[8] : 
                (N211)? mem[10] : 
                (N212)? mem[12] : 
                (N213)? mem[14] : 
                (N138)? mem[16] : 
                (N139)? mem[18] : 
                (N140)? mem[20] : 
                (N141)? mem[22] : 
                (N142)? mem[24] : 
                (N143)? mem[26] : 
                (N144)? mem[28] : 
                (N145)? mem[30] : 
                (N256)? mem[32] : 
                (N258)? mem[34] : 
                (N260)? mem[36] : 
                (N262)? mem[38] : 
                (N264)? mem[40] : 
                (N266)? mem[42] : 
                (N268)? mem[44] : 
                (N270)? mem[46] : 
                (N272)? mem[48] : 
                (N274)? mem[50] : 
                (N276)? mem[52] : 
                (N278)? mem[54] : 
                (N280)? mem[56] : 
                (N282)? mem[58] : 
                (N284)? mem[60] : 
                (N286)? mem[62] : 1'b0;
  assign N222 = (N255)? mem[1] : 
                (N257)? mem[3] : 
                (N259)? mem[5] : 
                (N261)? mem[7] : 
                (N263)? mem[9] : 
                (N265)? mem[11] : 
                (N267)? mem[13] : 
                (N269)? mem[15] : 
                (N271)? mem[17] : 
                (N273)? mem[19] : 
                (N275)? mem[21] : 
                (N277)? mem[23] : 
                (N279)? mem[25] : 
                (N281)? mem[27] : 
                (N283)? mem[29] : 
                (N285)? mem[31] : 
                (N256)? mem[33] : 
                (N258)? mem[35] : 
                (N260)? mem[37] : 
                (N262)? mem[39] : 
                (N264)? mem[41] : 
                (N266)? mem[43] : 
                (N268)? mem[45] : 
                (N270)? mem[47] : 
                (N272)? mem[49] : 
                (N274)? mem[51] : 
                (N276)? mem[53] : 
                (N278)? mem[55] : 
                (N280)? mem[57] : 
                (N282)? mem[59] : 
                (N284)? mem[61] : 
                (N286)? mem[63] : 1'b0;
  assign N223 = (N255)? mem[0] : 
                (N257)? mem[2] : 
                (N259)? mem[4] : 
                (N261)? mem[6] : 
                (N263)? mem[8] : 
                (N265)? mem[10] : 
                (N267)? mem[12] : 
                (N269)? mem[14] : 
                (N271)? mem[16] : 
                (N273)? mem[18] : 
                (N275)? mem[20] : 
                (N277)? mem[22] : 
                (N279)? mem[24] : 
                (N281)? mem[26] : 
                (N283)? mem[28] : 
                (N285)? mem[30] : 
                (N256)? mem[32] : 
                (N258)? mem[34] : 
                (N260)? mem[36] : 
                (N262)? mem[38] : 
                (N264)? mem[40] : 
                (N266)? mem[42] : 
                (N268)? mem[44] : 
                (N270)? mem[46] : 
                (N272)? mem[48] : 
                (N274)? mem[50] : 
                (N276)? mem[52] : 
                (N278)? mem[54] : 
                (N280)? mem[56] : 
                (N282)? mem[58] : 
                (N284)? mem[60] : 
                (N286)? mem[62] : 1'b0;
  assign N287 = (N255)? mem[1] : 
                (N257)? mem[3] : 
                (N259)? mem[5] : 
                (N261)? mem[7] : 
                (N263)? mem[9] : 
                (N265)? mem[11] : 
                (N267)? mem[13] : 
                (N269)? mem[15] : 
                (N271)? mem[17] : 
                (N273)? mem[19] : 
                (N275)? mem[21] : 
                (N277)? mem[23] : 
                (N279)? mem[25] : 
                (N281)? mem[27] : 
                (N283)? mem[29] : 
                (N285)? mem[31] : 
                (N256)? mem[33] : 
                (N258)? mem[35] : 
                (N260)? mem[37] : 
                (N262)? mem[39] : 
                (N264)? mem[41] : 
                (N266)? mem[43] : 
                (N268)? mem[45] : 
                (N270)? mem[47] : 
                (N272)? mem[49] : 
                (N274)? mem[51] : 
                (N276)? mem[53] : 
                (N278)? mem[55] : 
                (N280)? mem[57] : 
                (N282)? mem[59] : 
                (N284)? mem[61] : 
                (N286)? mem[63] : 1'b0;
  assign N288 = (N255)? mem[0] : 
                (N257)? mem[2] : 
                (N259)? mem[4] : 
                (N261)? mem[6] : 
                (N263)? mem[8] : 
                (N265)? mem[10] : 
                (N267)? mem[12] : 
                (N269)? mem[14] : 
                (N271)? mem[16] : 
                (N273)? mem[18] : 
                (N275)? mem[20] : 
                (N277)? mem[22] : 
                (N279)? mem[24] : 
                (N281)? mem[26] : 
                (N283)? mem[28] : 
                (N285)? mem[30] : 
                (N256)? mem[32] : 
                (N258)? mem[34] : 
                (N260)? mem[36] : 
                (N262)? mem[38] : 
                (N264)? mem[40] : 
                (N266)? mem[42] : 
                (N268)? mem[44] : 
                (N270)? mem[46] : 
                (N272)? mem[48] : 
                (N274)? mem[50] : 
                (N276)? mem[52] : 
                (N278)? mem[54] : 
                (N280)? mem[56] : 
                (N282)? mem[58] : 
                (N284)? mem[60] : 
                (N286)? mem[62] : 1'b0;
  assign N290 = (N255)? mem[1] : 
                (N257)? mem[3] : 
                (N259)? mem[5] : 
                (N261)? mem[7] : 
                (N263)? mem[9] : 
                (N265)? mem[11] : 
                (N267)? mem[13] : 
                (N269)? mem[15] : 
                (N271)? mem[17] : 
                (N273)? mem[19] : 
                (N275)? mem[21] : 
                (N277)? mem[23] : 
                (N279)? mem[25] : 
                (N281)? mem[27] : 
                (N283)? mem[29] : 
                (N285)? mem[31] : 
                (N256)? mem[33] : 
                (N258)? mem[35] : 
                (N260)? mem[37] : 
                (N262)? mem[39] : 
                (N264)? mem[41] : 
                (N266)? mem[43] : 
                (N268)? mem[45] : 
                (N270)? mem[47] : 
                (N272)? mem[49] : 
                (N274)? mem[51] : 
                (N276)? mem[53] : 
                (N278)? mem[55] : 
                (N280)? mem[57] : 
                (N282)? mem[59] : 
                (N284)? mem[61] : 
                (N286)? mem[63] : 1'b0;
  assign N291 = (N255)? mem[0] : 
                (N257)? mem[2] : 
                (N259)? mem[4] : 
                (N261)? mem[6] : 
                (N263)? mem[8] : 
                (N265)? mem[10] : 
                (N267)? mem[12] : 
                (N269)? mem[14] : 
                (N271)? mem[16] : 
                (N273)? mem[18] : 
                (N275)? mem[20] : 
                (N277)? mem[22] : 
                (N279)? mem[24] : 
                (N281)? mem[26] : 
                (N283)? mem[28] : 
                (N285)? mem[30] : 
                (N256)? mem[32] : 
                (N258)? mem[34] : 
                (N260)? mem[36] : 
                (N262)? mem[38] : 
                (N264)? mem[40] : 
                (N266)? mem[42] : 
                (N268)? mem[44] : 
                (N270)? mem[46] : 
                (N272)? mem[48] : 
                (N274)? mem[50] : 
                (N276)? mem[52] : 
                (N278)? mem[54] : 
                (N280)? mem[56] : 
                (N282)? mem[58] : 
                (N284)? mem[60] : 
                (N286)? mem[62] : 1'b0;
  assign N292 = (N255)? mem[1] : 
                (N257)? mem[3] : 
                (N259)? mem[5] : 
                (N261)? mem[7] : 
                (N263)? mem[9] : 
                (N265)? mem[11] : 
                (N267)? mem[13] : 
                (N269)? mem[15] : 
                (N271)? mem[17] : 
                (N273)? mem[19] : 
                (N275)? mem[21] : 
                (N277)? mem[23] : 
                (N279)? mem[25] : 
                (N281)? mem[27] : 
                (N283)? mem[29] : 
                (N285)? mem[31] : 
                (N256)? mem[33] : 
                (N258)? mem[35] : 
                (N260)? mem[37] : 
                (N262)? mem[39] : 
                (N264)? mem[41] : 
                (N266)? mem[43] : 
                (N268)? mem[45] : 
                (N270)? mem[47] : 
                (N272)? mem[49] : 
                (N274)? mem[51] : 
                (N276)? mem[53] : 
                (N278)? mem[55] : 
                (N280)? mem[57] : 
                (N282)? mem[59] : 
                (N284)? mem[61] : 
                (N286)? mem[63] : 1'b0;
  assign N293 = (N255)? mem[0] : 
                (N257)? mem[2] : 
                (N259)? mem[4] : 
                (N261)? mem[6] : 
                (N263)? mem[8] : 
                (N265)? mem[10] : 
                (N267)? mem[12] : 
                (N269)? mem[14] : 
                (N271)? mem[16] : 
                (N273)? mem[18] : 
                (N275)? mem[20] : 
                (N277)? mem[22] : 
                (N279)? mem[24] : 
                (N281)? mem[26] : 
                (N283)? mem[28] : 
                (N285)? mem[30] : 
                (N256)? mem[32] : 
                (N258)? mem[34] : 
                (N260)? mem[36] : 
                (N262)? mem[38] : 
                (N264)? mem[40] : 
                (N266)? mem[42] : 
                (N268)? mem[44] : 
                (N270)? mem[46] : 
                (N272)? mem[48] : 
                (N274)? mem[50] : 
                (N276)? mem[52] : 
                (N278)? mem[54] : 
                (N280)? mem[56] : 
                (N282)? mem[58] : 
                (N284)? mem[60] : 
                (N286)? mem[62] : 1'b0;
  assign N397 = idx_w_i[3] & idx_w_i[4];
  assign N398 = N0 & idx_w_i[4];
  assign N0 = ~idx_w_i[3];
  assign N399 = idx_w_i[3] & N1;
  assign N1 = ~idx_w_i[4];
  assign N400 = N2 & N3;
  assign N2 = ~idx_w_i[3];
  assign N3 = ~idx_w_i[4];
  assign N401 = ~idx_w_i[2];
  assign N402 = idx_w_i[0] & idx_w_i[1];
  assign N403 = N4 & idx_w_i[1];
  assign N4 = ~idx_w_i[0];
  assign N404 = idx_w_i[0] & N5;
  assign N5 = ~idx_w_i[1];
  assign N405 = N6 & N7;
  assign N6 = ~idx_w_i[0];
  assign N7 = ~idx_w_i[1];
  assign N406 = idx_w_i[2] & N402;
  assign N407 = idx_w_i[2] & N403;
  assign N408 = idx_w_i[2] & N404;
  assign N409 = idx_w_i[2] & N405;
  assign N410 = N401 & N402;
  assign N411 = N401 & N403;
  assign N412 = N401 & N404;
  assign N413 = N401 & N405;
  assign N195 = N397 & N406;
  assign N194 = N397 & N407;
  assign N193 = N397 & N408;
  assign N192 = N397 & N409;
  assign N191 = N397 & N410;
  assign N190 = N397 & N411;
  assign N189 = N397 & N412;
  assign N188 = N397 & N413;
  assign N187 = N398 & N406;
  assign N186 = N398 & N407;
  assign N185 = N398 & N408;
  assign N184 = N398 & N409;
  assign N183 = N398 & N410;
  assign N182 = N398 & N411;
  assign N181 = N398 & N412;
  assign N180 = N398 & N413;
  assign N179 = N399 & N406;
  assign N178 = N399 & N407;
  assign N177 = N399 & N408;
  assign N176 = N399 & N409;
  assign N175 = N399 & N410;
  assign N174 = N399 & N411;
  assign N173 = N399 & N412;
  assign N172 = N399 & N413;
  assign N171 = N400 & N406;
  assign N170 = N400 & N407;
  assign N169 = N400 & N408;
  assign N168 = N400 & N409;
  assign N167 = N400 & N410;
  assign N166 = N400 & N411;
  assign N165 = N400 & N412;
  assign N164 = N400 & N413;
  assign { N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N295 } = (N8)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } : 
                                                                                                                                                                                                              (N9)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } : 
                                                                                                                                                                                                              (N10)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } : 
                                                                                                                                                                                                              (N11)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } : 
                                                                                                                                                                                                              (N12)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } : 
                                                                                                                                                                                                              (N13)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } : 
                                                                                                                                                                                                              (N14)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } : 
                                                                                                                                                                                                              (N15)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } : 1'b0;
  assign N8 = N93;
  assign N9 = N96;
  assign N10 = N99;
  assign N11 = N101;
  assign N12 = N104;
  assign N13 = N106;
  assign N14 = N109;
  assign N15 = N111;
  assign { N297, N296 } = (N8)? { N196, 1'b1 } : 
                          (N9)? { N215, 1'b1 } : 
                          (N10)? { N218, 1'b1 } : 
                          (N11)? { N221, 1'b1 } : 
                          (N12)? { N222, N223 } : 
                          (N13)? { N287, N289 } : 
                          (N14)? { N290, N291 } : 
                          (N15)? { N292, N294 } : 1'b0;
  assign { N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N329 } = (N16)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                              (N396)? { N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N295 } : 
                                                                                                                                                                                                              (N86)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = reset_i;
  assign { N331, N330 } = (N16)? { 1'b0, 1'b1 } : 
                          (N396)? { N297, N296 } : 1'b0;
  assign { N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363 } = (N17)? { N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N329 } : 
                                                                                                                                                                                                              (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N17 = en_i;
  assign N18 = N84;
  assign N19 = ~idx_r_i[0];
  assign N20 = ~idx_r_i[1];
  assign N21 = N19 & N20;
  assign N22 = N19 & idx_r_i[1];
  assign N23 = idx_r_i[0] & N20;
  assign N24 = idx_r_i[0] & idx_r_i[1];
  assign N25 = ~idx_r_i[2];
  assign N26 = N21 & N25;
  assign N27 = N21 & idx_r_i[2];
  assign N28 = N23 & N25;
  assign N29 = N23 & idx_r_i[2];
  assign N30 = N22 & N25;
  assign N31 = N22 & idx_r_i[2];
  assign N32 = N24 & N25;
  assign N33 = N24 & idx_r_i[2];
  assign N34 = ~idx_r_i[3];
  assign N35 = N26 & N34;
  assign N36 = N26 & idx_r_i[3];
  assign N37 = N28 & N34;
  assign N38 = N28 & idx_r_i[3];
  assign N39 = N30 & N34;
  assign N40 = N30 & idx_r_i[3];
  assign N41 = N32 & N34;
  assign N42 = N32 & idx_r_i[3];
  assign N43 = N27 & N34;
  assign N44 = N27 & idx_r_i[3];
  assign N45 = N29 & N34;
  assign N46 = N29 & idx_r_i[3];
  assign N47 = N31 & N34;
  assign N48 = N31 & idx_r_i[3];
  assign N49 = N33 & N34;
  assign N50 = N33 & idx_r_i[3];
  assign N51 = ~idx_r_i[4];
  assign N52 = N35 & N51;
  assign N53 = N35 & idx_r_i[4];
  assign N54 = N37 & N51;
  assign N55 = N37 & idx_r_i[4];
  assign N56 = N39 & N51;
  assign N57 = N39 & idx_r_i[4];
  assign N58 = N41 & N51;
  assign N59 = N41 & idx_r_i[4];
  assign N60 = N43 & N51;
  assign N61 = N43 & idx_r_i[4];
  assign N62 = N45 & N51;
  assign N63 = N45 & idx_r_i[4];
  assign N64 = N47 & N51;
  assign N65 = N47 & idx_r_i[4];
  assign N66 = N49 & N51;
  assign N67 = N49 & idx_r_i[4];
  assign N68 = N36 & N51;
  assign N69 = N36 & idx_r_i[4];
  assign N70 = N38 & N51;
  assign N71 = N38 & idx_r_i[4];
  assign N72 = N40 & N51;
  assign N73 = N40 & idx_r_i[4];
  assign N74 = N42 & N51;
  assign N75 = N42 & idx_r_i[4];
  assign N76 = N44 & N51;
  assign N77 = N44 & idx_r_i[4];
  assign N78 = N46 & N51;
  assign N79 = N46 & idx_r_i[4];
  assign N80 = N48 & N51;
  assign N81 = N48 & idx_r_i[4];
  assign N82 = N50 & N51;
  assign N83 = N50 & idx_r_i[4];
  assign N84 = ~en_i;
  assign N85 = w_v_i | reset_i;
  assign N86 = ~N85;
  assign N89 = ~correct_i;
  assign N90 = ~N87;
  assign N91 = ~N88;
  assign N96 = ~N95;
  assign N99 = ~N98;
  assign N101 = ~N100;
  assign N104 = ~N103;
  assign N106 = ~N105;
  assign N109 = ~N108;
  assign N112 = ~idx_w_i[3];
  assign N113 = N231 & N112;
  assign N114 = N233 & N112;
  assign N115 = N235 & N112;
  assign N116 = N237 & N112;
  assign N117 = N232 & N112;
  assign N118 = N234 & N112;
  assign N119 = N236 & N112;
  assign N120 = N238 & N112;
  assign N121 = ~idx_w_i[4];
  assign N122 = N113 & N121;
  assign N123 = N113 & idx_w_i[4];
  assign N124 = N114 & N121;
  assign N125 = N114 & idx_w_i[4];
  assign N126 = N115 & N121;
  assign N127 = N115 & idx_w_i[4];
  assign N128 = N116 & N121;
  assign N129 = N116 & idx_w_i[4];
  assign N130 = N117 & N121;
  assign N131 = N117 & idx_w_i[4];
  assign N132 = N118 & N121;
  assign N133 = N118 & idx_w_i[4];
  assign N134 = N119 & N121;
  assign N135 = N119 & idx_w_i[4];
  assign N136 = N120 & N121;
  assign N137 = N120 & idx_w_i[4];
  assign N138 = N240 & N121;
  assign N139 = N242 & N121;
  assign N140 = N244 & N121;
  assign N141 = N246 & N121;
  assign N142 = N248 & N121;
  assign N143 = N250 & N121;
  assign N144 = N252 & N121;
  assign N145 = N254 & N121;
  assign N147 = N113 & N121;
  assign N148 = N114 & N121;
  assign N149 = N115 & N121;
  assign N150 = N116 & N121;
  assign N151 = N117 & N121;
  assign N152 = N118 & N121;
  assign N153 = N119 & N121;
  assign N154 = N120 & N121;
  assign N155 = N240 & N121;
  assign N156 = N242 & N121;
  assign N157 = N244 & N121;
  assign N158 = N246 & N121;
  assign N159 = N248 & N121;
  assign N160 = N250 & N121;
  assign N161 = N252 & N121;
  assign N162 = N254 & N121;
  assign N196 = N146 ^ N163;
  assign N197 = N239 & N121;
  assign N198 = N241 & N121;
  assign N199 = N243 & N121;
  assign N200 = N245 & N121;
  assign N201 = N247 & N121;
  assign N202 = N249 & N121;
  assign N203 = N251 & N121;
  assign N204 = N253 & N121;
  assign N206 = N239 & N121;
  assign N207 = N241 & N121;
  assign N208 = N243 & N121;
  assign N209 = N245 & N121;
  assign N210 = N247 & N121;
  assign N211 = N249 & N121;
  assign N212 = N251 & N121;
  assign N213 = N253 & N121;
  assign N215 = N205 ^ N214;
  assign N218 = N216 ^ N217;
  assign N221 = N219 ^ N220;
  assign N224 = ~idx_w_i[0];
  assign N225 = ~idx_w_i[1];
  assign N226 = N224 & N225;
  assign N227 = N224 & idx_w_i[1];
  assign N228 = idx_w_i[0] & N225;
  assign N229 = idx_w_i[0] & idx_w_i[1];
  assign N230 = ~idx_w_i[2];
  assign N231 = N226 & N230;
  assign N232 = N226 & idx_w_i[2];
  assign N233 = N228 & N230;
  assign N234 = N228 & idx_w_i[2];
  assign N235 = N227 & N230;
  assign N236 = N227 & idx_w_i[2];
  assign N237 = N229 & N230;
  assign N238 = N229 & idx_w_i[2];
  assign N239 = N231 & N112;
  assign N240 = N231 & idx_w_i[3];
  assign N241 = N233 & N112;
  assign N242 = N233 & idx_w_i[3];
  assign N243 = N235 & N112;
  assign N244 = N235 & idx_w_i[3];
  assign N245 = N237 & N112;
  assign N246 = N237 & idx_w_i[3];
  assign N247 = N232 & N112;
  assign N248 = N232 & idx_w_i[3];
  assign N249 = N234 & N112;
  assign N250 = N234 & idx_w_i[3];
  assign N251 = N236 & N112;
  assign N252 = N236 & idx_w_i[3];
  assign N253 = N238 & N112;
  assign N254 = N238 & idx_w_i[3];
  assign N255 = N239 & N121;
  assign N256 = N239 & idx_w_i[4];
  assign N257 = N241 & N121;
  assign N258 = N241 & idx_w_i[4];
  assign N259 = N243 & N121;
  assign N260 = N243 & idx_w_i[4];
  assign N261 = N245 & N121;
  assign N262 = N245 & idx_w_i[4];
  assign N263 = N247 & N121;
  assign N264 = N247 & idx_w_i[4];
  assign N265 = N249 & N121;
  assign N266 = N249 & idx_w_i[4];
  assign N267 = N251 & N121;
  assign N268 = N251 & idx_w_i[4];
  assign N269 = N253 & N121;
  assign N270 = N253 & idx_w_i[4];
  assign N271 = N240 & N121;
  assign N272 = N240 & idx_w_i[4];
  assign N273 = N242 & N121;
  assign N274 = N242 & idx_w_i[4];
  assign N275 = N244 & N121;
  assign N276 = N244 & idx_w_i[4];
  assign N277 = N246 & N121;
  assign N278 = N246 & idx_w_i[4];
  assign N279 = N248 & N121;
  assign N280 = N248 & idx_w_i[4];
  assign N281 = N250 & N121;
  assign N282 = N250 & idx_w_i[4];
  assign N283 = N252 & N121;
  assign N284 = N252 & idx_w_i[4];
  assign N285 = N254 & N121;
  assign N286 = N254 & idx_w_i[4];
  assign N289 = ~N288;
  assign N294 = ~N293;
  assign N395 = ~reset_i;
  assign N396 = w_v_i & N395;

  always @(posedge clk_i) begin
    if(N394) begin
      { mem[63:62] } <= { N331, N330 };
    end 
    if(N393) begin
      { mem[61:60] } <= { N331, N330 };
    end 
    if(N392) begin
      { mem[59:58] } <= { N331, N330 };
    end 
    if(N391) begin
      { mem[57:56] } <= { N331, N330 };
    end 
    if(N390) begin
      { mem[55:54] } <= { N331, N330 };
    end 
    if(N389) begin
      { mem[53:52] } <= { N331, N330 };
    end 
    if(N388) begin
      { mem[51:50] } <= { N331, N330 };
    end 
    if(N387) begin
      { mem[49:48] } <= { N331, N330 };
    end 
    if(N386) begin
      { mem[47:46] } <= { N331, N330 };
    end 
    if(N385) begin
      { mem[45:44] } <= { N331, N330 };
    end 
    if(N384) begin
      { mem[43:42] } <= { N331, N330 };
    end 
    if(N383) begin
      { mem[41:40] } <= { N331, N330 };
    end 
    if(N382) begin
      { mem[39:38] } <= { N331, N330 };
    end 
    if(N381) begin
      { mem[37:36] } <= { N331, N330 };
    end 
    if(N380) begin
      { mem[35:34] } <= { N331, N330 };
    end 
    if(N379) begin
      { mem[33:32] } <= { N331, N330 };
    end 
    if(N378) begin
      { mem[31:30] } <= { N331, N330 };
    end 
    if(N377) begin
      { mem[29:28] } <= { N331, N330 };
    end 
    if(N376) begin
      { mem[27:26] } <= { N331, N330 };
    end 
    if(N375) begin
      { mem[25:24] } <= { N331, N330 };
    end 
    if(N374) begin
      { mem[23:22] } <= { N331, N330 };
    end 
    if(N373) begin
      { mem[21:20] } <= { N331, N330 };
    end 
    if(N372) begin
      { mem[19:18] } <= { N331, N330 };
    end 
    if(N371) begin
      { mem[17:16] } <= { N331, N330 };
    end 
    if(N370) begin
      { mem[15:14] } <= { N331, N330 };
    end 
    if(N369) begin
      { mem[13:12] } <= { N331, N330 };
    end 
    if(N368) begin
      { mem[11:10] } <= { N331, N330 };
    end 
    if(N367) begin
      { mem[9:8] } <= { N331, N330 };
    end 
    if(N366) begin
      { mem[7:6] } <= { N331, N330 };
    end 
    if(N365) begin
      { mem[5:4] } <= { N331, N330 };
    end 
    if(N364) begin
      { mem[3:2] } <= { N331, N330 };
    end 
    if(N363) begin
      { mem[1:0] } <= { N331, N330 };
    end 
  end


endmodule



module bsg_mem_1rw_sync_width_p64_els_p512_addr_width_lp9
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_i,
  data_o
);

  input [63:0] data_i;
  input [8:0] addr_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [63:0] data_o;

  hard_mem_1rw_d512_w64_wrapper
  macro_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bp_fe_btb_bp_fe_pc_gen_btb_idx_width_lp9_eaddr_width_p64
(
  clk_i,
  reset_i,
  idx_w_i,
  idx_r_i,
  r_v_i,
  w_v_i,
  branch_target_i,
  branch_target_o,
  read_valid_o
);

  input [8:0] idx_w_i;
  input [8:0] idx_r_i;
  input [63:0] branch_target_i;
  output [63:0] branch_target_o;
  input clk_i;
  input reset_i;
  input r_v_i;
  input w_v_i;
  output read_valid_o;
  wire [63:0] branch_target_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,
  N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,
  N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,
  N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,
  N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,
  N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,
  N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,
  N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,
  N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,
  N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,
  N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,
  N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,
  N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,
  N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,
  N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,
  N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,
  N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,
  N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,
  N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,
  N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,
  N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,
  N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,
  N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,
  N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,
  N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,
  N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,
  N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,
  N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,
  N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,
  N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,
  N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,
  N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,
  N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,
  N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,
  N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,
  N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,
  N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,
  N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,
  N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,
  N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,
  N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,
  N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,
  N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,
  N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,
  N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,
  N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,
  N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,
  N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,
  N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,
  N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,
  N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,
  N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,
  N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,
  N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,
  N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,
  N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,
  N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,
  N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,
  N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,
  N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,
  N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,
  N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,
  N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,
  N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,
  N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,
  N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,
  N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,
  N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,
  N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,
  N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,
  N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153;
  wire [8:0] addr;
  reg [511:0] valid;
  reg read_valid_o;
  assign N2080 = (N1568)? valid[0] : 
                 (N1570)? valid[1] : 
                 (N1572)? valid[2] : 
                 (N1574)? valid[3] : 
                 (N1576)? valid[4] : 
                 (N1578)? valid[5] : 
                 (N1580)? valid[6] : 
                 (N1582)? valid[7] : 
                 (N1584)? valid[8] : 
                 (N1586)? valid[9] : 
                 (N1588)? valid[10] : 
                 (N1590)? valid[11] : 
                 (N1592)? valid[12] : 
                 (N1594)? valid[13] : 
                 (N1596)? valid[14] : 
                 (N1598)? valid[15] : 
                 (N1600)? valid[16] : 
                 (N1602)? valid[17] : 
                 (N1604)? valid[18] : 
                 (N1606)? valid[19] : 
                 (N1608)? valid[20] : 
                 (N1610)? valid[21] : 
                 (N1612)? valid[22] : 
                 (N1614)? valid[23] : 
                 (N1616)? valid[24] : 
                 (N1618)? valid[25] : 
                 (N1620)? valid[26] : 
                 (N1622)? valid[27] : 
                 (N1624)? valid[28] : 
                 (N1626)? valid[29] : 
                 (N1628)? valid[30] : 
                 (N1630)? valid[31] : 
                 (N1632)? valid[32] : 
                 (N1634)? valid[33] : 
                 (N1636)? valid[34] : 
                 (N1638)? valid[35] : 
                 (N1640)? valid[36] : 
                 (N1642)? valid[37] : 
                 (N1644)? valid[38] : 
                 (N1646)? valid[39] : 
                 (N1648)? valid[40] : 
                 (N1650)? valid[41] : 
                 (N1652)? valid[42] : 
                 (N1654)? valid[43] : 
                 (N1656)? valid[44] : 
                 (N1658)? valid[45] : 
                 (N1660)? valid[46] : 
                 (N1662)? valid[47] : 
                 (N1664)? valid[48] : 
                 (N1666)? valid[49] : 
                 (N1668)? valid[50] : 
                 (N1670)? valid[51] : 
                 (N1672)? valid[52] : 
                 (N1674)? valid[53] : 
                 (N1676)? valid[54] : 
                 (N1678)? valid[55] : 
                 (N1680)? valid[56] : 
                 (N1682)? valid[57] : 
                 (N1684)? valid[58] : 
                 (N1686)? valid[59] : 
                 (N1688)? valid[60] : 
                 (N1690)? valid[61] : 
                 (N1692)? valid[62] : 
                 (N1694)? valid[63] : 
                 (N1696)? valid[64] : 
                 (N1698)? valid[65] : 
                 (N1700)? valid[66] : 
                 (N1702)? valid[67] : 
                 (N1704)? valid[68] : 
                 (N1706)? valid[69] : 
                 (N1708)? valid[70] : 
                 (N1710)? valid[71] : 
                 (N1712)? valid[72] : 
                 (N1714)? valid[73] : 
                 (N1716)? valid[74] : 
                 (N1718)? valid[75] : 
                 (N1720)? valid[76] : 
                 (N1722)? valid[77] : 
                 (N1724)? valid[78] : 
                 (N1726)? valid[79] : 
                 (N1728)? valid[80] : 
                 (N1730)? valid[81] : 
                 (N1732)? valid[82] : 
                 (N1734)? valid[83] : 
                 (N1736)? valid[84] : 
                 (N1738)? valid[85] : 
                 (N1740)? valid[86] : 
                 (N1742)? valid[87] : 
                 (N1744)? valid[88] : 
                 (N1746)? valid[89] : 
                 (N1748)? valid[90] : 
                 (N1750)? valid[91] : 
                 (N1752)? valid[92] : 
                 (N1754)? valid[93] : 
                 (N1756)? valid[94] : 
                 (N1758)? valid[95] : 
                 (N1760)? valid[96] : 
                 (N1762)? valid[97] : 
                 (N1764)? valid[98] : 
                 (N1766)? valid[99] : 
                 (N1768)? valid[100] : 
                 (N1770)? valid[101] : 
                 (N1772)? valid[102] : 
                 (N1774)? valid[103] : 
                 (N1776)? valid[104] : 
                 (N1778)? valid[105] : 
                 (N1780)? valid[106] : 
                 (N1782)? valid[107] : 
                 (N1784)? valid[108] : 
                 (N1786)? valid[109] : 
                 (N1788)? valid[110] : 
                 (N1790)? valid[111] : 
                 (N1792)? valid[112] : 
                 (N1794)? valid[113] : 
                 (N1796)? valid[114] : 
                 (N1798)? valid[115] : 
                 (N1800)? valid[116] : 
                 (N1802)? valid[117] : 
                 (N1804)? valid[118] : 
                 (N1806)? valid[119] : 
                 (N1808)? valid[120] : 
                 (N1810)? valid[121] : 
                 (N1812)? valid[122] : 
                 (N1814)? valid[123] : 
                 (N1816)? valid[124] : 
                 (N1818)? valid[125] : 
                 (N1820)? valid[126] : 
                 (N1822)? valid[127] : 
                 (N1824)? valid[128] : 
                 (N1826)? valid[129] : 
                 (N1828)? valid[130] : 
                 (N1830)? valid[131] : 
                 (N1832)? valid[132] : 
                 (N1834)? valid[133] : 
                 (N1836)? valid[134] : 
                 (N1838)? valid[135] : 
                 (N1840)? valid[136] : 
                 (N1842)? valid[137] : 
                 (N1844)? valid[138] : 
                 (N1846)? valid[139] : 
                 (N1848)? valid[140] : 
                 (N1850)? valid[141] : 
                 (N1852)? valid[142] : 
                 (N1854)? valid[143] : 
                 (N1856)? valid[144] : 
                 (N1858)? valid[145] : 
                 (N1860)? valid[146] : 
                 (N1862)? valid[147] : 
                 (N1864)? valid[148] : 
                 (N1866)? valid[149] : 
                 (N1868)? valid[150] : 
                 (N1870)? valid[151] : 
                 (N1872)? valid[152] : 
                 (N1874)? valid[153] : 
                 (N1876)? valid[154] : 
                 (N1878)? valid[155] : 
                 (N1880)? valid[156] : 
                 (N1882)? valid[157] : 
                 (N1884)? valid[158] : 
                 (N1886)? valid[159] : 
                 (N1888)? valid[160] : 
                 (N1890)? valid[161] : 
                 (N1892)? valid[162] : 
                 (N1894)? valid[163] : 
                 (N1896)? valid[164] : 
                 (N1898)? valid[165] : 
                 (N1900)? valid[166] : 
                 (N1902)? valid[167] : 
                 (N1904)? valid[168] : 
                 (N1906)? valid[169] : 
                 (N1908)? valid[170] : 
                 (N1910)? valid[171] : 
                 (N1912)? valid[172] : 
                 (N1914)? valid[173] : 
                 (N1916)? valid[174] : 
                 (N1918)? valid[175] : 
                 (N1920)? valid[176] : 
                 (N1922)? valid[177] : 
                 (N1924)? valid[178] : 
                 (N1926)? valid[179] : 
                 (N1928)? valid[180] : 
                 (N1930)? valid[181] : 
                 (N1932)? valid[182] : 
                 (N1934)? valid[183] : 
                 (N1936)? valid[184] : 
                 (N1938)? valid[185] : 
                 (N1940)? valid[186] : 
                 (N1942)? valid[187] : 
                 (N1944)? valid[188] : 
                 (N1946)? valid[189] : 
                 (N1948)? valid[190] : 
                 (N1950)? valid[191] : 
                 (N1952)? valid[192] : 
                 (N1954)? valid[193] : 
                 (N1956)? valid[194] : 
                 (N1958)? valid[195] : 
                 (N1960)? valid[196] : 
                 (N1962)? valid[197] : 
                 (N1964)? valid[198] : 
                 (N1966)? valid[199] : 
                 (N1968)? valid[200] : 
                 (N1970)? valid[201] : 
                 (N1972)? valid[202] : 
                 (N1974)? valid[203] : 
                 (N1976)? valid[204] : 
                 (N1978)? valid[205] : 
                 (N1980)? valid[206] : 
                 (N1982)? valid[207] : 
                 (N1984)? valid[208] : 
                 (N1986)? valid[209] : 
                 (N1988)? valid[210] : 
                 (N1990)? valid[211] : 
                 (N1992)? valid[212] : 
                 (N1994)? valid[213] : 
                 (N1996)? valid[214] : 
                 (N1998)? valid[215] : 
                 (N2000)? valid[216] : 
                 (N2002)? valid[217] : 
                 (N2004)? valid[218] : 
                 (N2006)? valid[219] : 
                 (N2008)? valid[220] : 
                 (N2010)? valid[221] : 
                 (N2012)? valid[222] : 
                 (N2014)? valid[223] : 
                 (N2016)? valid[224] : 
                 (N2018)? valid[225] : 
                 (N2020)? valid[226] : 
                 (N2022)? valid[227] : 
                 (N2024)? valid[228] : 
                 (N2026)? valid[229] : 
                 (N2028)? valid[230] : 
                 (N2030)? valid[231] : 
                 (N2032)? valid[232] : 
                 (N2034)? valid[233] : 
                 (N2036)? valid[234] : 
                 (N2038)? valid[235] : 
                 (N2040)? valid[236] : 
                 (N2042)? valid[237] : 
                 (N2044)? valid[238] : 
                 (N2046)? valid[239] : 
                 (N2048)? valid[240] : 
                 (N2050)? valid[241] : 
                 (N2052)? valid[242] : 
                 (N2054)? valid[243] : 
                 (N2056)? valid[244] : 
                 (N2058)? valid[245] : 
                 (N2060)? valid[246] : 
                 (N2062)? valid[247] : 
                 (N2064)? valid[248] : 
                 (N2066)? valid[249] : 
                 (N2068)? valid[250] : 
                 (N2070)? valid[251] : 
                 (N2072)? valid[252] : 
                 (N2074)? valid[253] : 
                 (N2076)? valid[254] : 
                 (N2078)? valid[255] : 
                 (N1569)? valid[256] : 
                 (N1571)? valid[257] : 
                 (N1573)? valid[258] : 
                 (N1575)? valid[259] : 
                 (N1577)? valid[260] : 
                 (N1579)? valid[261] : 
                 (N1581)? valid[262] : 
                 (N1583)? valid[263] : 
                 (N1585)? valid[264] : 
                 (N1587)? valid[265] : 
                 (N1589)? valid[266] : 
                 (N1591)? valid[267] : 
                 (N1593)? valid[268] : 
                 (N1595)? valid[269] : 
                 (N1597)? valid[270] : 
                 (N1599)? valid[271] : 
                 (N1601)? valid[272] : 
                 (N1603)? valid[273] : 
                 (N1605)? valid[274] : 
                 (N1607)? valid[275] : 
                 (N1609)? valid[276] : 
                 (N1611)? valid[277] : 
                 (N1613)? valid[278] : 
                 (N1615)? valid[279] : 
                 (N1617)? valid[280] : 
                 (N1619)? valid[281] : 
                 (N1621)? valid[282] : 
                 (N1623)? valid[283] : 
                 (N1625)? valid[284] : 
                 (N1627)? valid[285] : 
                 (N1629)? valid[286] : 
                 (N1631)? valid[287] : 
                 (N1633)? valid[288] : 
                 (N1635)? valid[289] : 
                 (N1637)? valid[290] : 
                 (N1639)? valid[291] : 
                 (N1641)? valid[292] : 
                 (N1643)? valid[293] : 
                 (N1645)? valid[294] : 
                 (N1647)? valid[295] : 
                 (N1649)? valid[296] : 
                 (N1651)? valid[297] : 
                 (N1653)? valid[298] : 
                 (N1655)? valid[299] : 
                 (N1657)? valid[300] : 
                 (N1659)? valid[301] : 
                 (N1661)? valid[302] : 
                 (N1663)? valid[303] : 
                 (N1665)? valid[304] : 
                 (N1667)? valid[305] : 
                 (N1669)? valid[306] : 
                 (N1671)? valid[307] : 
                 (N1673)? valid[308] : 
                 (N1675)? valid[309] : 
                 (N1677)? valid[310] : 
                 (N1679)? valid[311] : 
                 (N1681)? valid[312] : 
                 (N1683)? valid[313] : 
                 (N1685)? valid[314] : 
                 (N1687)? valid[315] : 
                 (N1689)? valid[316] : 
                 (N1691)? valid[317] : 
                 (N1693)? valid[318] : 
                 (N1695)? valid[319] : 
                 (N1697)? valid[320] : 
                 (N1699)? valid[321] : 
                 (N1701)? valid[322] : 
                 (N1703)? valid[323] : 
                 (N1705)? valid[324] : 
                 (N1707)? valid[325] : 
                 (N1709)? valid[326] : 
                 (N1711)? valid[327] : 
                 (N1713)? valid[328] : 
                 (N1715)? valid[329] : 
                 (N1717)? valid[330] : 
                 (N1719)? valid[331] : 
                 (N1721)? valid[332] : 
                 (N1723)? valid[333] : 
                 (N1725)? valid[334] : 
                 (N1727)? valid[335] : 
                 (N1729)? valid[336] : 
                 (N1731)? valid[337] : 
                 (N1733)? valid[338] : 
                 (N1735)? valid[339] : 
                 (N1737)? valid[340] : 
                 (N1739)? valid[341] : 
                 (N1741)? valid[342] : 
                 (N1743)? valid[343] : 
                 (N1745)? valid[344] : 
                 (N1747)? valid[345] : 
                 (N1749)? valid[346] : 
                 (N1751)? valid[347] : 
                 (N1753)? valid[348] : 
                 (N1755)? valid[349] : 
                 (N1757)? valid[350] : 
                 (N1759)? valid[351] : 
                 (N1761)? valid[352] : 
                 (N1763)? valid[353] : 
                 (N1765)? valid[354] : 
                 (N1767)? valid[355] : 
                 (N1769)? valid[356] : 
                 (N1771)? valid[357] : 
                 (N1773)? valid[358] : 
                 (N1775)? valid[359] : 
                 (N1777)? valid[360] : 
                 (N1779)? valid[361] : 
                 (N1781)? valid[362] : 
                 (N1783)? valid[363] : 
                 (N1785)? valid[364] : 
                 (N1787)? valid[365] : 
                 (N1789)? valid[366] : 
                 (N1791)? valid[367] : 
                 (N1793)? valid[368] : 
                 (N1795)? valid[369] : 
                 (N1797)? valid[370] : 
                 (N1799)? valid[371] : 
                 (N1801)? valid[372] : 
                 (N1803)? valid[373] : 
                 (N1805)? valid[374] : 
                 (N1807)? valid[375] : 
                 (N1809)? valid[376] : 
                 (N1811)? valid[377] : 
                 (N1813)? valid[378] : 
                 (N1815)? valid[379] : 
                 (N1817)? valid[380] : 
                 (N1819)? valid[381] : 
                 (N1821)? valid[382] : 
                 (N1823)? valid[383] : 
                 (N1825)? valid[384] : 
                 (N1827)? valid[385] : 
                 (N1829)? valid[386] : 
                 (N1831)? valid[387] : 
                 (N1833)? valid[388] : 
                 (N1835)? valid[389] : 
                 (N1837)? valid[390] : 
                 (N1839)? valid[391] : 
                 (N1841)? valid[392] : 
                 (N1843)? valid[393] : 
                 (N1845)? valid[394] : 
                 (N1847)? valid[395] : 
                 (N1849)? valid[396] : 
                 (N1851)? valid[397] : 
                 (N1853)? valid[398] : 
                 (N1855)? valid[399] : 
                 (N1857)? valid[400] : 
                 (N1859)? valid[401] : 
                 (N1861)? valid[402] : 
                 (N1863)? valid[403] : 
                 (N1865)? valid[404] : 
                 (N1867)? valid[405] : 
                 (N1869)? valid[406] : 
                 (N1871)? valid[407] : 
                 (N1873)? valid[408] : 
                 (N1875)? valid[409] : 
                 (N1877)? valid[410] : 
                 (N1879)? valid[411] : 
                 (N1881)? valid[412] : 
                 (N1883)? valid[413] : 
                 (N1885)? valid[414] : 
                 (N1887)? valid[415] : 
                 (N1889)? valid[416] : 
                 (N1891)? valid[417] : 
                 (N1893)? valid[418] : 
                 (N1895)? valid[419] : 
                 (N1897)? valid[420] : 
                 (N1899)? valid[421] : 
                 (N1901)? valid[422] : 
                 (N1903)? valid[423] : 
                 (N1905)? valid[424] : 
                 (N1907)? valid[425] : 
                 (N1909)? valid[426] : 
                 (N1911)? valid[427] : 
                 (N1913)? valid[428] : 
                 (N1915)? valid[429] : 
                 (N1917)? valid[430] : 
                 (N1919)? valid[431] : 
                 (N1921)? valid[432] : 
                 (N1923)? valid[433] : 
                 (N1925)? valid[434] : 
                 (N1927)? valid[435] : 
                 (N1929)? valid[436] : 
                 (N1931)? valid[437] : 
                 (N1933)? valid[438] : 
                 (N1935)? valid[439] : 
                 (N1937)? valid[440] : 
                 (N1939)? valid[441] : 
                 (N1941)? valid[442] : 
                 (N1943)? valid[443] : 
                 (N1945)? valid[444] : 
                 (N1947)? valid[445] : 
                 (N1949)? valid[446] : 
                 (N1951)? valid[447] : 
                 (N1953)? valid[448] : 
                 (N1955)? valid[449] : 
                 (N1957)? valid[450] : 
                 (N1959)? valid[451] : 
                 (N1961)? valid[452] : 
                 (N1963)? valid[453] : 
                 (N1965)? valid[454] : 
                 (N1967)? valid[455] : 
                 (N1969)? valid[456] : 
                 (N1971)? valid[457] : 
                 (N1973)? valid[458] : 
                 (N1975)? valid[459] : 
                 (N1977)? valid[460] : 
                 (N1979)? valid[461] : 
                 (N1981)? valid[462] : 
                 (N1983)? valid[463] : 
                 (N1985)? valid[464] : 
                 (N1987)? valid[465] : 
                 (N1989)? valid[466] : 
                 (N1991)? valid[467] : 
                 (N1993)? valid[468] : 
                 (N1995)? valid[469] : 
                 (N1997)? valid[470] : 
                 (N1999)? valid[471] : 
                 (N2001)? valid[472] : 
                 (N2003)? valid[473] : 
                 (N2005)? valid[474] : 
                 (N2007)? valid[475] : 
                 (N2009)? valid[476] : 
                 (N2011)? valid[477] : 
                 (N2013)? valid[478] : 
                 (N2015)? valid[479] : 
                 (N2017)? valid[480] : 
                 (N2019)? valid[481] : 
                 (N2021)? valid[482] : 
                 (N2023)? valid[483] : 
                 (N2025)? valid[484] : 
                 (N2027)? valid[485] : 
                 (N2029)? valid[486] : 
                 (N2031)? valid[487] : 
                 (N2033)? valid[488] : 
                 (N2035)? valid[489] : 
                 (N2037)? valid[490] : 
                 (N2039)? valid[491] : 
                 (N2041)? valid[492] : 
                 (N2043)? valid[493] : 
                 (N2045)? valid[494] : 
                 (N2047)? valid[495] : 
                 (N2049)? valid[496] : 
                 (N2051)? valid[497] : 
                 (N2053)? valid[498] : 
                 (N2055)? valid[499] : 
                 (N2057)? valid[500] : 
                 (N2059)? valid[501] : 
                 (N2061)? valid[502] : 
                 (N2063)? valid[503] : 
                 (N2065)? valid[504] : 
                 (N2067)? valid[505] : 
                 (N2069)? valid[506] : 
                 (N2071)? valid[507] : 
                 (N2073)? valid[508] : 
                 (N2075)? valid[509] : 
                 (N2077)? valid[510] : 
                 (N2079)? valid[511] : 1'b0;

  bsg_mem_1rw_sync_width_p64_els_p512_addr_width_lp9
  btb_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(branch_target_i),
    .addr_i(addr),
    .v_i(1'b1),
    .w_i(w_v_i),
    .data_o(branch_target_o)
  );

  assign N2081 = idx_w_i[7] & idx_w_i[8];
  assign N2082 = N0 & idx_w_i[8];
  assign N0 = ~idx_w_i[7];
  assign N2083 = idx_w_i[7] & N1;
  assign N1 = ~idx_w_i[8];
  assign N2084 = N2 & N3;
  assign N2 = ~idx_w_i[7];
  assign N3 = ~idx_w_i[8];
  assign N2085 = idx_w_i[5] & idx_w_i[6];
  assign N2086 = N4 & idx_w_i[6];
  assign N4 = ~idx_w_i[5];
  assign N2087 = idx_w_i[5] & N5;
  assign N5 = ~idx_w_i[6];
  assign N2088 = N6 & N7;
  assign N6 = ~idx_w_i[5];
  assign N7 = ~idx_w_i[6];
  assign N2089 = N2081 & N2085;
  assign N2090 = N2081 & N2086;
  assign N2091 = N2081 & N2087;
  assign N2092 = N2081 & N2088;
  assign N2093 = N2082 & N2085;
  assign N2094 = N2082 & N2086;
  assign N2095 = N2082 & N2087;
  assign N2096 = N2082 & N2088;
  assign N2097 = N2083 & N2085;
  assign N2098 = N2083 & N2086;
  assign N2099 = N2083 & N2087;
  assign N2100 = N2083 & N2088;
  assign N2101 = N2084 & N2085;
  assign N2102 = N2084 & N2086;
  assign N2103 = N2084 & N2087;
  assign N2104 = N2084 & N2088;
  assign N2105 = idx_w_i[3] & idx_w_i[4];
  assign N2106 = N8 & idx_w_i[4];
  assign N8 = ~idx_w_i[3];
  assign N2107 = idx_w_i[3] & N9;
  assign N9 = ~idx_w_i[4];
  assign N2108 = N10 & N11;
  assign N10 = ~idx_w_i[3];
  assign N11 = ~idx_w_i[4];
  assign N2109 = ~idx_w_i[2];
  assign N2110 = idx_w_i[0] & idx_w_i[1];
  assign N2111 = N12 & idx_w_i[1];
  assign N12 = ~idx_w_i[0];
  assign N2112 = idx_w_i[0] & N13;
  assign N13 = ~idx_w_i[1];
  assign N2113 = N14 & N15;
  assign N14 = ~idx_w_i[0];
  assign N15 = ~idx_w_i[1];
  assign N2114 = idx_w_i[2] & N2110;
  assign N2115 = idx_w_i[2] & N2111;
  assign N2116 = idx_w_i[2] & N2112;
  assign N2117 = idx_w_i[2] & N2113;
  assign N2118 = N2109 & N2110;
  assign N2119 = N2109 & N2111;
  assign N2120 = N2109 & N2112;
  assign N2121 = N2109 & N2113;
  assign N2122 = N2105 & N2114;
  assign N2123 = N2105 & N2115;
  assign N2124 = N2105 & N2116;
  assign N2125 = N2105 & N2117;
  assign N2126 = N2105 & N2118;
  assign N2127 = N2105 & N2119;
  assign N2128 = N2105 & N2120;
  assign N2129 = N2105 & N2121;
  assign N2130 = N2106 & N2114;
  assign N2131 = N2106 & N2115;
  assign N2132 = N2106 & N2116;
  assign N2133 = N2106 & N2117;
  assign N2134 = N2106 & N2118;
  assign N2135 = N2106 & N2119;
  assign N2136 = N2106 & N2120;
  assign N2137 = N2106 & N2121;
  assign N2138 = N2107 & N2114;
  assign N2139 = N2107 & N2115;
  assign N2140 = N2107 & N2116;
  assign N2141 = N2107 & N2117;
  assign N2142 = N2107 & N2118;
  assign N2143 = N2107 & N2119;
  assign N2144 = N2107 & N2120;
  assign N2145 = N2107 & N2121;
  assign N2146 = N2108 & N2114;
  assign N2147 = N2108 & N2115;
  assign N2148 = N2108 & N2116;
  assign N2149 = N2108 & N2117;
  assign N2150 = N2108 & N2118;
  assign N2151 = N2108 & N2119;
  assign N2152 = N2108 & N2120;
  assign N2153 = N2108 & N2121;
  assign N534 = N2089 & N2122;
  assign N533 = N2089 & N2123;
  assign N532 = N2089 & N2124;
  assign N531 = N2089 & N2125;
  assign N530 = N2089 & N2126;
  assign N529 = N2089 & N2127;
  assign N528 = N2089 & N2128;
  assign N527 = N2089 & N2129;
  assign N526 = N2089 & N2130;
  assign N525 = N2089 & N2131;
  assign N524 = N2089 & N2132;
  assign N523 = N2089 & N2133;
  assign N522 = N2089 & N2134;
  assign N521 = N2089 & N2135;
  assign N520 = N2089 & N2136;
  assign N519 = N2089 & N2137;
  assign N518 = N2089 & N2138;
  assign N517 = N2089 & N2139;
  assign N516 = N2089 & N2140;
  assign N515 = N2089 & N2141;
  assign N514 = N2089 & N2142;
  assign N513 = N2089 & N2143;
  assign N512 = N2089 & N2144;
  assign N511 = N2089 & N2145;
  assign N510 = N2089 & N2146;
  assign N509 = N2089 & N2147;
  assign N508 = N2089 & N2148;
  assign N507 = N2089 & N2149;
  assign N506 = N2089 & N2150;
  assign N505 = N2089 & N2151;
  assign N504 = N2089 & N2152;
  assign N503 = N2089 & N2153;
  assign N502 = N2090 & N2122;
  assign N501 = N2090 & N2123;
  assign N500 = N2090 & N2124;
  assign N499 = N2090 & N2125;
  assign N498 = N2090 & N2126;
  assign N497 = N2090 & N2127;
  assign N496 = N2090 & N2128;
  assign N495 = N2090 & N2129;
  assign N494 = N2090 & N2130;
  assign N493 = N2090 & N2131;
  assign N492 = N2090 & N2132;
  assign N491 = N2090 & N2133;
  assign N490 = N2090 & N2134;
  assign N489 = N2090 & N2135;
  assign N488 = N2090 & N2136;
  assign N487 = N2090 & N2137;
  assign N486 = N2090 & N2138;
  assign N485 = N2090 & N2139;
  assign N484 = N2090 & N2140;
  assign N483 = N2090 & N2141;
  assign N482 = N2090 & N2142;
  assign N481 = N2090 & N2143;
  assign N480 = N2090 & N2144;
  assign N479 = N2090 & N2145;
  assign N478 = N2090 & N2146;
  assign N477 = N2090 & N2147;
  assign N476 = N2090 & N2148;
  assign N475 = N2090 & N2149;
  assign N474 = N2090 & N2150;
  assign N473 = N2090 & N2151;
  assign N472 = N2090 & N2152;
  assign N471 = N2090 & N2153;
  assign N470 = N2091 & N2122;
  assign N469 = N2091 & N2123;
  assign N468 = N2091 & N2124;
  assign N467 = N2091 & N2125;
  assign N466 = N2091 & N2126;
  assign N465 = N2091 & N2127;
  assign N464 = N2091 & N2128;
  assign N463 = N2091 & N2129;
  assign N462 = N2091 & N2130;
  assign N461 = N2091 & N2131;
  assign N460 = N2091 & N2132;
  assign N459 = N2091 & N2133;
  assign N458 = N2091 & N2134;
  assign N457 = N2091 & N2135;
  assign N456 = N2091 & N2136;
  assign N455 = N2091 & N2137;
  assign N454 = N2091 & N2138;
  assign N453 = N2091 & N2139;
  assign N452 = N2091 & N2140;
  assign N451 = N2091 & N2141;
  assign N450 = N2091 & N2142;
  assign N449 = N2091 & N2143;
  assign N448 = N2091 & N2144;
  assign N447 = N2091 & N2145;
  assign N446 = N2091 & N2146;
  assign N445 = N2091 & N2147;
  assign N444 = N2091 & N2148;
  assign N443 = N2091 & N2149;
  assign N442 = N2091 & N2150;
  assign N441 = N2091 & N2151;
  assign N440 = N2091 & N2152;
  assign N439 = N2091 & N2153;
  assign N438 = N2092 & N2122;
  assign N437 = N2092 & N2123;
  assign N436 = N2092 & N2124;
  assign N435 = N2092 & N2125;
  assign N434 = N2092 & N2126;
  assign N433 = N2092 & N2127;
  assign N432 = N2092 & N2128;
  assign N431 = N2092 & N2129;
  assign N430 = N2092 & N2130;
  assign N429 = N2092 & N2131;
  assign N428 = N2092 & N2132;
  assign N427 = N2092 & N2133;
  assign N426 = N2092 & N2134;
  assign N425 = N2092 & N2135;
  assign N424 = N2092 & N2136;
  assign N423 = N2092 & N2137;
  assign N422 = N2092 & N2138;
  assign N421 = N2092 & N2139;
  assign N420 = N2092 & N2140;
  assign N419 = N2092 & N2141;
  assign N418 = N2092 & N2142;
  assign N417 = N2092 & N2143;
  assign N416 = N2092 & N2144;
  assign N415 = N2092 & N2145;
  assign N414 = N2092 & N2146;
  assign N413 = N2092 & N2147;
  assign N412 = N2092 & N2148;
  assign N411 = N2092 & N2149;
  assign N410 = N2092 & N2150;
  assign N409 = N2092 & N2151;
  assign N408 = N2092 & N2152;
  assign N407 = N2092 & N2153;
  assign N406 = N2093 & N2122;
  assign N405 = N2093 & N2123;
  assign N404 = N2093 & N2124;
  assign N403 = N2093 & N2125;
  assign N402 = N2093 & N2126;
  assign N401 = N2093 & N2127;
  assign N400 = N2093 & N2128;
  assign N399 = N2093 & N2129;
  assign N398 = N2093 & N2130;
  assign N397 = N2093 & N2131;
  assign N396 = N2093 & N2132;
  assign N395 = N2093 & N2133;
  assign N394 = N2093 & N2134;
  assign N393 = N2093 & N2135;
  assign N392 = N2093 & N2136;
  assign N391 = N2093 & N2137;
  assign N390 = N2093 & N2138;
  assign N389 = N2093 & N2139;
  assign N388 = N2093 & N2140;
  assign N387 = N2093 & N2141;
  assign N386 = N2093 & N2142;
  assign N385 = N2093 & N2143;
  assign N384 = N2093 & N2144;
  assign N383 = N2093 & N2145;
  assign N382 = N2093 & N2146;
  assign N381 = N2093 & N2147;
  assign N380 = N2093 & N2148;
  assign N379 = N2093 & N2149;
  assign N378 = N2093 & N2150;
  assign N377 = N2093 & N2151;
  assign N376 = N2093 & N2152;
  assign N375 = N2093 & N2153;
  assign N374 = N2094 & N2122;
  assign N373 = N2094 & N2123;
  assign N372 = N2094 & N2124;
  assign N371 = N2094 & N2125;
  assign N370 = N2094 & N2126;
  assign N369 = N2094 & N2127;
  assign N368 = N2094 & N2128;
  assign N367 = N2094 & N2129;
  assign N366 = N2094 & N2130;
  assign N365 = N2094 & N2131;
  assign N364 = N2094 & N2132;
  assign N363 = N2094 & N2133;
  assign N362 = N2094 & N2134;
  assign N361 = N2094 & N2135;
  assign N360 = N2094 & N2136;
  assign N359 = N2094 & N2137;
  assign N358 = N2094 & N2138;
  assign N357 = N2094 & N2139;
  assign N356 = N2094 & N2140;
  assign N355 = N2094 & N2141;
  assign N354 = N2094 & N2142;
  assign N353 = N2094 & N2143;
  assign N352 = N2094 & N2144;
  assign N351 = N2094 & N2145;
  assign N350 = N2094 & N2146;
  assign N349 = N2094 & N2147;
  assign N348 = N2094 & N2148;
  assign N347 = N2094 & N2149;
  assign N346 = N2094 & N2150;
  assign N345 = N2094 & N2151;
  assign N344 = N2094 & N2152;
  assign N343 = N2094 & N2153;
  assign N342 = N2095 & N2122;
  assign N341 = N2095 & N2123;
  assign N340 = N2095 & N2124;
  assign N339 = N2095 & N2125;
  assign N338 = N2095 & N2126;
  assign N337 = N2095 & N2127;
  assign N336 = N2095 & N2128;
  assign N335 = N2095 & N2129;
  assign N334 = N2095 & N2130;
  assign N333 = N2095 & N2131;
  assign N332 = N2095 & N2132;
  assign N331 = N2095 & N2133;
  assign N330 = N2095 & N2134;
  assign N329 = N2095 & N2135;
  assign N328 = N2095 & N2136;
  assign N327 = N2095 & N2137;
  assign N326 = N2095 & N2138;
  assign N325 = N2095 & N2139;
  assign N324 = N2095 & N2140;
  assign N323 = N2095 & N2141;
  assign N322 = N2095 & N2142;
  assign N321 = N2095 & N2143;
  assign N320 = N2095 & N2144;
  assign N319 = N2095 & N2145;
  assign N318 = N2095 & N2146;
  assign N317 = N2095 & N2147;
  assign N316 = N2095 & N2148;
  assign N315 = N2095 & N2149;
  assign N314 = N2095 & N2150;
  assign N313 = N2095 & N2151;
  assign N312 = N2095 & N2152;
  assign N311 = N2095 & N2153;
  assign N310 = N2096 & N2122;
  assign N309 = N2096 & N2123;
  assign N308 = N2096 & N2124;
  assign N307 = N2096 & N2125;
  assign N306 = N2096 & N2126;
  assign N305 = N2096 & N2127;
  assign N304 = N2096 & N2128;
  assign N303 = N2096 & N2129;
  assign N302 = N2096 & N2130;
  assign N301 = N2096 & N2131;
  assign N300 = N2096 & N2132;
  assign N299 = N2096 & N2133;
  assign N298 = N2096 & N2134;
  assign N297 = N2096 & N2135;
  assign N296 = N2096 & N2136;
  assign N295 = N2096 & N2137;
  assign N294 = N2096 & N2138;
  assign N293 = N2096 & N2139;
  assign N292 = N2096 & N2140;
  assign N291 = N2096 & N2141;
  assign N290 = N2096 & N2142;
  assign N289 = N2096 & N2143;
  assign N288 = N2096 & N2144;
  assign N287 = N2096 & N2145;
  assign N286 = N2096 & N2146;
  assign N285 = N2096 & N2147;
  assign N284 = N2096 & N2148;
  assign N283 = N2096 & N2149;
  assign N282 = N2096 & N2150;
  assign N281 = N2096 & N2151;
  assign N280 = N2096 & N2152;
  assign N279 = N2096 & N2153;
  assign N278 = N2097 & N2122;
  assign N277 = N2097 & N2123;
  assign N276 = N2097 & N2124;
  assign N275 = N2097 & N2125;
  assign N274 = N2097 & N2126;
  assign N273 = N2097 & N2127;
  assign N272 = N2097 & N2128;
  assign N271 = N2097 & N2129;
  assign N270 = N2097 & N2130;
  assign N269 = N2097 & N2131;
  assign N268 = N2097 & N2132;
  assign N267 = N2097 & N2133;
  assign N266 = N2097 & N2134;
  assign N265 = N2097 & N2135;
  assign N264 = N2097 & N2136;
  assign N263 = N2097 & N2137;
  assign N262 = N2097 & N2138;
  assign N261 = N2097 & N2139;
  assign N260 = N2097 & N2140;
  assign N259 = N2097 & N2141;
  assign N258 = N2097 & N2142;
  assign N257 = N2097 & N2143;
  assign N256 = N2097 & N2144;
  assign N255 = N2097 & N2145;
  assign N254 = N2097 & N2146;
  assign N253 = N2097 & N2147;
  assign N252 = N2097 & N2148;
  assign N251 = N2097 & N2149;
  assign N250 = N2097 & N2150;
  assign N249 = N2097 & N2151;
  assign N248 = N2097 & N2152;
  assign N247 = N2097 & N2153;
  assign N246 = N2098 & N2122;
  assign N245 = N2098 & N2123;
  assign N244 = N2098 & N2124;
  assign N243 = N2098 & N2125;
  assign N242 = N2098 & N2126;
  assign N241 = N2098 & N2127;
  assign N240 = N2098 & N2128;
  assign N239 = N2098 & N2129;
  assign N238 = N2098 & N2130;
  assign N237 = N2098 & N2131;
  assign N236 = N2098 & N2132;
  assign N235 = N2098 & N2133;
  assign N234 = N2098 & N2134;
  assign N233 = N2098 & N2135;
  assign N232 = N2098 & N2136;
  assign N231 = N2098 & N2137;
  assign N230 = N2098 & N2138;
  assign N229 = N2098 & N2139;
  assign N228 = N2098 & N2140;
  assign N227 = N2098 & N2141;
  assign N226 = N2098 & N2142;
  assign N225 = N2098 & N2143;
  assign N224 = N2098 & N2144;
  assign N223 = N2098 & N2145;
  assign N222 = N2098 & N2146;
  assign N221 = N2098 & N2147;
  assign N220 = N2098 & N2148;
  assign N219 = N2098 & N2149;
  assign N218 = N2098 & N2150;
  assign N217 = N2098 & N2151;
  assign N216 = N2098 & N2152;
  assign N215 = N2098 & N2153;
  assign N214 = N2099 & N2122;
  assign N213 = N2099 & N2123;
  assign N212 = N2099 & N2124;
  assign N211 = N2099 & N2125;
  assign N210 = N2099 & N2126;
  assign N209 = N2099 & N2127;
  assign N208 = N2099 & N2128;
  assign N207 = N2099 & N2129;
  assign N206 = N2099 & N2130;
  assign N205 = N2099 & N2131;
  assign N204 = N2099 & N2132;
  assign N203 = N2099 & N2133;
  assign N202 = N2099 & N2134;
  assign N201 = N2099 & N2135;
  assign N200 = N2099 & N2136;
  assign N199 = N2099 & N2137;
  assign N198 = N2099 & N2138;
  assign N197 = N2099 & N2139;
  assign N196 = N2099 & N2140;
  assign N195 = N2099 & N2141;
  assign N194 = N2099 & N2142;
  assign N193 = N2099 & N2143;
  assign N192 = N2099 & N2144;
  assign N191 = N2099 & N2145;
  assign N190 = N2099 & N2146;
  assign N189 = N2099 & N2147;
  assign N188 = N2099 & N2148;
  assign N187 = N2099 & N2149;
  assign N186 = N2099 & N2150;
  assign N185 = N2099 & N2151;
  assign N184 = N2099 & N2152;
  assign N183 = N2099 & N2153;
  assign N182 = N2100 & N2122;
  assign N181 = N2100 & N2123;
  assign N180 = N2100 & N2124;
  assign N179 = N2100 & N2125;
  assign N178 = N2100 & N2126;
  assign N177 = N2100 & N2127;
  assign N176 = N2100 & N2128;
  assign N175 = N2100 & N2129;
  assign N174 = N2100 & N2130;
  assign N173 = N2100 & N2131;
  assign N172 = N2100 & N2132;
  assign N171 = N2100 & N2133;
  assign N170 = N2100 & N2134;
  assign N169 = N2100 & N2135;
  assign N168 = N2100 & N2136;
  assign N167 = N2100 & N2137;
  assign N166 = N2100 & N2138;
  assign N165 = N2100 & N2139;
  assign N164 = N2100 & N2140;
  assign N163 = N2100 & N2141;
  assign N162 = N2100 & N2142;
  assign N161 = N2100 & N2143;
  assign N160 = N2100 & N2144;
  assign N159 = N2100 & N2145;
  assign N158 = N2100 & N2146;
  assign N157 = N2100 & N2147;
  assign N156 = N2100 & N2148;
  assign N155 = N2100 & N2149;
  assign N154 = N2100 & N2150;
  assign N153 = N2100 & N2151;
  assign N152 = N2100 & N2152;
  assign N151 = N2100 & N2153;
  assign N150 = N2101 & N2122;
  assign N149 = N2101 & N2123;
  assign N148 = N2101 & N2124;
  assign N147 = N2101 & N2125;
  assign N146 = N2101 & N2126;
  assign N145 = N2101 & N2127;
  assign N144 = N2101 & N2128;
  assign N143 = N2101 & N2129;
  assign N142 = N2101 & N2130;
  assign N141 = N2101 & N2131;
  assign N140 = N2101 & N2132;
  assign N139 = N2101 & N2133;
  assign N138 = N2101 & N2134;
  assign N137 = N2101 & N2135;
  assign N136 = N2101 & N2136;
  assign N135 = N2101 & N2137;
  assign N134 = N2101 & N2138;
  assign N133 = N2101 & N2139;
  assign N132 = N2101 & N2140;
  assign N131 = N2101 & N2141;
  assign N130 = N2101 & N2142;
  assign N129 = N2101 & N2143;
  assign N128 = N2101 & N2144;
  assign N127 = N2101 & N2145;
  assign N126 = N2101 & N2146;
  assign N125 = N2101 & N2147;
  assign N124 = N2101 & N2148;
  assign N123 = N2101 & N2149;
  assign N122 = N2101 & N2150;
  assign N121 = N2101 & N2151;
  assign N120 = N2101 & N2152;
  assign N119 = N2101 & N2153;
  assign N118 = N2102 & N2122;
  assign N117 = N2102 & N2123;
  assign N116 = N2102 & N2124;
  assign N115 = N2102 & N2125;
  assign N114 = N2102 & N2126;
  assign N113 = N2102 & N2127;
  assign N112 = N2102 & N2128;
  assign N111 = N2102 & N2129;
  assign N110 = N2102 & N2130;
  assign N109 = N2102 & N2131;
  assign N108 = N2102 & N2132;
  assign N107 = N2102 & N2133;
  assign N106 = N2102 & N2134;
  assign N105 = N2102 & N2135;
  assign N104 = N2102 & N2136;
  assign N103 = N2102 & N2137;
  assign N102 = N2102 & N2138;
  assign N101 = N2102 & N2139;
  assign N100 = N2102 & N2140;
  assign N99 = N2102 & N2141;
  assign N98 = N2102 & N2142;
  assign N97 = N2102 & N2143;
  assign N96 = N2102 & N2144;
  assign N95 = N2102 & N2145;
  assign N94 = N2102 & N2146;
  assign N93 = N2102 & N2147;
  assign N92 = N2102 & N2148;
  assign N91 = N2102 & N2149;
  assign N90 = N2102 & N2150;
  assign N89 = N2102 & N2151;
  assign N88 = N2102 & N2152;
  assign N87 = N2102 & N2153;
  assign N86 = N2103 & N2122;
  assign N85 = N2103 & N2123;
  assign N84 = N2103 & N2124;
  assign N83 = N2103 & N2125;
  assign N82 = N2103 & N2126;
  assign N81 = N2103 & N2127;
  assign N80 = N2103 & N2128;
  assign N79 = N2103 & N2129;
  assign N78 = N2103 & N2130;
  assign N77 = N2103 & N2131;
  assign N76 = N2103 & N2132;
  assign N75 = N2103 & N2133;
  assign N74 = N2103 & N2134;
  assign N73 = N2103 & N2135;
  assign N72 = N2103 & N2136;
  assign N71 = N2103 & N2137;
  assign N70 = N2103 & N2138;
  assign N69 = N2103 & N2139;
  assign N68 = N2103 & N2140;
  assign N67 = N2103 & N2141;
  assign N66 = N2103 & N2142;
  assign N65 = N2103 & N2143;
  assign N64 = N2103 & N2144;
  assign N63 = N2103 & N2145;
  assign N62 = N2103 & N2146;
  assign N61 = N2103 & N2147;
  assign N60 = N2103 & N2148;
  assign N59 = N2103 & N2149;
  assign N58 = N2103 & N2150;
  assign N57 = N2103 & N2151;
  assign N56 = N2103 & N2152;
  assign N55 = N2103 & N2153;
  assign N54 = N2104 & N2122;
  assign N53 = N2104 & N2123;
  assign N52 = N2104 & N2124;
  assign N51 = N2104 & N2125;
  assign N50 = N2104 & N2126;
  assign N49 = N2104 & N2127;
  assign N48 = N2104 & N2128;
  assign N47 = N2104 & N2129;
  assign N46 = N2104 & N2130;
  assign N45 = N2104 & N2131;
  assign N44 = N2104 & N2132;
  assign N43 = N2104 & N2133;
  assign N42 = N2104 & N2134;
  assign N41 = N2104 & N2135;
  assign N40 = N2104 & N2136;
  assign N39 = N2104 & N2137;
  assign N38 = N2104 & N2138;
  assign N37 = N2104 & N2139;
  assign N36 = N2104 & N2140;
  assign N35 = N2104 & N2141;
  assign N34 = N2104 & N2142;
  assign N33 = N2104 & N2143;
  assign N32 = N2104 & N2144;
  assign N31 = N2104 & N2145;
  assign N30 = N2104 & N2146;
  assign N29 = N2104 & N2147;
  assign N28 = N2104 & N2148;
  assign N27 = N2104 & N2149;
  assign N26 = N2104 & N2150;
  assign N25 = N2104 & N2151;
  assign N24 = N2104 & N2152;
  assign N23 = N2104 & N2153;
  assign { N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N540, N539, N538, N537, N536, N535 } = (N16)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N541)? { N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = N19;
  assign addr = (N17)? idx_w_i : 
                (N18)? idx_r_i : 1'b0;
  assign N17 = N1050;
  assign N18 = N1049;
  assign N19 = reset_i;
  assign N20 = w_v_i;
  assign N21 = N20 | N19;
  assign N22 = ~N21;
  assign N1048 = ~N19;
  assign N541 = N20 & N1048;
  assign N1049 = ~w_v_i;
  assign N1050 = w_v_i;
  assign N1051 = ~idx_r_i[0];
  assign N1052 = ~idx_r_i[1];
  assign N1053 = N1051 & N1052;
  assign N1054 = N1051 & idx_r_i[1];
  assign N1055 = idx_r_i[0] & N1052;
  assign N1056 = idx_r_i[0] & idx_r_i[1];
  assign N1057 = ~idx_r_i[2];
  assign N1058 = N1053 & N1057;
  assign N1059 = N1053 & idx_r_i[2];
  assign N1060 = N1055 & N1057;
  assign N1061 = N1055 & idx_r_i[2];
  assign N1062 = N1054 & N1057;
  assign N1063 = N1054 & idx_r_i[2];
  assign N1064 = N1056 & N1057;
  assign N1065 = N1056 & idx_r_i[2];
  assign N1066 = ~idx_r_i[3];
  assign N1067 = N1058 & N1066;
  assign N1068 = N1058 & idx_r_i[3];
  assign N1069 = N1060 & N1066;
  assign N1070 = N1060 & idx_r_i[3];
  assign N1071 = N1062 & N1066;
  assign N1072 = N1062 & idx_r_i[3];
  assign N1073 = N1064 & N1066;
  assign N1074 = N1064 & idx_r_i[3];
  assign N1075 = N1059 & N1066;
  assign N1076 = N1059 & idx_r_i[3];
  assign N1077 = N1061 & N1066;
  assign N1078 = N1061 & idx_r_i[3];
  assign N1079 = N1063 & N1066;
  assign N1080 = N1063 & idx_r_i[3];
  assign N1081 = N1065 & N1066;
  assign N1082 = N1065 & idx_r_i[3];
  assign N1083 = ~idx_r_i[4];
  assign N1084 = N1067 & N1083;
  assign N1085 = N1067 & idx_r_i[4];
  assign N1086 = N1069 & N1083;
  assign N1087 = N1069 & idx_r_i[4];
  assign N1088 = N1071 & N1083;
  assign N1089 = N1071 & idx_r_i[4];
  assign N1090 = N1073 & N1083;
  assign N1091 = N1073 & idx_r_i[4];
  assign N1092 = N1075 & N1083;
  assign N1093 = N1075 & idx_r_i[4];
  assign N1094 = N1077 & N1083;
  assign N1095 = N1077 & idx_r_i[4];
  assign N1096 = N1079 & N1083;
  assign N1097 = N1079 & idx_r_i[4];
  assign N1098 = N1081 & N1083;
  assign N1099 = N1081 & idx_r_i[4];
  assign N1100 = N1068 & N1083;
  assign N1101 = N1068 & idx_r_i[4];
  assign N1102 = N1070 & N1083;
  assign N1103 = N1070 & idx_r_i[4];
  assign N1104 = N1072 & N1083;
  assign N1105 = N1072 & idx_r_i[4];
  assign N1106 = N1074 & N1083;
  assign N1107 = N1074 & idx_r_i[4];
  assign N1108 = N1076 & N1083;
  assign N1109 = N1076 & idx_r_i[4];
  assign N1110 = N1078 & N1083;
  assign N1111 = N1078 & idx_r_i[4];
  assign N1112 = N1080 & N1083;
  assign N1113 = N1080 & idx_r_i[4];
  assign N1114 = N1082 & N1083;
  assign N1115 = N1082 & idx_r_i[4];
  assign N1116 = ~idx_r_i[5];
  assign N1117 = N1084 & N1116;
  assign N1118 = N1084 & idx_r_i[5];
  assign N1119 = N1086 & N1116;
  assign N1120 = N1086 & idx_r_i[5];
  assign N1121 = N1088 & N1116;
  assign N1122 = N1088 & idx_r_i[5];
  assign N1123 = N1090 & N1116;
  assign N1124 = N1090 & idx_r_i[5];
  assign N1125 = N1092 & N1116;
  assign N1126 = N1092 & idx_r_i[5];
  assign N1127 = N1094 & N1116;
  assign N1128 = N1094 & idx_r_i[5];
  assign N1129 = N1096 & N1116;
  assign N1130 = N1096 & idx_r_i[5];
  assign N1131 = N1098 & N1116;
  assign N1132 = N1098 & idx_r_i[5];
  assign N1133 = N1100 & N1116;
  assign N1134 = N1100 & idx_r_i[5];
  assign N1135 = N1102 & N1116;
  assign N1136 = N1102 & idx_r_i[5];
  assign N1137 = N1104 & N1116;
  assign N1138 = N1104 & idx_r_i[5];
  assign N1139 = N1106 & N1116;
  assign N1140 = N1106 & idx_r_i[5];
  assign N1141 = N1108 & N1116;
  assign N1142 = N1108 & idx_r_i[5];
  assign N1143 = N1110 & N1116;
  assign N1144 = N1110 & idx_r_i[5];
  assign N1145 = N1112 & N1116;
  assign N1146 = N1112 & idx_r_i[5];
  assign N1147 = N1114 & N1116;
  assign N1148 = N1114 & idx_r_i[5];
  assign N1149 = N1085 & N1116;
  assign N1150 = N1085 & idx_r_i[5];
  assign N1151 = N1087 & N1116;
  assign N1152 = N1087 & idx_r_i[5];
  assign N1153 = N1089 & N1116;
  assign N1154 = N1089 & idx_r_i[5];
  assign N1155 = N1091 & N1116;
  assign N1156 = N1091 & idx_r_i[5];
  assign N1157 = N1093 & N1116;
  assign N1158 = N1093 & idx_r_i[5];
  assign N1159 = N1095 & N1116;
  assign N1160 = N1095 & idx_r_i[5];
  assign N1161 = N1097 & N1116;
  assign N1162 = N1097 & idx_r_i[5];
  assign N1163 = N1099 & N1116;
  assign N1164 = N1099 & idx_r_i[5];
  assign N1165 = N1101 & N1116;
  assign N1166 = N1101 & idx_r_i[5];
  assign N1167 = N1103 & N1116;
  assign N1168 = N1103 & idx_r_i[5];
  assign N1169 = N1105 & N1116;
  assign N1170 = N1105 & idx_r_i[5];
  assign N1171 = N1107 & N1116;
  assign N1172 = N1107 & idx_r_i[5];
  assign N1173 = N1109 & N1116;
  assign N1174 = N1109 & idx_r_i[5];
  assign N1175 = N1111 & N1116;
  assign N1176 = N1111 & idx_r_i[5];
  assign N1177 = N1113 & N1116;
  assign N1178 = N1113 & idx_r_i[5];
  assign N1179 = N1115 & N1116;
  assign N1180 = N1115 & idx_r_i[5];
  assign N1181 = ~idx_r_i[6];
  assign N1182 = N1117 & N1181;
  assign N1183 = N1117 & idx_r_i[6];
  assign N1184 = N1119 & N1181;
  assign N1185 = N1119 & idx_r_i[6];
  assign N1186 = N1121 & N1181;
  assign N1187 = N1121 & idx_r_i[6];
  assign N1188 = N1123 & N1181;
  assign N1189 = N1123 & idx_r_i[6];
  assign N1190 = N1125 & N1181;
  assign N1191 = N1125 & idx_r_i[6];
  assign N1192 = N1127 & N1181;
  assign N1193 = N1127 & idx_r_i[6];
  assign N1194 = N1129 & N1181;
  assign N1195 = N1129 & idx_r_i[6];
  assign N1196 = N1131 & N1181;
  assign N1197 = N1131 & idx_r_i[6];
  assign N1198 = N1133 & N1181;
  assign N1199 = N1133 & idx_r_i[6];
  assign N1200 = N1135 & N1181;
  assign N1201 = N1135 & idx_r_i[6];
  assign N1202 = N1137 & N1181;
  assign N1203 = N1137 & idx_r_i[6];
  assign N1204 = N1139 & N1181;
  assign N1205 = N1139 & idx_r_i[6];
  assign N1206 = N1141 & N1181;
  assign N1207 = N1141 & idx_r_i[6];
  assign N1208 = N1143 & N1181;
  assign N1209 = N1143 & idx_r_i[6];
  assign N1210 = N1145 & N1181;
  assign N1211 = N1145 & idx_r_i[6];
  assign N1212 = N1147 & N1181;
  assign N1213 = N1147 & idx_r_i[6];
  assign N1214 = N1149 & N1181;
  assign N1215 = N1149 & idx_r_i[6];
  assign N1216 = N1151 & N1181;
  assign N1217 = N1151 & idx_r_i[6];
  assign N1218 = N1153 & N1181;
  assign N1219 = N1153 & idx_r_i[6];
  assign N1220 = N1155 & N1181;
  assign N1221 = N1155 & idx_r_i[6];
  assign N1222 = N1157 & N1181;
  assign N1223 = N1157 & idx_r_i[6];
  assign N1224 = N1159 & N1181;
  assign N1225 = N1159 & idx_r_i[6];
  assign N1226 = N1161 & N1181;
  assign N1227 = N1161 & idx_r_i[6];
  assign N1228 = N1163 & N1181;
  assign N1229 = N1163 & idx_r_i[6];
  assign N1230 = N1165 & N1181;
  assign N1231 = N1165 & idx_r_i[6];
  assign N1232 = N1167 & N1181;
  assign N1233 = N1167 & idx_r_i[6];
  assign N1234 = N1169 & N1181;
  assign N1235 = N1169 & idx_r_i[6];
  assign N1236 = N1171 & N1181;
  assign N1237 = N1171 & idx_r_i[6];
  assign N1238 = N1173 & N1181;
  assign N1239 = N1173 & idx_r_i[6];
  assign N1240 = N1175 & N1181;
  assign N1241 = N1175 & idx_r_i[6];
  assign N1242 = N1177 & N1181;
  assign N1243 = N1177 & idx_r_i[6];
  assign N1244 = N1179 & N1181;
  assign N1245 = N1179 & idx_r_i[6];
  assign N1246 = N1118 & N1181;
  assign N1247 = N1118 & idx_r_i[6];
  assign N1248 = N1120 & N1181;
  assign N1249 = N1120 & idx_r_i[6];
  assign N1250 = N1122 & N1181;
  assign N1251 = N1122 & idx_r_i[6];
  assign N1252 = N1124 & N1181;
  assign N1253 = N1124 & idx_r_i[6];
  assign N1254 = N1126 & N1181;
  assign N1255 = N1126 & idx_r_i[6];
  assign N1256 = N1128 & N1181;
  assign N1257 = N1128 & idx_r_i[6];
  assign N1258 = N1130 & N1181;
  assign N1259 = N1130 & idx_r_i[6];
  assign N1260 = N1132 & N1181;
  assign N1261 = N1132 & idx_r_i[6];
  assign N1262 = N1134 & N1181;
  assign N1263 = N1134 & idx_r_i[6];
  assign N1264 = N1136 & N1181;
  assign N1265 = N1136 & idx_r_i[6];
  assign N1266 = N1138 & N1181;
  assign N1267 = N1138 & idx_r_i[6];
  assign N1268 = N1140 & N1181;
  assign N1269 = N1140 & idx_r_i[6];
  assign N1270 = N1142 & N1181;
  assign N1271 = N1142 & idx_r_i[6];
  assign N1272 = N1144 & N1181;
  assign N1273 = N1144 & idx_r_i[6];
  assign N1274 = N1146 & N1181;
  assign N1275 = N1146 & idx_r_i[6];
  assign N1276 = N1148 & N1181;
  assign N1277 = N1148 & idx_r_i[6];
  assign N1278 = N1150 & N1181;
  assign N1279 = N1150 & idx_r_i[6];
  assign N1280 = N1152 & N1181;
  assign N1281 = N1152 & idx_r_i[6];
  assign N1282 = N1154 & N1181;
  assign N1283 = N1154 & idx_r_i[6];
  assign N1284 = N1156 & N1181;
  assign N1285 = N1156 & idx_r_i[6];
  assign N1286 = N1158 & N1181;
  assign N1287 = N1158 & idx_r_i[6];
  assign N1288 = N1160 & N1181;
  assign N1289 = N1160 & idx_r_i[6];
  assign N1290 = N1162 & N1181;
  assign N1291 = N1162 & idx_r_i[6];
  assign N1292 = N1164 & N1181;
  assign N1293 = N1164 & idx_r_i[6];
  assign N1294 = N1166 & N1181;
  assign N1295 = N1166 & idx_r_i[6];
  assign N1296 = N1168 & N1181;
  assign N1297 = N1168 & idx_r_i[6];
  assign N1298 = N1170 & N1181;
  assign N1299 = N1170 & idx_r_i[6];
  assign N1300 = N1172 & N1181;
  assign N1301 = N1172 & idx_r_i[6];
  assign N1302 = N1174 & N1181;
  assign N1303 = N1174 & idx_r_i[6];
  assign N1304 = N1176 & N1181;
  assign N1305 = N1176 & idx_r_i[6];
  assign N1306 = N1178 & N1181;
  assign N1307 = N1178 & idx_r_i[6];
  assign N1308 = N1180 & N1181;
  assign N1309 = N1180 & idx_r_i[6];
  assign N1310 = ~idx_r_i[7];
  assign N1311 = N1182 & N1310;
  assign N1312 = N1182 & idx_r_i[7];
  assign N1313 = N1184 & N1310;
  assign N1314 = N1184 & idx_r_i[7];
  assign N1315 = N1186 & N1310;
  assign N1316 = N1186 & idx_r_i[7];
  assign N1317 = N1188 & N1310;
  assign N1318 = N1188 & idx_r_i[7];
  assign N1319 = N1190 & N1310;
  assign N1320 = N1190 & idx_r_i[7];
  assign N1321 = N1192 & N1310;
  assign N1322 = N1192 & idx_r_i[7];
  assign N1323 = N1194 & N1310;
  assign N1324 = N1194 & idx_r_i[7];
  assign N1325 = N1196 & N1310;
  assign N1326 = N1196 & idx_r_i[7];
  assign N1327 = N1198 & N1310;
  assign N1328 = N1198 & idx_r_i[7];
  assign N1329 = N1200 & N1310;
  assign N1330 = N1200 & idx_r_i[7];
  assign N1331 = N1202 & N1310;
  assign N1332 = N1202 & idx_r_i[7];
  assign N1333 = N1204 & N1310;
  assign N1334 = N1204 & idx_r_i[7];
  assign N1335 = N1206 & N1310;
  assign N1336 = N1206 & idx_r_i[7];
  assign N1337 = N1208 & N1310;
  assign N1338 = N1208 & idx_r_i[7];
  assign N1339 = N1210 & N1310;
  assign N1340 = N1210 & idx_r_i[7];
  assign N1341 = N1212 & N1310;
  assign N1342 = N1212 & idx_r_i[7];
  assign N1343 = N1214 & N1310;
  assign N1344 = N1214 & idx_r_i[7];
  assign N1345 = N1216 & N1310;
  assign N1346 = N1216 & idx_r_i[7];
  assign N1347 = N1218 & N1310;
  assign N1348 = N1218 & idx_r_i[7];
  assign N1349 = N1220 & N1310;
  assign N1350 = N1220 & idx_r_i[7];
  assign N1351 = N1222 & N1310;
  assign N1352 = N1222 & idx_r_i[7];
  assign N1353 = N1224 & N1310;
  assign N1354 = N1224 & idx_r_i[7];
  assign N1355 = N1226 & N1310;
  assign N1356 = N1226 & idx_r_i[7];
  assign N1357 = N1228 & N1310;
  assign N1358 = N1228 & idx_r_i[7];
  assign N1359 = N1230 & N1310;
  assign N1360 = N1230 & idx_r_i[7];
  assign N1361 = N1232 & N1310;
  assign N1362 = N1232 & idx_r_i[7];
  assign N1363 = N1234 & N1310;
  assign N1364 = N1234 & idx_r_i[7];
  assign N1365 = N1236 & N1310;
  assign N1366 = N1236 & idx_r_i[7];
  assign N1367 = N1238 & N1310;
  assign N1368 = N1238 & idx_r_i[7];
  assign N1369 = N1240 & N1310;
  assign N1370 = N1240 & idx_r_i[7];
  assign N1371 = N1242 & N1310;
  assign N1372 = N1242 & idx_r_i[7];
  assign N1373 = N1244 & N1310;
  assign N1374 = N1244 & idx_r_i[7];
  assign N1375 = N1246 & N1310;
  assign N1376 = N1246 & idx_r_i[7];
  assign N1377 = N1248 & N1310;
  assign N1378 = N1248 & idx_r_i[7];
  assign N1379 = N1250 & N1310;
  assign N1380 = N1250 & idx_r_i[7];
  assign N1381 = N1252 & N1310;
  assign N1382 = N1252 & idx_r_i[7];
  assign N1383 = N1254 & N1310;
  assign N1384 = N1254 & idx_r_i[7];
  assign N1385 = N1256 & N1310;
  assign N1386 = N1256 & idx_r_i[7];
  assign N1387 = N1258 & N1310;
  assign N1388 = N1258 & idx_r_i[7];
  assign N1389 = N1260 & N1310;
  assign N1390 = N1260 & idx_r_i[7];
  assign N1391 = N1262 & N1310;
  assign N1392 = N1262 & idx_r_i[7];
  assign N1393 = N1264 & N1310;
  assign N1394 = N1264 & idx_r_i[7];
  assign N1395 = N1266 & N1310;
  assign N1396 = N1266 & idx_r_i[7];
  assign N1397 = N1268 & N1310;
  assign N1398 = N1268 & idx_r_i[7];
  assign N1399 = N1270 & N1310;
  assign N1400 = N1270 & idx_r_i[7];
  assign N1401 = N1272 & N1310;
  assign N1402 = N1272 & idx_r_i[7];
  assign N1403 = N1274 & N1310;
  assign N1404 = N1274 & idx_r_i[7];
  assign N1405 = N1276 & N1310;
  assign N1406 = N1276 & idx_r_i[7];
  assign N1407 = N1278 & N1310;
  assign N1408 = N1278 & idx_r_i[7];
  assign N1409 = N1280 & N1310;
  assign N1410 = N1280 & idx_r_i[7];
  assign N1411 = N1282 & N1310;
  assign N1412 = N1282 & idx_r_i[7];
  assign N1413 = N1284 & N1310;
  assign N1414 = N1284 & idx_r_i[7];
  assign N1415 = N1286 & N1310;
  assign N1416 = N1286 & idx_r_i[7];
  assign N1417 = N1288 & N1310;
  assign N1418 = N1288 & idx_r_i[7];
  assign N1419 = N1290 & N1310;
  assign N1420 = N1290 & idx_r_i[7];
  assign N1421 = N1292 & N1310;
  assign N1422 = N1292 & idx_r_i[7];
  assign N1423 = N1294 & N1310;
  assign N1424 = N1294 & idx_r_i[7];
  assign N1425 = N1296 & N1310;
  assign N1426 = N1296 & idx_r_i[7];
  assign N1427 = N1298 & N1310;
  assign N1428 = N1298 & idx_r_i[7];
  assign N1429 = N1300 & N1310;
  assign N1430 = N1300 & idx_r_i[7];
  assign N1431 = N1302 & N1310;
  assign N1432 = N1302 & idx_r_i[7];
  assign N1433 = N1304 & N1310;
  assign N1434 = N1304 & idx_r_i[7];
  assign N1435 = N1306 & N1310;
  assign N1436 = N1306 & idx_r_i[7];
  assign N1437 = N1308 & N1310;
  assign N1438 = N1308 & idx_r_i[7];
  assign N1439 = N1183 & N1310;
  assign N1440 = N1183 & idx_r_i[7];
  assign N1441 = N1185 & N1310;
  assign N1442 = N1185 & idx_r_i[7];
  assign N1443 = N1187 & N1310;
  assign N1444 = N1187 & idx_r_i[7];
  assign N1445 = N1189 & N1310;
  assign N1446 = N1189 & idx_r_i[7];
  assign N1447 = N1191 & N1310;
  assign N1448 = N1191 & idx_r_i[7];
  assign N1449 = N1193 & N1310;
  assign N1450 = N1193 & idx_r_i[7];
  assign N1451 = N1195 & N1310;
  assign N1452 = N1195 & idx_r_i[7];
  assign N1453 = N1197 & N1310;
  assign N1454 = N1197 & idx_r_i[7];
  assign N1455 = N1199 & N1310;
  assign N1456 = N1199 & idx_r_i[7];
  assign N1457 = N1201 & N1310;
  assign N1458 = N1201 & idx_r_i[7];
  assign N1459 = N1203 & N1310;
  assign N1460 = N1203 & idx_r_i[7];
  assign N1461 = N1205 & N1310;
  assign N1462 = N1205 & idx_r_i[7];
  assign N1463 = N1207 & N1310;
  assign N1464 = N1207 & idx_r_i[7];
  assign N1465 = N1209 & N1310;
  assign N1466 = N1209 & idx_r_i[7];
  assign N1467 = N1211 & N1310;
  assign N1468 = N1211 & idx_r_i[7];
  assign N1469 = N1213 & N1310;
  assign N1470 = N1213 & idx_r_i[7];
  assign N1471 = N1215 & N1310;
  assign N1472 = N1215 & idx_r_i[7];
  assign N1473 = N1217 & N1310;
  assign N1474 = N1217 & idx_r_i[7];
  assign N1475 = N1219 & N1310;
  assign N1476 = N1219 & idx_r_i[7];
  assign N1477 = N1221 & N1310;
  assign N1478 = N1221 & idx_r_i[7];
  assign N1479 = N1223 & N1310;
  assign N1480 = N1223 & idx_r_i[7];
  assign N1481 = N1225 & N1310;
  assign N1482 = N1225 & idx_r_i[7];
  assign N1483 = N1227 & N1310;
  assign N1484 = N1227 & idx_r_i[7];
  assign N1485 = N1229 & N1310;
  assign N1486 = N1229 & idx_r_i[7];
  assign N1487 = N1231 & N1310;
  assign N1488 = N1231 & idx_r_i[7];
  assign N1489 = N1233 & N1310;
  assign N1490 = N1233 & idx_r_i[7];
  assign N1491 = N1235 & N1310;
  assign N1492 = N1235 & idx_r_i[7];
  assign N1493 = N1237 & N1310;
  assign N1494 = N1237 & idx_r_i[7];
  assign N1495 = N1239 & N1310;
  assign N1496 = N1239 & idx_r_i[7];
  assign N1497 = N1241 & N1310;
  assign N1498 = N1241 & idx_r_i[7];
  assign N1499 = N1243 & N1310;
  assign N1500 = N1243 & idx_r_i[7];
  assign N1501 = N1245 & N1310;
  assign N1502 = N1245 & idx_r_i[7];
  assign N1503 = N1247 & N1310;
  assign N1504 = N1247 & idx_r_i[7];
  assign N1505 = N1249 & N1310;
  assign N1506 = N1249 & idx_r_i[7];
  assign N1507 = N1251 & N1310;
  assign N1508 = N1251 & idx_r_i[7];
  assign N1509 = N1253 & N1310;
  assign N1510 = N1253 & idx_r_i[7];
  assign N1511 = N1255 & N1310;
  assign N1512 = N1255 & idx_r_i[7];
  assign N1513 = N1257 & N1310;
  assign N1514 = N1257 & idx_r_i[7];
  assign N1515 = N1259 & N1310;
  assign N1516 = N1259 & idx_r_i[7];
  assign N1517 = N1261 & N1310;
  assign N1518 = N1261 & idx_r_i[7];
  assign N1519 = N1263 & N1310;
  assign N1520 = N1263 & idx_r_i[7];
  assign N1521 = N1265 & N1310;
  assign N1522 = N1265 & idx_r_i[7];
  assign N1523 = N1267 & N1310;
  assign N1524 = N1267 & idx_r_i[7];
  assign N1525 = N1269 & N1310;
  assign N1526 = N1269 & idx_r_i[7];
  assign N1527 = N1271 & N1310;
  assign N1528 = N1271 & idx_r_i[7];
  assign N1529 = N1273 & N1310;
  assign N1530 = N1273 & idx_r_i[7];
  assign N1531 = N1275 & N1310;
  assign N1532 = N1275 & idx_r_i[7];
  assign N1533 = N1277 & N1310;
  assign N1534 = N1277 & idx_r_i[7];
  assign N1535 = N1279 & N1310;
  assign N1536 = N1279 & idx_r_i[7];
  assign N1537 = N1281 & N1310;
  assign N1538 = N1281 & idx_r_i[7];
  assign N1539 = N1283 & N1310;
  assign N1540 = N1283 & idx_r_i[7];
  assign N1541 = N1285 & N1310;
  assign N1542 = N1285 & idx_r_i[7];
  assign N1543 = N1287 & N1310;
  assign N1544 = N1287 & idx_r_i[7];
  assign N1545 = N1289 & N1310;
  assign N1546 = N1289 & idx_r_i[7];
  assign N1547 = N1291 & N1310;
  assign N1548 = N1291 & idx_r_i[7];
  assign N1549 = N1293 & N1310;
  assign N1550 = N1293 & idx_r_i[7];
  assign N1551 = N1295 & N1310;
  assign N1552 = N1295 & idx_r_i[7];
  assign N1553 = N1297 & N1310;
  assign N1554 = N1297 & idx_r_i[7];
  assign N1555 = N1299 & N1310;
  assign N1556 = N1299 & idx_r_i[7];
  assign N1557 = N1301 & N1310;
  assign N1558 = N1301 & idx_r_i[7];
  assign N1559 = N1303 & N1310;
  assign N1560 = N1303 & idx_r_i[7];
  assign N1561 = N1305 & N1310;
  assign N1562 = N1305 & idx_r_i[7];
  assign N1563 = N1307 & N1310;
  assign N1564 = N1307 & idx_r_i[7];
  assign N1565 = N1309 & N1310;
  assign N1566 = N1309 & idx_r_i[7];
  assign N1567 = ~idx_r_i[8];
  assign N1568 = N1311 & N1567;
  assign N1569 = N1311 & idx_r_i[8];
  assign N1570 = N1313 & N1567;
  assign N1571 = N1313 & idx_r_i[8];
  assign N1572 = N1315 & N1567;
  assign N1573 = N1315 & idx_r_i[8];
  assign N1574 = N1317 & N1567;
  assign N1575 = N1317 & idx_r_i[8];
  assign N1576 = N1319 & N1567;
  assign N1577 = N1319 & idx_r_i[8];
  assign N1578 = N1321 & N1567;
  assign N1579 = N1321 & idx_r_i[8];
  assign N1580 = N1323 & N1567;
  assign N1581 = N1323 & idx_r_i[8];
  assign N1582 = N1325 & N1567;
  assign N1583 = N1325 & idx_r_i[8];
  assign N1584 = N1327 & N1567;
  assign N1585 = N1327 & idx_r_i[8];
  assign N1586 = N1329 & N1567;
  assign N1587 = N1329 & idx_r_i[8];
  assign N1588 = N1331 & N1567;
  assign N1589 = N1331 & idx_r_i[8];
  assign N1590 = N1333 & N1567;
  assign N1591 = N1333 & idx_r_i[8];
  assign N1592 = N1335 & N1567;
  assign N1593 = N1335 & idx_r_i[8];
  assign N1594 = N1337 & N1567;
  assign N1595 = N1337 & idx_r_i[8];
  assign N1596 = N1339 & N1567;
  assign N1597 = N1339 & idx_r_i[8];
  assign N1598 = N1341 & N1567;
  assign N1599 = N1341 & idx_r_i[8];
  assign N1600 = N1343 & N1567;
  assign N1601 = N1343 & idx_r_i[8];
  assign N1602 = N1345 & N1567;
  assign N1603 = N1345 & idx_r_i[8];
  assign N1604 = N1347 & N1567;
  assign N1605 = N1347 & idx_r_i[8];
  assign N1606 = N1349 & N1567;
  assign N1607 = N1349 & idx_r_i[8];
  assign N1608 = N1351 & N1567;
  assign N1609 = N1351 & idx_r_i[8];
  assign N1610 = N1353 & N1567;
  assign N1611 = N1353 & idx_r_i[8];
  assign N1612 = N1355 & N1567;
  assign N1613 = N1355 & idx_r_i[8];
  assign N1614 = N1357 & N1567;
  assign N1615 = N1357 & idx_r_i[8];
  assign N1616 = N1359 & N1567;
  assign N1617 = N1359 & idx_r_i[8];
  assign N1618 = N1361 & N1567;
  assign N1619 = N1361 & idx_r_i[8];
  assign N1620 = N1363 & N1567;
  assign N1621 = N1363 & idx_r_i[8];
  assign N1622 = N1365 & N1567;
  assign N1623 = N1365 & idx_r_i[8];
  assign N1624 = N1367 & N1567;
  assign N1625 = N1367 & idx_r_i[8];
  assign N1626 = N1369 & N1567;
  assign N1627 = N1369 & idx_r_i[8];
  assign N1628 = N1371 & N1567;
  assign N1629 = N1371 & idx_r_i[8];
  assign N1630 = N1373 & N1567;
  assign N1631 = N1373 & idx_r_i[8];
  assign N1632 = N1375 & N1567;
  assign N1633 = N1375 & idx_r_i[8];
  assign N1634 = N1377 & N1567;
  assign N1635 = N1377 & idx_r_i[8];
  assign N1636 = N1379 & N1567;
  assign N1637 = N1379 & idx_r_i[8];
  assign N1638 = N1381 & N1567;
  assign N1639 = N1381 & idx_r_i[8];
  assign N1640 = N1383 & N1567;
  assign N1641 = N1383 & idx_r_i[8];
  assign N1642 = N1385 & N1567;
  assign N1643 = N1385 & idx_r_i[8];
  assign N1644 = N1387 & N1567;
  assign N1645 = N1387 & idx_r_i[8];
  assign N1646 = N1389 & N1567;
  assign N1647 = N1389 & idx_r_i[8];
  assign N1648 = N1391 & N1567;
  assign N1649 = N1391 & idx_r_i[8];
  assign N1650 = N1393 & N1567;
  assign N1651 = N1393 & idx_r_i[8];
  assign N1652 = N1395 & N1567;
  assign N1653 = N1395 & idx_r_i[8];
  assign N1654 = N1397 & N1567;
  assign N1655 = N1397 & idx_r_i[8];
  assign N1656 = N1399 & N1567;
  assign N1657 = N1399 & idx_r_i[8];
  assign N1658 = N1401 & N1567;
  assign N1659 = N1401 & idx_r_i[8];
  assign N1660 = N1403 & N1567;
  assign N1661 = N1403 & idx_r_i[8];
  assign N1662 = N1405 & N1567;
  assign N1663 = N1405 & idx_r_i[8];
  assign N1664 = N1407 & N1567;
  assign N1665 = N1407 & idx_r_i[8];
  assign N1666 = N1409 & N1567;
  assign N1667 = N1409 & idx_r_i[8];
  assign N1668 = N1411 & N1567;
  assign N1669 = N1411 & idx_r_i[8];
  assign N1670 = N1413 & N1567;
  assign N1671 = N1413 & idx_r_i[8];
  assign N1672 = N1415 & N1567;
  assign N1673 = N1415 & idx_r_i[8];
  assign N1674 = N1417 & N1567;
  assign N1675 = N1417 & idx_r_i[8];
  assign N1676 = N1419 & N1567;
  assign N1677 = N1419 & idx_r_i[8];
  assign N1678 = N1421 & N1567;
  assign N1679 = N1421 & idx_r_i[8];
  assign N1680 = N1423 & N1567;
  assign N1681 = N1423 & idx_r_i[8];
  assign N1682 = N1425 & N1567;
  assign N1683 = N1425 & idx_r_i[8];
  assign N1684 = N1427 & N1567;
  assign N1685 = N1427 & idx_r_i[8];
  assign N1686 = N1429 & N1567;
  assign N1687 = N1429 & idx_r_i[8];
  assign N1688 = N1431 & N1567;
  assign N1689 = N1431 & idx_r_i[8];
  assign N1690 = N1433 & N1567;
  assign N1691 = N1433 & idx_r_i[8];
  assign N1692 = N1435 & N1567;
  assign N1693 = N1435 & idx_r_i[8];
  assign N1694 = N1437 & N1567;
  assign N1695 = N1437 & idx_r_i[8];
  assign N1696 = N1439 & N1567;
  assign N1697 = N1439 & idx_r_i[8];
  assign N1698 = N1441 & N1567;
  assign N1699 = N1441 & idx_r_i[8];
  assign N1700 = N1443 & N1567;
  assign N1701 = N1443 & idx_r_i[8];
  assign N1702 = N1445 & N1567;
  assign N1703 = N1445 & idx_r_i[8];
  assign N1704 = N1447 & N1567;
  assign N1705 = N1447 & idx_r_i[8];
  assign N1706 = N1449 & N1567;
  assign N1707 = N1449 & idx_r_i[8];
  assign N1708 = N1451 & N1567;
  assign N1709 = N1451 & idx_r_i[8];
  assign N1710 = N1453 & N1567;
  assign N1711 = N1453 & idx_r_i[8];
  assign N1712 = N1455 & N1567;
  assign N1713 = N1455 & idx_r_i[8];
  assign N1714 = N1457 & N1567;
  assign N1715 = N1457 & idx_r_i[8];
  assign N1716 = N1459 & N1567;
  assign N1717 = N1459 & idx_r_i[8];
  assign N1718 = N1461 & N1567;
  assign N1719 = N1461 & idx_r_i[8];
  assign N1720 = N1463 & N1567;
  assign N1721 = N1463 & idx_r_i[8];
  assign N1722 = N1465 & N1567;
  assign N1723 = N1465 & idx_r_i[8];
  assign N1724 = N1467 & N1567;
  assign N1725 = N1467 & idx_r_i[8];
  assign N1726 = N1469 & N1567;
  assign N1727 = N1469 & idx_r_i[8];
  assign N1728 = N1471 & N1567;
  assign N1729 = N1471 & idx_r_i[8];
  assign N1730 = N1473 & N1567;
  assign N1731 = N1473 & idx_r_i[8];
  assign N1732 = N1475 & N1567;
  assign N1733 = N1475 & idx_r_i[8];
  assign N1734 = N1477 & N1567;
  assign N1735 = N1477 & idx_r_i[8];
  assign N1736 = N1479 & N1567;
  assign N1737 = N1479 & idx_r_i[8];
  assign N1738 = N1481 & N1567;
  assign N1739 = N1481 & idx_r_i[8];
  assign N1740 = N1483 & N1567;
  assign N1741 = N1483 & idx_r_i[8];
  assign N1742 = N1485 & N1567;
  assign N1743 = N1485 & idx_r_i[8];
  assign N1744 = N1487 & N1567;
  assign N1745 = N1487 & idx_r_i[8];
  assign N1746 = N1489 & N1567;
  assign N1747 = N1489 & idx_r_i[8];
  assign N1748 = N1491 & N1567;
  assign N1749 = N1491 & idx_r_i[8];
  assign N1750 = N1493 & N1567;
  assign N1751 = N1493 & idx_r_i[8];
  assign N1752 = N1495 & N1567;
  assign N1753 = N1495 & idx_r_i[8];
  assign N1754 = N1497 & N1567;
  assign N1755 = N1497 & idx_r_i[8];
  assign N1756 = N1499 & N1567;
  assign N1757 = N1499 & idx_r_i[8];
  assign N1758 = N1501 & N1567;
  assign N1759 = N1501 & idx_r_i[8];
  assign N1760 = N1503 & N1567;
  assign N1761 = N1503 & idx_r_i[8];
  assign N1762 = N1505 & N1567;
  assign N1763 = N1505 & idx_r_i[8];
  assign N1764 = N1507 & N1567;
  assign N1765 = N1507 & idx_r_i[8];
  assign N1766 = N1509 & N1567;
  assign N1767 = N1509 & idx_r_i[8];
  assign N1768 = N1511 & N1567;
  assign N1769 = N1511 & idx_r_i[8];
  assign N1770 = N1513 & N1567;
  assign N1771 = N1513 & idx_r_i[8];
  assign N1772 = N1515 & N1567;
  assign N1773 = N1515 & idx_r_i[8];
  assign N1774 = N1517 & N1567;
  assign N1775 = N1517 & idx_r_i[8];
  assign N1776 = N1519 & N1567;
  assign N1777 = N1519 & idx_r_i[8];
  assign N1778 = N1521 & N1567;
  assign N1779 = N1521 & idx_r_i[8];
  assign N1780 = N1523 & N1567;
  assign N1781 = N1523 & idx_r_i[8];
  assign N1782 = N1525 & N1567;
  assign N1783 = N1525 & idx_r_i[8];
  assign N1784 = N1527 & N1567;
  assign N1785 = N1527 & idx_r_i[8];
  assign N1786 = N1529 & N1567;
  assign N1787 = N1529 & idx_r_i[8];
  assign N1788 = N1531 & N1567;
  assign N1789 = N1531 & idx_r_i[8];
  assign N1790 = N1533 & N1567;
  assign N1791 = N1533 & idx_r_i[8];
  assign N1792 = N1535 & N1567;
  assign N1793 = N1535 & idx_r_i[8];
  assign N1794 = N1537 & N1567;
  assign N1795 = N1537 & idx_r_i[8];
  assign N1796 = N1539 & N1567;
  assign N1797 = N1539 & idx_r_i[8];
  assign N1798 = N1541 & N1567;
  assign N1799 = N1541 & idx_r_i[8];
  assign N1800 = N1543 & N1567;
  assign N1801 = N1543 & idx_r_i[8];
  assign N1802 = N1545 & N1567;
  assign N1803 = N1545 & idx_r_i[8];
  assign N1804 = N1547 & N1567;
  assign N1805 = N1547 & idx_r_i[8];
  assign N1806 = N1549 & N1567;
  assign N1807 = N1549 & idx_r_i[8];
  assign N1808 = N1551 & N1567;
  assign N1809 = N1551 & idx_r_i[8];
  assign N1810 = N1553 & N1567;
  assign N1811 = N1553 & idx_r_i[8];
  assign N1812 = N1555 & N1567;
  assign N1813 = N1555 & idx_r_i[8];
  assign N1814 = N1557 & N1567;
  assign N1815 = N1557 & idx_r_i[8];
  assign N1816 = N1559 & N1567;
  assign N1817 = N1559 & idx_r_i[8];
  assign N1818 = N1561 & N1567;
  assign N1819 = N1561 & idx_r_i[8];
  assign N1820 = N1563 & N1567;
  assign N1821 = N1563 & idx_r_i[8];
  assign N1822 = N1565 & N1567;
  assign N1823 = N1565 & idx_r_i[8];
  assign N1824 = N1312 & N1567;
  assign N1825 = N1312 & idx_r_i[8];
  assign N1826 = N1314 & N1567;
  assign N1827 = N1314 & idx_r_i[8];
  assign N1828 = N1316 & N1567;
  assign N1829 = N1316 & idx_r_i[8];
  assign N1830 = N1318 & N1567;
  assign N1831 = N1318 & idx_r_i[8];
  assign N1832 = N1320 & N1567;
  assign N1833 = N1320 & idx_r_i[8];
  assign N1834 = N1322 & N1567;
  assign N1835 = N1322 & idx_r_i[8];
  assign N1836 = N1324 & N1567;
  assign N1837 = N1324 & idx_r_i[8];
  assign N1838 = N1326 & N1567;
  assign N1839 = N1326 & idx_r_i[8];
  assign N1840 = N1328 & N1567;
  assign N1841 = N1328 & idx_r_i[8];
  assign N1842 = N1330 & N1567;
  assign N1843 = N1330 & idx_r_i[8];
  assign N1844 = N1332 & N1567;
  assign N1845 = N1332 & idx_r_i[8];
  assign N1846 = N1334 & N1567;
  assign N1847 = N1334 & idx_r_i[8];
  assign N1848 = N1336 & N1567;
  assign N1849 = N1336 & idx_r_i[8];
  assign N1850 = N1338 & N1567;
  assign N1851 = N1338 & idx_r_i[8];
  assign N1852 = N1340 & N1567;
  assign N1853 = N1340 & idx_r_i[8];
  assign N1854 = N1342 & N1567;
  assign N1855 = N1342 & idx_r_i[8];
  assign N1856 = N1344 & N1567;
  assign N1857 = N1344 & idx_r_i[8];
  assign N1858 = N1346 & N1567;
  assign N1859 = N1346 & idx_r_i[8];
  assign N1860 = N1348 & N1567;
  assign N1861 = N1348 & idx_r_i[8];
  assign N1862 = N1350 & N1567;
  assign N1863 = N1350 & idx_r_i[8];
  assign N1864 = N1352 & N1567;
  assign N1865 = N1352 & idx_r_i[8];
  assign N1866 = N1354 & N1567;
  assign N1867 = N1354 & idx_r_i[8];
  assign N1868 = N1356 & N1567;
  assign N1869 = N1356 & idx_r_i[8];
  assign N1870 = N1358 & N1567;
  assign N1871 = N1358 & idx_r_i[8];
  assign N1872 = N1360 & N1567;
  assign N1873 = N1360 & idx_r_i[8];
  assign N1874 = N1362 & N1567;
  assign N1875 = N1362 & idx_r_i[8];
  assign N1876 = N1364 & N1567;
  assign N1877 = N1364 & idx_r_i[8];
  assign N1878 = N1366 & N1567;
  assign N1879 = N1366 & idx_r_i[8];
  assign N1880 = N1368 & N1567;
  assign N1881 = N1368 & idx_r_i[8];
  assign N1882 = N1370 & N1567;
  assign N1883 = N1370 & idx_r_i[8];
  assign N1884 = N1372 & N1567;
  assign N1885 = N1372 & idx_r_i[8];
  assign N1886 = N1374 & N1567;
  assign N1887 = N1374 & idx_r_i[8];
  assign N1888 = N1376 & N1567;
  assign N1889 = N1376 & idx_r_i[8];
  assign N1890 = N1378 & N1567;
  assign N1891 = N1378 & idx_r_i[8];
  assign N1892 = N1380 & N1567;
  assign N1893 = N1380 & idx_r_i[8];
  assign N1894 = N1382 & N1567;
  assign N1895 = N1382 & idx_r_i[8];
  assign N1896 = N1384 & N1567;
  assign N1897 = N1384 & idx_r_i[8];
  assign N1898 = N1386 & N1567;
  assign N1899 = N1386 & idx_r_i[8];
  assign N1900 = N1388 & N1567;
  assign N1901 = N1388 & idx_r_i[8];
  assign N1902 = N1390 & N1567;
  assign N1903 = N1390 & idx_r_i[8];
  assign N1904 = N1392 & N1567;
  assign N1905 = N1392 & idx_r_i[8];
  assign N1906 = N1394 & N1567;
  assign N1907 = N1394 & idx_r_i[8];
  assign N1908 = N1396 & N1567;
  assign N1909 = N1396 & idx_r_i[8];
  assign N1910 = N1398 & N1567;
  assign N1911 = N1398 & idx_r_i[8];
  assign N1912 = N1400 & N1567;
  assign N1913 = N1400 & idx_r_i[8];
  assign N1914 = N1402 & N1567;
  assign N1915 = N1402 & idx_r_i[8];
  assign N1916 = N1404 & N1567;
  assign N1917 = N1404 & idx_r_i[8];
  assign N1918 = N1406 & N1567;
  assign N1919 = N1406 & idx_r_i[8];
  assign N1920 = N1408 & N1567;
  assign N1921 = N1408 & idx_r_i[8];
  assign N1922 = N1410 & N1567;
  assign N1923 = N1410 & idx_r_i[8];
  assign N1924 = N1412 & N1567;
  assign N1925 = N1412 & idx_r_i[8];
  assign N1926 = N1414 & N1567;
  assign N1927 = N1414 & idx_r_i[8];
  assign N1928 = N1416 & N1567;
  assign N1929 = N1416 & idx_r_i[8];
  assign N1930 = N1418 & N1567;
  assign N1931 = N1418 & idx_r_i[8];
  assign N1932 = N1420 & N1567;
  assign N1933 = N1420 & idx_r_i[8];
  assign N1934 = N1422 & N1567;
  assign N1935 = N1422 & idx_r_i[8];
  assign N1936 = N1424 & N1567;
  assign N1937 = N1424 & idx_r_i[8];
  assign N1938 = N1426 & N1567;
  assign N1939 = N1426 & idx_r_i[8];
  assign N1940 = N1428 & N1567;
  assign N1941 = N1428 & idx_r_i[8];
  assign N1942 = N1430 & N1567;
  assign N1943 = N1430 & idx_r_i[8];
  assign N1944 = N1432 & N1567;
  assign N1945 = N1432 & idx_r_i[8];
  assign N1946 = N1434 & N1567;
  assign N1947 = N1434 & idx_r_i[8];
  assign N1948 = N1436 & N1567;
  assign N1949 = N1436 & idx_r_i[8];
  assign N1950 = N1438 & N1567;
  assign N1951 = N1438 & idx_r_i[8];
  assign N1952 = N1440 & N1567;
  assign N1953 = N1440 & idx_r_i[8];
  assign N1954 = N1442 & N1567;
  assign N1955 = N1442 & idx_r_i[8];
  assign N1956 = N1444 & N1567;
  assign N1957 = N1444 & idx_r_i[8];
  assign N1958 = N1446 & N1567;
  assign N1959 = N1446 & idx_r_i[8];
  assign N1960 = N1448 & N1567;
  assign N1961 = N1448 & idx_r_i[8];
  assign N1962 = N1450 & N1567;
  assign N1963 = N1450 & idx_r_i[8];
  assign N1964 = N1452 & N1567;
  assign N1965 = N1452 & idx_r_i[8];
  assign N1966 = N1454 & N1567;
  assign N1967 = N1454 & idx_r_i[8];
  assign N1968 = N1456 & N1567;
  assign N1969 = N1456 & idx_r_i[8];
  assign N1970 = N1458 & N1567;
  assign N1971 = N1458 & idx_r_i[8];
  assign N1972 = N1460 & N1567;
  assign N1973 = N1460 & idx_r_i[8];
  assign N1974 = N1462 & N1567;
  assign N1975 = N1462 & idx_r_i[8];
  assign N1976 = N1464 & N1567;
  assign N1977 = N1464 & idx_r_i[8];
  assign N1978 = N1466 & N1567;
  assign N1979 = N1466 & idx_r_i[8];
  assign N1980 = N1468 & N1567;
  assign N1981 = N1468 & idx_r_i[8];
  assign N1982 = N1470 & N1567;
  assign N1983 = N1470 & idx_r_i[8];
  assign N1984 = N1472 & N1567;
  assign N1985 = N1472 & idx_r_i[8];
  assign N1986 = N1474 & N1567;
  assign N1987 = N1474 & idx_r_i[8];
  assign N1988 = N1476 & N1567;
  assign N1989 = N1476 & idx_r_i[8];
  assign N1990 = N1478 & N1567;
  assign N1991 = N1478 & idx_r_i[8];
  assign N1992 = N1480 & N1567;
  assign N1993 = N1480 & idx_r_i[8];
  assign N1994 = N1482 & N1567;
  assign N1995 = N1482 & idx_r_i[8];
  assign N1996 = N1484 & N1567;
  assign N1997 = N1484 & idx_r_i[8];
  assign N1998 = N1486 & N1567;
  assign N1999 = N1486 & idx_r_i[8];
  assign N2000 = N1488 & N1567;
  assign N2001 = N1488 & idx_r_i[8];
  assign N2002 = N1490 & N1567;
  assign N2003 = N1490 & idx_r_i[8];
  assign N2004 = N1492 & N1567;
  assign N2005 = N1492 & idx_r_i[8];
  assign N2006 = N1494 & N1567;
  assign N2007 = N1494 & idx_r_i[8];
  assign N2008 = N1496 & N1567;
  assign N2009 = N1496 & idx_r_i[8];
  assign N2010 = N1498 & N1567;
  assign N2011 = N1498 & idx_r_i[8];
  assign N2012 = N1500 & N1567;
  assign N2013 = N1500 & idx_r_i[8];
  assign N2014 = N1502 & N1567;
  assign N2015 = N1502 & idx_r_i[8];
  assign N2016 = N1504 & N1567;
  assign N2017 = N1504 & idx_r_i[8];
  assign N2018 = N1506 & N1567;
  assign N2019 = N1506 & idx_r_i[8];
  assign N2020 = N1508 & N1567;
  assign N2021 = N1508 & idx_r_i[8];
  assign N2022 = N1510 & N1567;
  assign N2023 = N1510 & idx_r_i[8];
  assign N2024 = N1512 & N1567;
  assign N2025 = N1512 & idx_r_i[8];
  assign N2026 = N1514 & N1567;
  assign N2027 = N1514 & idx_r_i[8];
  assign N2028 = N1516 & N1567;
  assign N2029 = N1516 & idx_r_i[8];
  assign N2030 = N1518 & N1567;
  assign N2031 = N1518 & idx_r_i[8];
  assign N2032 = N1520 & N1567;
  assign N2033 = N1520 & idx_r_i[8];
  assign N2034 = N1522 & N1567;
  assign N2035 = N1522 & idx_r_i[8];
  assign N2036 = N1524 & N1567;
  assign N2037 = N1524 & idx_r_i[8];
  assign N2038 = N1526 & N1567;
  assign N2039 = N1526 & idx_r_i[8];
  assign N2040 = N1528 & N1567;
  assign N2041 = N1528 & idx_r_i[8];
  assign N2042 = N1530 & N1567;
  assign N2043 = N1530 & idx_r_i[8];
  assign N2044 = N1532 & N1567;
  assign N2045 = N1532 & idx_r_i[8];
  assign N2046 = N1534 & N1567;
  assign N2047 = N1534 & idx_r_i[8];
  assign N2048 = N1536 & N1567;
  assign N2049 = N1536 & idx_r_i[8];
  assign N2050 = N1538 & N1567;
  assign N2051 = N1538 & idx_r_i[8];
  assign N2052 = N1540 & N1567;
  assign N2053 = N1540 & idx_r_i[8];
  assign N2054 = N1542 & N1567;
  assign N2055 = N1542 & idx_r_i[8];
  assign N2056 = N1544 & N1567;
  assign N2057 = N1544 & idx_r_i[8];
  assign N2058 = N1546 & N1567;
  assign N2059 = N1546 & idx_r_i[8];
  assign N2060 = N1548 & N1567;
  assign N2061 = N1548 & idx_r_i[8];
  assign N2062 = N1550 & N1567;
  assign N2063 = N1550 & idx_r_i[8];
  assign N2064 = N1552 & N1567;
  assign N2065 = N1552 & idx_r_i[8];
  assign N2066 = N1554 & N1567;
  assign N2067 = N1554 & idx_r_i[8];
  assign N2068 = N1556 & N1567;
  assign N2069 = N1556 & idx_r_i[8];
  assign N2070 = N1558 & N1567;
  assign N2071 = N1558 & idx_r_i[8];
  assign N2072 = N1560 & N1567;
  assign N2073 = N1560 & idx_r_i[8];
  assign N2074 = N1562 & N1567;
  assign N2075 = N1562 & idx_r_i[8];
  assign N2076 = N1564 & N1567;
  assign N2077 = N1564 & idx_r_i[8];
  assign N2078 = N1566 & N1567;
  assign N2079 = N1566 & idx_r_i[8];

  always @(posedge clk_i) begin
    if(N1047) begin
      { valid[511:511] } <= { N541 };
    end 
    if(N1046) begin
      { valid[510:510] } <= { N541 };
    end 
    if(N1045) begin
      { valid[509:509] } <= { N541 };
    end 
    if(N1044) begin
      { valid[508:508] } <= { N541 };
    end 
    if(N1043) begin
      { valid[507:507] } <= { N541 };
    end 
    if(N1042) begin
      { valid[506:506] } <= { N541 };
    end 
    if(N1041) begin
      { valid[505:505] } <= { N541 };
    end 
    if(N1040) begin
      { valid[504:504] } <= { N541 };
    end 
    if(N1039) begin
      { valid[503:503] } <= { N541 };
    end 
    if(N1038) begin
      { valid[502:502] } <= { N541 };
    end 
    if(N1037) begin
      { valid[501:501] } <= { N541 };
    end 
    if(N1036) begin
      { valid[500:500] } <= { N541 };
    end 
    if(N1035) begin
      { valid[499:499] } <= { N541 };
    end 
    if(N1034) begin
      { valid[498:498] } <= { N541 };
    end 
    if(N1033) begin
      { valid[497:497] } <= { N541 };
    end 
    if(N1032) begin
      { valid[496:496] } <= { N541 };
    end 
    if(N1031) begin
      { valid[495:495] } <= { N541 };
    end 
    if(N1030) begin
      { valid[494:494] } <= { N541 };
    end 
    if(N1029) begin
      { valid[493:493] } <= { N541 };
    end 
    if(N1028) begin
      { valid[492:492] } <= { N541 };
    end 
    if(N1027) begin
      { valid[491:491] } <= { N541 };
    end 
    if(N1026) begin
      { valid[490:490] } <= { N541 };
    end 
    if(N1025) begin
      { valid[489:489] } <= { N541 };
    end 
    if(N1024) begin
      { valid[488:488] } <= { N541 };
    end 
    if(N1023) begin
      { valid[487:487] } <= { N541 };
    end 
    if(N1022) begin
      { valid[486:486] } <= { N541 };
    end 
    if(N1021) begin
      { valid[485:485] } <= { N541 };
    end 
    if(N1020) begin
      { valid[484:484] } <= { N541 };
    end 
    if(N1019) begin
      { valid[483:483] } <= { N541 };
    end 
    if(N1018) begin
      { valid[482:482] } <= { N541 };
    end 
    if(N1017) begin
      { valid[481:481] } <= { N541 };
    end 
    if(N1016) begin
      { valid[480:480] } <= { N541 };
    end 
    if(N1015) begin
      { valid[479:479] } <= { N541 };
    end 
    if(N1014) begin
      { valid[478:478] } <= { N541 };
    end 
    if(N1013) begin
      { valid[477:477] } <= { N541 };
    end 
    if(N1012) begin
      { valid[476:476] } <= { N541 };
    end 
    if(N1011) begin
      { valid[475:475] } <= { N541 };
    end 
    if(N1010) begin
      { valid[474:474] } <= { N541 };
    end 
    if(N1009) begin
      { valid[473:473] } <= { N541 };
    end 
    if(N1008) begin
      { valid[472:472] } <= { N541 };
    end 
    if(N1007) begin
      { valid[471:471] } <= { N541 };
    end 
    if(N1006) begin
      { valid[470:470] } <= { N541 };
    end 
    if(N1005) begin
      { valid[469:469] } <= { N541 };
    end 
    if(N1004) begin
      { valid[468:468] } <= { N541 };
    end 
    if(N1003) begin
      { valid[467:467] } <= { N541 };
    end 
    if(N1002) begin
      { valid[466:466] } <= { N541 };
    end 
    if(N1001) begin
      { valid[465:465] } <= { N541 };
    end 
    if(N1000) begin
      { valid[464:464] } <= { N541 };
    end 
    if(N999) begin
      { valid[463:463] } <= { N541 };
    end 
    if(N998) begin
      { valid[462:462] } <= { N541 };
    end 
    if(N997) begin
      { valid[461:461] } <= { N541 };
    end 
    if(N996) begin
      { valid[460:460] } <= { N541 };
    end 
    if(N995) begin
      { valid[459:459] } <= { N541 };
    end 
    if(N994) begin
      { valid[458:458] } <= { N541 };
    end 
    if(N993) begin
      { valid[457:457] } <= { N541 };
    end 
    if(N992) begin
      { valid[456:456] } <= { N541 };
    end 
    if(N991) begin
      { valid[455:455] } <= { N541 };
    end 
    if(N990) begin
      { valid[454:454] } <= { N541 };
    end 
    if(N989) begin
      { valid[453:453] } <= { N541 };
    end 
    if(N988) begin
      { valid[452:452] } <= { N541 };
    end 
    if(N987) begin
      { valid[451:451] } <= { N541 };
    end 
    if(N986) begin
      { valid[450:450] } <= { N541 };
    end 
    if(N985) begin
      { valid[449:449] } <= { N541 };
    end 
    if(N984) begin
      { valid[448:448] } <= { N541 };
    end 
    if(N983) begin
      { valid[447:447] } <= { N541 };
    end 
    if(N982) begin
      { valid[446:446] } <= { N541 };
    end 
    if(N981) begin
      { valid[445:445] } <= { N541 };
    end 
    if(N980) begin
      { valid[444:444] } <= { N541 };
    end 
    if(N979) begin
      { valid[443:443] } <= { N541 };
    end 
    if(N978) begin
      { valid[442:442] } <= { N541 };
    end 
    if(N977) begin
      { valid[441:441] } <= { N541 };
    end 
    if(N976) begin
      { valid[440:440] } <= { N541 };
    end 
    if(N975) begin
      { valid[439:439] } <= { N541 };
    end 
    if(N974) begin
      { valid[438:438] } <= { N541 };
    end 
    if(N973) begin
      { valid[437:437] } <= { N541 };
    end 
    if(N972) begin
      { valid[436:436] } <= { N541 };
    end 
    if(N971) begin
      { valid[435:435] } <= { N541 };
    end 
    if(N970) begin
      { valid[434:434] } <= { N541 };
    end 
    if(N969) begin
      { valid[433:433] } <= { N541 };
    end 
    if(N968) begin
      { valid[432:432] } <= { N541 };
    end 
    if(N967) begin
      { valid[431:431] } <= { N541 };
    end 
    if(N966) begin
      { valid[430:430] } <= { N541 };
    end 
    if(N965) begin
      { valid[429:429] } <= { N541 };
    end 
    if(N964) begin
      { valid[428:428] } <= { N541 };
    end 
    if(N963) begin
      { valid[427:427] } <= { N541 };
    end 
    if(N962) begin
      { valid[426:426] } <= { N541 };
    end 
    if(N961) begin
      { valid[425:425] } <= { N541 };
    end 
    if(N960) begin
      { valid[424:424] } <= { N541 };
    end 
    if(N959) begin
      { valid[423:423] } <= { N541 };
    end 
    if(N958) begin
      { valid[422:422] } <= { N541 };
    end 
    if(N957) begin
      { valid[421:421] } <= { N541 };
    end 
    if(N956) begin
      { valid[420:420] } <= { N541 };
    end 
    if(N955) begin
      { valid[419:419] } <= { N541 };
    end 
    if(N954) begin
      { valid[418:418] } <= { N541 };
    end 
    if(N953) begin
      { valid[417:417] } <= { N541 };
    end 
    if(N952) begin
      { valid[416:416] } <= { N541 };
    end 
    if(N951) begin
      { valid[415:415] } <= { N541 };
    end 
    if(N950) begin
      { valid[414:414] } <= { N541 };
    end 
    if(N949) begin
      { valid[413:413] } <= { N541 };
    end 
    if(N948) begin
      { valid[412:412] } <= { N541 };
    end 
    if(N947) begin
      { valid[411:411] } <= { N541 };
    end 
    if(N946) begin
      { valid[410:410] } <= { N541 };
    end 
    if(N945) begin
      { valid[409:409] } <= { N541 };
    end 
    if(N944) begin
      { valid[408:408] } <= { N541 };
    end 
    if(N943) begin
      { valid[407:407] } <= { N541 };
    end 
    if(N942) begin
      { valid[406:406] } <= { N541 };
    end 
    if(N941) begin
      { valid[405:405] } <= { N541 };
    end 
    if(N940) begin
      { valid[404:404] } <= { N541 };
    end 
    if(N939) begin
      { valid[403:403] } <= { N541 };
    end 
    if(N938) begin
      { valid[402:402] } <= { N541 };
    end 
    if(N937) begin
      { valid[401:401] } <= { N541 };
    end 
    if(N936) begin
      { valid[400:400] } <= { N541 };
    end 
    if(N935) begin
      { valid[399:399] } <= { N541 };
    end 
    if(N934) begin
      { valid[398:398] } <= { N541 };
    end 
    if(N933) begin
      { valid[397:397] } <= { N541 };
    end 
    if(N932) begin
      { valid[396:396] } <= { N541 };
    end 
    if(N931) begin
      { valid[395:395] } <= { N541 };
    end 
    if(N930) begin
      { valid[394:394] } <= { N541 };
    end 
    if(N929) begin
      { valid[393:393] } <= { N541 };
    end 
    if(N928) begin
      { valid[392:392] } <= { N541 };
    end 
    if(N927) begin
      { valid[391:391] } <= { N541 };
    end 
    if(N926) begin
      { valid[390:390] } <= { N541 };
    end 
    if(N925) begin
      { valid[389:389] } <= { N541 };
    end 
    if(N924) begin
      { valid[388:388] } <= { N541 };
    end 
    if(N923) begin
      { valid[387:387] } <= { N541 };
    end 
    if(N922) begin
      { valid[386:386] } <= { N541 };
    end 
    if(N921) begin
      { valid[385:385] } <= { N541 };
    end 
    if(N920) begin
      { valid[384:384] } <= { N541 };
    end 
    if(N919) begin
      { valid[383:383] } <= { N541 };
    end 
    if(N918) begin
      { valid[382:382] } <= { N541 };
    end 
    if(N917) begin
      { valid[381:381] } <= { N541 };
    end 
    if(N916) begin
      { valid[380:380] } <= { N541 };
    end 
    if(N915) begin
      { valid[379:379] } <= { N541 };
    end 
    if(N914) begin
      { valid[378:378] } <= { N541 };
    end 
    if(N913) begin
      { valid[377:377] } <= { N541 };
    end 
    if(N912) begin
      { valid[376:376] } <= { N541 };
    end 
    if(N911) begin
      { valid[375:375] } <= { N541 };
    end 
    if(N910) begin
      { valid[374:374] } <= { N541 };
    end 
    if(N909) begin
      { valid[373:373] } <= { N541 };
    end 
    if(N908) begin
      { valid[372:372] } <= { N541 };
    end 
    if(N907) begin
      { valid[371:371] } <= { N541 };
    end 
    if(N906) begin
      { valid[370:370] } <= { N541 };
    end 
    if(N905) begin
      { valid[369:369] } <= { N541 };
    end 
    if(N904) begin
      { valid[368:368] } <= { N541 };
    end 
    if(N903) begin
      { valid[367:367] } <= { N541 };
    end 
    if(N902) begin
      { valid[366:366] } <= { N541 };
    end 
    if(N901) begin
      { valid[365:365] } <= { N541 };
    end 
    if(N900) begin
      { valid[364:364] } <= { N541 };
    end 
    if(N899) begin
      { valid[363:363] } <= { N541 };
    end 
    if(N898) begin
      { valid[362:362] } <= { N541 };
    end 
    if(N897) begin
      { valid[361:361] } <= { N541 };
    end 
    if(N896) begin
      { valid[360:360] } <= { N541 };
    end 
    if(N895) begin
      { valid[359:359] } <= { N541 };
    end 
    if(N894) begin
      { valid[358:358] } <= { N541 };
    end 
    if(N893) begin
      { valid[357:357] } <= { N541 };
    end 
    if(N892) begin
      { valid[356:356] } <= { N541 };
    end 
    if(N891) begin
      { valid[355:355] } <= { N541 };
    end 
    if(N890) begin
      { valid[354:354] } <= { N541 };
    end 
    if(N889) begin
      { valid[353:353] } <= { N541 };
    end 
    if(N888) begin
      { valid[352:352] } <= { N541 };
    end 
    if(N887) begin
      { valid[351:351] } <= { N541 };
    end 
    if(N886) begin
      { valid[350:350] } <= { N541 };
    end 
    if(N885) begin
      { valid[349:349] } <= { N541 };
    end 
    if(N884) begin
      { valid[348:348] } <= { N541 };
    end 
    if(N883) begin
      { valid[347:347] } <= { N541 };
    end 
    if(N882) begin
      { valid[346:346] } <= { N541 };
    end 
    if(N881) begin
      { valid[345:345] } <= { N541 };
    end 
    if(N880) begin
      { valid[344:344] } <= { N541 };
    end 
    if(N879) begin
      { valid[343:343] } <= { N541 };
    end 
    if(N878) begin
      { valid[342:342] } <= { N541 };
    end 
    if(N877) begin
      { valid[341:341] } <= { N541 };
    end 
    if(N876) begin
      { valid[340:340] } <= { N541 };
    end 
    if(N875) begin
      { valid[339:339] } <= { N541 };
    end 
    if(N874) begin
      { valid[338:338] } <= { N541 };
    end 
    if(N873) begin
      { valid[337:337] } <= { N541 };
    end 
    if(N872) begin
      { valid[336:336] } <= { N541 };
    end 
    if(N871) begin
      { valid[335:335] } <= { N541 };
    end 
    if(N870) begin
      { valid[334:334] } <= { N541 };
    end 
    if(N869) begin
      { valid[333:333] } <= { N541 };
    end 
    if(N868) begin
      { valid[332:332] } <= { N541 };
    end 
    if(N867) begin
      { valid[331:331] } <= { N541 };
    end 
    if(N866) begin
      { valid[330:330] } <= { N541 };
    end 
    if(N865) begin
      { valid[329:329] } <= { N541 };
    end 
    if(N864) begin
      { valid[328:328] } <= { N541 };
    end 
    if(N863) begin
      { valid[327:327] } <= { N541 };
    end 
    if(N862) begin
      { valid[326:326] } <= { N541 };
    end 
    if(N861) begin
      { valid[325:325] } <= { N541 };
    end 
    if(N860) begin
      { valid[324:324] } <= { N541 };
    end 
    if(N859) begin
      { valid[323:323] } <= { N541 };
    end 
    if(N858) begin
      { valid[322:322] } <= { N541 };
    end 
    if(N857) begin
      { valid[321:321] } <= { N541 };
    end 
    if(N856) begin
      { valid[320:320] } <= { N541 };
    end 
    if(N855) begin
      { valid[319:319] } <= { N541 };
    end 
    if(N854) begin
      { valid[318:318] } <= { N541 };
    end 
    if(N853) begin
      { valid[317:317] } <= { N541 };
    end 
    if(N852) begin
      { valid[316:316] } <= { N541 };
    end 
    if(N851) begin
      { valid[315:315] } <= { N541 };
    end 
    if(N850) begin
      { valid[314:314] } <= { N541 };
    end 
    if(N849) begin
      { valid[313:313] } <= { N541 };
    end 
    if(N848) begin
      { valid[312:312] } <= { N541 };
    end 
    if(N847) begin
      { valid[311:311] } <= { N541 };
    end 
    if(N846) begin
      { valid[310:310] } <= { N541 };
    end 
    if(N845) begin
      { valid[309:309] } <= { N541 };
    end 
    if(N844) begin
      { valid[308:308] } <= { N541 };
    end 
    if(N843) begin
      { valid[307:307] } <= { N541 };
    end 
    if(N842) begin
      { valid[306:306] } <= { N541 };
    end 
    if(N841) begin
      { valid[305:305] } <= { N541 };
    end 
    if(N840) begin
      { valid[304:304] } <= { N541 };
    end 
    if(N839) begin
      { valid[303:303] } <= { N541 };
    end 
    if(N838) begin
      { valid[302:302] } <= { N541 };
    end 
    if(N837) begin
      { valid[301:301] } <= { N541 };
    end 
    if(N836) begin
      { valid[300:300] } <= { N541 };
    end 
    if(N835) begin
      { valid[299:299] } <= { N541 };
    end 
    if(N834) begin
      { valid[298:298] } <= { N541 };
    end 
    if(N833) begin
      { valid[297:297] } <= { N541 };
    end 
    if(N832) begin
      { valid[296:296] } <= { N541 };
    end 
    if(N831) begin
      { valid[295:295] } <= { N541 };
    end 
    if(N830) begin
      { valid[294:294] } <= { N541 };
    end 
    if(N829) begin
      { valid[293:293] } <= { N541 };
    end 
    if(N828) begin
      { valid[292:292] } <= { N541 };
    end 
    if(N827) begin
      { valid[291:291] } <= { N541 };
    end 
    if(N826) begin
      { valid[290:290] } <= { N541 };
    end 
    if(N825) begin
      { valid[289:289] } <= { N541 };
    end 
    if(N824) begin
      { valid[288:288] } <= { N541 };
    end 
    if(N823) begin
      { valid[287:287] } <= { N541 };
    end 
    if(N822) begin
      { valid[286:286] } <= { N541 };
    end 
    if(N821) begin
      { valid[285:285] } <= { N541 };
    end 
    if(N820) begin
      { valid[284:284] } <= { N541 };
    end 
    if(N819) begin
      { valid[283:283] } <= { N541 };
    end 
    if(N818) begin
      { valid[282:282] } <= { N541 };
    end 
    if(N817) begin
      { valid[281:281] } <= { N541 };
    end 
    if(N816) begin
      { valid[280:280] } <= { N541 };
    end 
    if(N815) begin
      { valid[279:279] } <= { N541 };
    end 
    if(N814) begin
      { valid[278:278] } <= { N541 };
    end 
    if(N813) begin
      { valid[277:277] } <= { N541 };
    end 
    if(N812) begin
      { valid[276:276] } <= { N541 };
    end 
    if(N811) begin
      { valid[275:275] } <= { N541 };
    end 
    if(N810) begin
      { valid[274:274] } <= { N541 };
    end 
    if(N809) begin
      { valid[273:273] } <= { N541 };
    end 
    if(N808) begin
      { valid[272:272] } <= { N541 };
    end 
    if(N807) begin
      { valid[271:271] } <= { N541 };
    end 
    if(N806) begin
      { valid[270:270] } <= { N541 };
    end 
    if(N805) begin
      { valid[269:269] } <= { N541 };
    end 
    if(N804) begin
      { valid[268:268] } <= { N541 };
    end 
    if(N803) begin
      { valid[267:267] } <= { N541 };
    end 
    if(N802) begin
      { valid[266:266] } <= { N541 };
    end 
    if(N801) begin
      { valid[265:265] } <= { N541 };
    end 
    if(N800) begin
      { valid[264:264] } <= { N541 };
    end 
    if(N799) begin
      { valid[263:263] } <= { N541 };
    end 
    if(N798) begin
      { valid[262:262] } <= { N541 };
    end 
    if(N797) begin
      { valid[261:261] } <= { N541 };
    end 
    if(N796) begin
      { valid[260:260] } <= { N541 };
    end 
    if(N795) begin
      { valid[259:259] } <= { N541 };
    end 
    if(N794) begin
      { valid[258:258] } <= { N541 };
    end 
    if(N793) begin
      { valid[257:257] } <= { N541 };
    end 
    if(N792) begin
      { valid[256:256] } <= { N541 };
    end 
    if(N791) begin
      { valid[255:255] } <= { N541 };
    end 
    if(N790) begin
      { valid[254:254] } <= { N541 };
    end 
    if(N789) begin
      { valid[253:253] } <= { N541 };
    end 
    if(N788) begin
      { valid[252:252] } <= { N541 };
    end 
    if(N787) begin
      { valid[251:251] } <= { N541 };
    end 
    if(N786) begin
      { valid[250:250] } <= { N541 };
    end 
    if(N785) begin
      { valid[249:249] } <= { N541 };
    end 
    if(N784) begin
      { valid[248:248] } <= { N541 };
    end 
    if(N783) begin
      { valid[247:247] } <= { N541 };
    end 
    if(N782) begin
      { valid[246:246] } <= { N541 };
    end 
    if(N781) begin
      { valid[245:245] } <= { N541 };
    end 
    if(N780) begin
      { valid[244:244] } <= { N541 };
    end 
    if(N779) begin
      { valid[243:243] } <= { N541 };
    end 
    if(N778) begin
      { valid[242:242] } <= { N541 };
    end 
    if(N777) begin
      { valid[241:241] } <= { N541 };
    end 
    if(N776) begin
      { valid[240:240] } <= { N541 };
    end 
    if(N775) begin
      { valid[239:239] } <= { N541 };
    end 
    if(N774) begin
      { valid[238:238] } <= { N541 };
    end 
    if(N773) begin
      { valid[237:237] } <= { N541 };
    end 
    if(N772) begin
      { valid[236:236] } <= { N541 };
    end 
    if(N771) begin
      { valid[235:235] } <= { N541 };
    end 
    if(N770) begin
      { valid[234:234] } <= { N541 };
    end 
    if(N769) begin
      { valid[233:233] } <= { N541 };
    end 
    if(N768) begin
      { valid[232:232] } <= { N541 };
    end 
    if(N767) begin
      { valid[231:231] } <= { N541 };
    end 
    if(N766) begin
      { valid[230:230] } <= { N541 };
    end 
    if(N765) begin
      { valid[229:229] } <= { N541 };
    end 
    if(N764) begin
      { valid[228:228] } <= { N541 };
    end 
    if(N763) begin
      { valid[227:227] } <= { N541 };
    end 
    if(N762) begin
      { valid[226:226] } <= { N541 };
    end 
    if(N761) begin
      { valid[225:225] } <= { N541 };
    end 
    if(N760) begin
      { valid[224:224] } <= { N541 };
    end 
    if(N759) begin
      { valid[223:223] } <= { N541 };
    end 
    if(N758) begin
      { valid[222:222] } <= { N541 };
    end 
    if(N757) begin
      { valid[221:221] } <= { N541 };
    end 
    if(N756) begin
      { valid[220:220] } <= { N541 };
    end 
    if(N755) begin
      { valid[219:219] } <= { N541 };
    end 
    if(N754) begin
      { valid[218:218] } <= { N541 };
    end 
    if(N753) begin
      { valid[217:217] } <= { N541 };
    end 
    if(N752) begin
      { valid[216:216] } <= { N541 };
    end 
    if(N751) begin
      { valid[215:215] } <= { N541 };
    end 
    if(N750) begin
      { valid[214:214] } <= { N541 };
    end 
    if(N749) begin
      { valid[213:213] } <= { N541 };
    end 
    if(N748) begin
      { valid[212:212] } <= { N541 };
    end 
    if(N747) begin
      { valid[211:211] } <= { N541 };
    end 
    if(N746) begin
      { valid[210:210] } <= { N541 };
    end 
    if(N745) begin
      { valid[209:209] } <= { N541 };
    end 
    if(N744) begin
      { valid[208:208] } <= { N541 };
    end 
    if(N743) begin
      { valid[207:207] } <= { N541 };
    end 
    if(N742) begin
      { valid[206:206] } <= { N541 };
    end 
    if(N741) begin
      { valid[205:205] } <= { N541 };
    end 
    if(N740) begin
      { valid[204:204] } <= { N541 };
    end 
    if(N739) begin
      { valid[203:203] } <= { N541 };
    end 
    if(N738) begin
      { valid[202:202] } <= { N541 };
    end 
    if(N737) begin
      { valid[201:201] } <= { N541 };
    end 
    if(N736) begin
      { valid[200:200] } <= { N541 };
    end 
    if(N735) begin
      { valid[199:199] } <= { N541 };
    end 
    if(N734) begin
      { valid[198:198] } <= { N541 };
    end 
    if(N733) begin
      { valid[197:197] } <= { N541 };
    end 
    if(N732) begin
      { valid[196:196] } <= { N541 };
    end 
    if(N731) begin
      { valid[195:195] } <= { N541 };
    end 
    if(N730) begin
      { valid[194:194] } <= { N541 };
    end 
    if(N729) begin
      { valid[193:193] } <= { N541 };
    end 
    if(N728) begin
      { valid[192:192] } <= { N541 };
    end 
    if(N727) begin
      { valid[191:191] } <= { N541 };
    end 
    if(N726) begin
      { valid[190:190] } <= { N541 };
    end 
    if(N725) begin
      { valid[189:189] } <= { N541 };
    end 
    if(N724) begin
      { valid[188:188] } <= { N541 };
    end 
    if(N723) begin
      { valid[187:187] } <= { N541 };
    end 
    if(N722) begin
      { valid[186:186] } <= { N541 };
    end 
    if(N721) begin
      { valid[185:185] } <= { N541 };
    end 
    if(N720) begin
      { valid[184:184] } <= { N541 };
    end 
    if(N719) begin
      { valid[183:183] } <= { N541 };
    end 
    if(N718) begin
      { valid[182:182] } <= { N541 };
    end 
    if(N717) begin
      { valid[181:181] } <= { N541 };
    end 
    if(N716) begin
      { valid[180:180] } <= { N541 };
    end 
    if(N715) begin
      { valid[179:179] } <= { N541 };
    end 
    if(N714) begin
      { valid[178:178] } <= { N541 };
    end 
    if(N713) begin
      { valid[177:177] } <= { N541 };
    end 
    if(N712) begin
      { valid[176:176] } <= { N541 };
    end 
    if(N711) begin
      { valid[175:175] } <= { N541 };
    end 
    if(N710) begin
      { valid[174:174] } <= { N541 };
    end 
    if(N709) begin
      { valid[173:173] } <= { N541 };
    end 
    if(N708) begin
      { valid[172:172] } <= { N541 };
    end 
    if(N707) begin
      { valid[171:171] } <= { N541 };
    end 
    if(N706) begin
      { valid[170:170] } <= { N541 };
    end 
    if(N705) begin
      { valid[169:169] } <= { N541 };
    end 
    if(N704) begin
      { valid[168:168] } <= { N541 };
    end 
    if(N703) begin
      { valid[167:167] } <= { N541 };
    end 
    if(N702) begin
      { valid[166:166] } <= { N541 };
    end 
    if(N701) begin
      { valid[165:165] } <= { N541 };
    end 
    if(N700) begin
      { valid[164:164] } <= { N541 };
    end 
    if(N699) begin
      { valid[163:163] } <= { N541 };
    end 
    if(N698) begin
      { valid[162:162] } <= { N541 };
    end 
    if(N697) begin
      { valid[161:161] } <= { N541 };
    end 
    if(N696) begin
      { valid[160:160] } <= { N541 };
    end 
    if(N695) begin
      { valid[159:159] } <= { N541 };
    end 
    if(N694) begin
      { valid[158:158] } <= { N541 };
    end 
    if(N693) begin
      { valid[157:157] } <= { N541 };
    end 
    if(N692) begin
      { valid[156:156] } <= { N541 };
    end 
    if(N691) begin
      { valid[155:155] } <= { N541 };
    end 
    if(N690) begin
      { valid[154:154] } <= { N541 };
    end 
    if(N689) begin
      { valid[153:153] } <= { N541 };
    end 
    if(N688) begin
      { valid[152:152] } <= { N541 };
    end 
    if(N687) begin
      { valid[151:151] } <= { N541 };
    end 
    if(N686) begin
      { valid[150:150] } <= { N541 };
    end 
    if(N685) begin
      { valid[149:149] } <= { N541 };
    end 
    if(N684) begin
      { valid[148:148] } <= { N541 };
    end 
    if(N683) begin
      { valid[147:147] } <= { N541 };
    end 
    if(N682) begin
      { valid[146:146] } <= { N541 };
    end 
    if(N681) begin
      { valid[145:145] } <= { N541 };
    end 
    if(N680) begin
      { valid[144:144] } <= { N541 };
    end 
    if(N679) begin
      { valid[143:143] } <= { N541 };
    end 
    if(N678) begin
      { valid[142:142] } <= { N541 };
    end 
    if(N677) begin
      { valid[141:141] } <= { N541 };
    end 
    if(N676) begin
      { valid[140:140] } <= { N541 };
    end 
    if(N675) begin
      { valid[139:139] } <= { N541 };
    end 
    if(N674) begin
      { valid[138:138] } <= { N541 };
    end 
    if(N673) begin
      { valid[137:137] } <= { N541 };
    end 
    if(N672) begin
      { valid[136:136] } <= { N541 };
    end 
    if(N671) begin
      { valid[135:135] } <= { N541 };
    end 
    if(N670) begin
      { valid[134:134] } <= { N541 };
    end 
    if(N669) begin
      { valid[133:133] } <= { N541 };
    end 
    if(N668) begin
      { valid[132:132] } <= { N541 };
    end 
    if(N667) begin
      { valid[131:131] } <= { N541 };
    end 
    if(N666) begin
      { valid[130:130] } <= { N541 };
    end 
    if(N665) begin
      { valid[129:129] } <= { N541 };
    end 
    if(N664) begin
      { valid[128:128] } <= { N541 };
    end 
    if(N663) begin
      { valid[127:127] } <= { N541 };
    end 
    if(N662) begin
      { valid[126:126] } <= { N541 };
    end 
    if(N661) begin
      { valid[125:125] } <= { N541 };
    end 
    if(N660) begin
      { valid[124:124] } <= { N541 };
    end 
    if(N659) begin
      { valid[123:123] } <= { N541 };
    end 
    if(N658) begin
      { valid[122:122] } <= { N541 };
    end 
    if(N657) begin
      { valid[121:121] } <= { N541 };
    end 
    if(N656) begin
      { valid[120:120] } <= { N541 };
    end 
    if(N655) begin
      { valid[119:119] } <= { N541 };
    end 
    if(N654) begin
      { valid[118:118] } <= { N541 };
    end 
    if(N653) begin
      { valid[117:117] } <= { N541 };
    end 
    if(N652) begin
      { valid[116:116] } <= { N541 };
    end 
    if(N651) begin
      { valid[115:115] } <= { N541 };
    end 
    if(N650) begin
      { valid[114:114] } <= { N541 };
    end 
    if(N649) begin
      { valid[113:113] } <= { N541 };
    end 
    if(N648) begin
      { valid[112:112] } <= { N541 };
    end 
    if(N647) begin
      { valid[111:111] } <= { N541 };
    end 
    if(N646) begin
      { valid[110:110] } <= { N541 };
    end 
    if(N645) begin
      { valid[109:109] } <= { N541 };
    end 
    if(N644) begin
      { valid[108:108] } <= { N541 };
    end 
    if(N643) begin
      { valid[107:107] } <= { N541 };
    end 
    if(N642) begin
      { valid[106:106] } <= { N541 };
    end 
    if(N641) begin
      { valid[105:105] } <= { N541 };
    end 
    if(N640) begin
      { valid[104:104] } <= { N541 };
    end 
    if(N639) begin
      { valid[103:103] } <= { N541 };
    end 
    if(N638) begin
      { valid[102:102] } <= { N541 };
    end 
    if(N637) begin
      { valid[101:101] } <= { N541 };
    end 
    if(N636) begin
      { valid[100:100] } <= { N541 };
    end 
    if(N635) begin
      { valid[99:99] } <= { N541 };
    end 
    if(N634) begin
      { valid[98:98] } <= { N541 };
    end 
    if(N633) begin
      { valid[97:97] } <= { N541 };
    end 
    if(N632) begin
      { valid[96:96] } <= { N541 };
    end 
    if(N631) begin
      { valid[95:95] } <= { N541 };
    end 
    if(N630) begin
      { valid[94:94] } <= { N541 };
    end 
    if(N629) begin
      { valid[93:93] } <= { N541 };
    end 
    if(N628) begin
      { valid[92:92] } <= { N541 };
    end 
    if(N627) begin
      { valid[91:91] } <= { N541 };
    end 
    if(N626) begin
      { valid[90:90] } <= { N541 };
    end 
    if(N625) begin
      { valid[89:89] } <= { N541 };
    end 
    if(N624) begin
      { valid[88:88] } <= { N541 };
    end 
    if(N623) begin
      { valid[87:87] } <= { N541 };
    end 
    if(N622) begin
      { valid[86:86] } <= { N541 };
    end 
    if(N621) begin
      { valid[85:85] } <= { N541 };
    end 
    if(N620) begin
      { valid[84:84] } <= { N541 };
    end 
    if(N619) begin
      { valid[83:83] } <= { N541 };
    end 
    if(N618) begin
      { valid[82:82] } <= { N541 };
    end 
    if(N617) begin
      { valid[81:81] } <= { N541 };
    end 
    if(N616) begin
      { valid[80:80] } <= { N541 };
    end 
    if(N615) begin
      { valid[79:79] } <= { N541 };
    end 
    if(N614) begin
      { valid[78:78] } <= { N541 };
    end 
    if(N613) begin
      { valid[77:77] } <= { N541 };
    end 
    if(N612) begin
      { valid[76:76] } <= { N541 };
    end 
    if(N611) begin
      { valid[75:75] } <= { N541 };
    end 
    if(N610) begin
      { valid[74:74] } <= { N541 };
    end 
    if(N609) begin
      { valid[73:73] } <= { N541 };
    end 
    if(N608) begin
      { valid[72:72] } <= { N541 };
    end 
    if(N607) begin
      { valid[71:71] } <= { N541 };
    end 
    if(N606) begin
      { valid[70:70] } <= { N541 };
    end 
    if(N605) begin
      { valid[69:69] } <= { N541 };
    end 
    if(N604) begin
      { valid[68:68] } <= { N541 };
    end 
    if(N603) begin
      { valid[67:67] } <= { N541 };
    end 
    if(N602) begin
      { valid[66:66] } <= { N541 };
    end 
    if(N601) begin
      { valid[65:65] } <= { N541 };
    end 
    if(N600) begin
      { valid[64:64] } <= { N541 };
    end 
    if(N599) begin
      { valid[63:63] } <= { N541 };
    end 
    if(N598) begin
      { valid[62:62] } <= { N541 };
    end 
    if(N597) begin
      { valid[61:61] } <= { N541 };
    end 
    if(N596) begin
      { valid[60:60] } <= { N541 };
    end 
    if(N595) begin
      { valid[59:59] } <= { N541 };
    end 
    if(N594) begin
      { valid[58:58] } <= { N541 };
    end 
    if(N593) begin
      { valid[57:57] } <= { N541 };
    end 
    if(N592) begin
      { valid[56:56] } <= { N541 };
    end 
    if(N591) begin
      { valid[55:55] } <= { N541 };
    end 
    if(N590) begin
      { valid[54:54] } <= { N541 };
    end 
    if(N589) begin
      { valid[53:53] } <= { N541 };
    end 
    if(N588) begin
      { valid[52:52] } <= { N541 };
    end 
    if(N587) begin
      { valid[51:51] } <= { N541 };
    end 
    if(N586) begin
      { valid[50:50] } <= { N541 };
    end 
    if(N585) begin
      { valid[49:49] } <= { N541 };
    end 
    if(N584) begin
      { valid[48:48] } <= { N541 };
    end 
    if(N583) begin
      { valid[47:47] } <= { N541 };
    end 
    if(N582) begin
      { valid[46:46] } <= { N541 };
    end 
    if(N581) begin
      { valid[45:45] } <= { N541 };
    end 
    if(N580) begin
      { valid[44:44] } <= { N541 };
    end 
    if(N579) begin
      { valid[43:43] } <= { N541 };
    end 
    if(N578) begin
      { valid[42:42] } <= { N541 };
    end 
    if(N577) begin
      { valid[41:41] } <= { N541 };
    end 
    if(N576) begin
      { valid[40:40] } <= { N541 };
    end 
    if(N575) begin
      { valid[39:39] } <= { N541 };
    end 
    if(N574) begin
      { valid[38:38] } <= { N541 };
    end 
    if(N573) begin
      { valid[37:37] } <= { N541 };
    end 
    if(N572) begin
      { valid[36:36] } <= { N541 };
    end 
    if(N571) begin
      { valid[35:35] } <= { N541 };
    end 
    if(N570) begin
      { valid[34:34] } <= { N541 };
    end 
    if(N569) begin
      { valid[33:33] } <= { N541 };
    end 
    if(N568) begin
      { valid[32:32] } <= { N541 };
    end 
    if(N567) begin
      { valid[31:31] } <= { N541 };
    end 
    if(N566) begin
      { valid[30:30] } <= { N541 };
    end 
    if(N565) begin
      { valid[29:29] } <= { N541 };
    end 
    if(N564) begin
      { valid[28:28] } <= { N541 };
    end 
    if(N563) begin
      { valid[27:27] } <= { N541 };
    end 
    if(N562) begin
      { valid[26:26] } <= { N541 };
    end 
    if(N561) begin
      { valid[25:25] } <= { N541 };
    end 
    if(N560) begin
      { valid[24:24] } <= { N541 };
    end 
    if(N559) begin
      { valid[23:23] } <= { N541 };
    end 
    if(N558) begin
      { valid[22:22] } <= { N541 };
    end 
    if(N557) begin
      { valid[21:21] } <= { N541 };
    end 
    if(N556) begin
      { valid[20:20] } <= { N541 };
    end 
    if(N555) begin
      { valid[19:19] } <= { N541 };
    end 
    if(N554) begin
      { valid[18:18] } <= { N541 };
    end 
    if(N553) begin
      { valid[17:17] } <= { N541 };
    end 
    if(N552) begin
      { valid[16:16] } <= { N541 };
    end 
    if(N551) begin
      { valid[15:15] } <= { N541 };
    end 
    if(N550) begin
      { valid[14:14] } <= { N541 };
    end 
    if(N549) begin
      { valid[13:13] } <= { N541 };
    end 
    if(N548) begin
      { valid[12:12] } <= { N541 };
    end 
    if(N547) begin
      { valid[11:11] } <= { N541 };
    end 
    if(N546) begin
      { valid[10:10] } <= { N541 };
    end 
    if(N545) begin
      { valid[9:9] } <= { N541 };
    end 
    if(N544) begin
      { valid[8:8] } <= { N541 };
    end 
    if(N543) begin
      { valid[7:7] } <= { N541 };
    end 
    if(N542) begin
      { valid[6:6] } <= { N541 };
    end 
    if(N540) begin
      { valid[5:5] } <= { N541 };
    end 
    if(N539) begin
      { valid[4:4] } <= { N541 };
    end 
    if(N538) begin
      { valid[3:3] } <= { N541 };
    end 
    if(N537) begin
      { valid[2:2] } <= { N541 };
    end 
    if(N536) begin
      { valid[1:1] } <= { N541 };
    end 
    if(N535) begin
      { valid[0:0] } <= { N541 };
    end 
    if(1'b1) begin
      read_valid_o <= N2080;
    end 
  end


endmodule



module bp_fe_branch_predictor_eaddr_width_p64_btb_indx_width_p9_bht_indx_width_p5_ras_addr_width_p22
(
  clk_i,
  reset_i,
  attaboy_i,
  r_v_i,
  w_v_i,
  pc_queue_i,
  pc_cmd_i,
  pc_fwd_i,
  branch_metadata_fwd_i,
  predict_o,
  pc_o,
  branch_metadata_fwd_o
);

  input [63:0] pc_queue_i;
  input [63:0] pc_cmd_i;
  input [63:0] pc_fwd_i;
  input [35:0] branch_metadata_fwd_i;
  output [63:0] pc_o;
  output [35:0] branch_metadata_fwd_o;
  input clk_i;
  input reset_i;
  input attaboy_i;
  input r_v_i;
  input w_v_i;
  output predict_o;
  wire [63:0] pc_o;
  wire [35:0] branch_metadata_fwd_o;
  wire predict_o,predict,read_valid;
  assign branch_metadata_fwd_o[0] = 1'b0;
  assign branch_metadata_fwd_o[1] = 1'b0;
  assign branch_metadata_fwd_o[2] = 1'b0;
  assign branch_metadata_fwd_o[3] = 1'b0;
  assign branch_metadata_fwd_o[4] = 1'b0;
  assign branch_metadata_fwd_o[5] = 1'b0;
  assign branch_metadata_fwd_o[6] = 1'b0;
  assign branch_metadata_fwd_o[7] = 1'b0;
  assign branch_metadata_fwd_o[8] = 1'b0;
  assign branch_metadata_fwd_o[9] = 1'b0;
  assign branch_metadata_fwd_o[10] = 1'b0;
  assign branch_metadata_fwd_o[11] = 1'b0;
  assign branch_metadata_fwd_o[12] = 1'b0;
  assign branch_metadata_fwd_o[13] = 1'b0;
  assign branch_metadata_fwd_o[14] = 1'b0;
  assign branch_metadata_fwd_o[15] = 1'b0;
  assign branch_metadata_fwd_o[16] = 1'b0;
  assign branch_metadata_fwd_o[17] = 1'b0;
  assign branch_metadata_fwd_o[18] = 1'b0;
  assign branch_metadata_fwd_o[19] = 1'b0;
  assign branch_metadata_fwd_o[20] = 1'b0;
  assign branch_metadata_fwd_o[21] = 1'b0;
  assign branch_metadata_fwd_o[35] = pc_fwd_i[8];
  assign branch_metadata_fwd_o[34] = pc_fwd_i[7];
  assign branch_metadata_fwd_o[33] = pc_fwd_i[6];
  assign branch_metadata_fwd_o[32] = pc_fwd_i[5];
  assign branch_metadata_fwd_o[26] = pc_fwd_i[4];
  assign branch_metadata_fwd_o[31] = pc_fwd_i[4];
  assign branch_metadata_fwd_o[25] = pc_fwd_i[3];
  assign branch_metadata_fwd_o[30] = pc_fwd_i[3];
  assign branch_metadata_fwd_o[24] = pc_fwd_i[2];
  assign branch_metadata_fwd_o[29] = pc_fwd_i[2];
  assign branch_metadata_fwd_o[23] = pc_fwd_i[1];
  assign branch_metadata_fwd_o[28] = pc_fwd_i[1];
  assign branch_metadata_fwd_o[22] = pc_fwd_i[0];
  assign branch_metadata_fwd_o[27] = pc_fwd_i[0];

  bp_fe_bht_bht_indx_width_p5
  bht_1
  (
    .clk_i(clk_i),
    .en_i(1'b1),
    .reset_i(reset_i),
    .idx_r_i(pc_fwd_i[4:0]),
    .idx_w_i(branch_metadata_fwd_i[26:22]),
    .r_v_i(r_v_i),
    .w_v_i(w_v_i),
    .correct_i(attaboy_i),
    .predict_o(predict)
  );


  bp_fe_btb_bp_fe_pc_gen_btb_idx_width_lp9_eaddr_width_p64
  btb_1
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .idx_w_i(branch_metadata_fwd_i[35:27]),
    .idx_r_i(pc_queue_i[8:0]),
    .r_v_i(r_v_i),
    .w_v_i(w_v_i),
    .branch_target_i(pc_cmd_i),
    .branch_target_o(pc_o),
    .read_valid_o(read_valid)
  );

  assign predict_o = predict & read_valid;

endmodule



module bp_fe_pc_gen_56_22_64_9_5_22_32_10_80000124_1
(
  clk_i,
  reset_i,
  v_i,
  pc_gen_icache_o,
  pc_gen_icache_v_o,
  pc_gen_icache_ready_i,
  icache_pc_gen_i,
  icache_pc_gen_v_i,
  icache_pc_gen_ready_o,
  icache_miss_i,
  pc_gen_itlb_o,
  pc_gen_itlb_v_o,
  pc_gen_itlb_ready_i,
  pc_gen_fe_o,
  pc_gen_fe_v_o,
  pc_gen_fe_ready_i,
  fe_pc_gen_i,
  fe_pc_gen_v_i,
  fe_pc_gen_ready_o
);

  output [63:0] pc_gen_icache_o;
  input [95:0] icache_pc_gen_i;
  output [63:0] pc_gen_itlb_o;
  output [202:0] pc_gen_fe_o;
  input [101:0] fe_pc_gen_i;
  input clk_i;
  input reset_i;
  input v_i;
  input pc_gen_icache_ready_i;
  input icache_pc_gen_v_i;
  input icache_miss_i;
  input pc_gen_itlb_ready_i;
  input pc_gen_fe_ready_i;
  input fe_pc_gen_v_i;
  output pc_gen_icache_v_o;
  output icache_pc_gen_ready_o;
  output pc_gen_itlb_v_o;
  output pc_gen_fe_v_o;
  output fe_pc_gen_ready_o;
  wire [63:0] pc_gen_itlb_o,next_pc,btb_target;
  wire [202:0] pc_gen_fe_o;
  wire pc_gen_icache_v_o,icache_pc_gen_ready_o,pc_gen_itlb_v_o,pc_gen_fe_v_o,
  fe_pc_gen_ready_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,misalignment,N12,
  pc_gen_exception_exception_code__1_,pc_gen_fetch_branch_metadata_fwd__35_,
  pc_gen_fetch_branch_metadata_fwd__34_,pc_gen_fetch_branch_metadata_fwd__33_,
  pc_gen_fetch_branch_metadata_fwd__32_,pc_gen_fetch_branch_metadata_fwd__31_,
  pc_gen_fetch_branch_metadata_fwd__30_,pc_gen_fetch_branch_metadata_fwd__29_,
  pc_gen_fetch_branch_metadata_fwd__28_,pc_gen_fetch_branch_metadata_fwd__27_,pc_gen_fetch_branch_metadata_fwd__26_,
  pc_gen_fetch_branch_metadata_fwd__25_,pc_gen_fetch_branch_metadata_fwd__24_,
  pc_gen_fetch_branch_metadata_fwd__23_,pc_gen_fetch_branch_metadata_fwd__22_,
  pc_gen_fetch_branch_metadata_fwd__21_,pc_gen_fetch_branch_metadata_fwd__20_,
  pc_gen_fetch_branch_metadata_fwd__19_,pc_gen_fetch_branch_metadata_fwd__18_,
  pc_gen_fetch_branch_metadata_fwd__17_,pc_gen_fetch_branch_metadata_fwd__16_,
  pc_gen_fetch_branch_metadata_fwd__15_,pc_gen_fetch_branch_metadata_fwd__14_,
  pc_gen_fetch_branch_metadata_fwd__13_,pc_gen_fetch_branch_metadata_fwd__12_,
  pc_gen_fetch_branch_metadata_fwd__11_,pc_gen_fetch_branch_metadata_fwd__10_,
  pc_gen_fetch_branch_metadata_fwd__9_,pc_gen_fetch_branch_metadata_fwd__8_,pc_gen_fetch_branch_metadata_fwd__7_,
  pc_gen_fetch_branch_metadata_fwd__6_,pc_gen_fetch_branch_metadata_fwd__5_,
  pc_gen_fetch_branch_metadata_fwd__4_,pc_gen_fetch_branch_metadata_fwd__3_,
  pc_gen_fetch_branch_metadata_fwd__2_,pc_gen_fetch_branch_metadata_fwd__1_,
  pc_gen_fetch_branch_metadata_fwd__0_,N13,N14,N15,N16,N17,predict,scan_instr_is_compressed_,
  scan_instr_instr_scan_class__3_,scan_instr_instr_scan_class__2_,
  scan_instr_instr_scan_class__1_,scan_instr_instr_scan_class__0_,scan_instr_imm__63_,scan_instr_imm__62_,
  scan_instr_imm__61_,scan_instr_imm__60_,scan_instr_imm__59_,scan_instr_imm__58_,
  scan_instr_imm__57_,scan_instr_imm__56_,scan_instr_imm__55_,scan_instr_imm__54_,
  scan_instr_imm__53_,scan_instr_imm__52_,scan_instr_imm__51_,scan_instr_imm__50_,
  scan_instr_imm__49_,scan_instr_imm__48_,scan_instr_imm__47_,scan_instr_imm__46_,
  scan_instr_imm__45_,scan_instr_imm__44_,scan_instr_imm__43_,scan_instr_imm__42_,
  scan_instr_imm__41_,scan_instr_imm__40_,scan_instr_imm__39_,scan_instr_imm__38_,
  scan_instr_imm__37_,scan_instr_imm__36_,scan_instr_imm__35_,scan_instr_imm__34_,
  scan_instr_imm__33_,scan_instr_imm__32_,scan_instr_imm__31_,scan_instr_imm__30_,
  scan_instr_imm__29_,scan_instr_imm__28_,scan_instr_imm__27_,scan_instr_imm__26_,
  scan_instr_imm__25_,scan_instr_imm__24_,scan_instr_imm__23_,scan_instr_imm__22_,
  scan_instr_imm__21_,scan_instr_imm__20_,scan_instr_imm__19_,scan_instr_imm__18_,
  scan_instr_imm__17_,scan_instr_imm__16_,scan_instr_imm__15_,scan_instr_imm__14_,
  scan_instr_imm__13_,scan_instr_imm__12_,scan_instr_imm__11_,scan_instr_imm__10_,
  scan_instr_imm__9_,scan_instr_imm__8_,scan_instr_imm__7_,scan_instr_imm__6_,
  scan_instr_imm__5_,scan_instr_imm__4_,scan_instr_imm__3_,scan_instr_imm__2_,
  scan_instr_imm__1_,scan_instr_imm__0_,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,
  N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,
  N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,
  N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,
  N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,
  N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,
  N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,
  N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,
  N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,
  N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,
  N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,
  N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,
  N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,
  N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,
  N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,
  N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,
  N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,
  N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,
  N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,
  N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,
  N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,
  N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,
  N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,
  N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,
  N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,
  N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,
  stalled_pc_redirect_n,N444,N445,N446,bht_r_v_branch_jalr_inst,N447,N448,N449,N450,
  N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,
  N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,
  N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,
  N499,N500,N501,N502,N503;
  reg [63:0] icache_miss_pc,pc_gen_icache_o,last_pc,pc_redirect;
  reg stalled_pc_redirect;
  assign pc_gen_fe_o[0] = 1'b0;
  assign pc_gen_itlb_v_o = 1'b0;
  assign icache_pc_gen_ready_o = 1'b0;
  assign pc_gen_itlb_o[63] = pc_gen_icache_o[63];
  assign pc_gen_itlb_o[62] = pc_gen_icache_o[62];
  assign pc_gen_itlb_o[61] = pc_gen_icache_o[61];
  assign pc_gen_itlb_o[60] = pc_gen_icache_o[60];
  assign pc_gen_itlb_o[59] = pc_gen_icache_o[59];
  assign pc_gen_itlb_o[58] = pc_gen_icache_o[58];
  assign pc_gen_itlb_o[57] = pc_gen_icache_o[57];
  assign pc_gen_itlb_o[56] = pc_gen_icache_o[56];
  assign pc_gen_itlb_o[55] = pc_gen_icache_o[55];
  assign pc_gen_itlb_o[54] = pc_gen_icache_o[54];
  assign pc_gen_itlb_o[53] = pc_gen_icache_o[53];
  assign pc_gen_itlb_o[52] = pc_gen_icache_o[52];
  assign pc_gen_itlb_o[51] = pc_gen_icache_o[51];
  assign pc_gen_itlb_o[50] = pc_gen_icache_o[50];
  assign pc_gen_itlb_o[49] = pc_gen_icache_o[49];
  assign pc_gen_itlb_o[48] = pc_gen_icache_o[48];
  assign pc_gen_itlb_o[47] = pc_gen_icache_o[47];
  assign pc_gen_itlb_o[46] = pc_gen_icache_o[46];
  assign pc_gen_itlb_o[45] = pc_gen_icache_o[45];
  assign pc_gen_itlb_o[44] = pc_gen_icache_o[44];
  assign pc_gen_itlb_o[43] = pc_gen_icache_o[43];
  assign pc_gen_itlb_o[42] = pc_gen_icache_o[42];
  assign pc_gen_itlb_o[41] = pc_gen_icache_o[41];
  assign pc_gen_itlb_o[40] = pc_gen_icache_o[40];
  assign pc_gen_itlb_o[39] = pc_gen_icache_o[39];
  assign pc_gen_itlb_o[38] = pc_gen_icache_o[38];
  assign pc_gen_itlb_o[37] = pc_gen_icache_o[37];
  assign pc_gen_itlb_o[36] = pc_gen_icache_o[36];
  assign pc_gen_itlb_o[35] = pc_gen_icache_o[35];
  assign pc_gen_itlb_o[34] = pc_gen_icache_o[34];
  assign pc_gen_itlb_o[33] = pc_gen_icache_o[33];
  assign pc_gen_itlb_o[32] = pc_gen_icache_o[32];
  assign pc_gen_itlb_o[31] = pc_gen_icache_o[31];
  assign pc_gen_itlb_o[30] = pc_gen_icache_o[30];
  assign pc_gen_itlb_o[29] = pc_gen_icache_o[29];
  assign pc_gen_itlb_o[28] = pc_gen_icache_o[28];
  assign pc_gen_itlb_o[27] = pc_gen_icache_o[27];
  assign pc_gen_itlb_o[26] = pc_gen_icache_o[26];
  assign pc_gen_itlb_o[25] = pc_gen_icache_o[25];
  assign pc_gen_itlb_o[24] = pc_gen_icache_o[24];
  assign pc_gen_itlb_o[23] = pc_gen_icache_o[23];
  assign pc_gen_itlb_o[22] = pc_gen_icache_o[22];
  assign pc_gen_itlb_o[21] = pc_gen_icache_o[21];
  assign pc_gen_itlb_o[20] = pc_gen_icache_o[20];
  assign pc_gen_itlb_o[19] = pc_gen_icache_o[19];
  assign pc_gen_itlb_o[18] = pc_gen_icache_o[18];
  assign pc_gen_itlb_o[17] = pc_gen_icache_o[17];
  assign pc_gen_itlb_o[16] = pc_gen_icache_o[16];
  assign pc_gen_itlb_o[15] = pc_gen_icache_o[15];
  assign pc_gen_itlb_o[14] = pc_gen_icache_o[14];
  assign pc_gen_itlb_o[13] = pc_gen_icache_o[13];
  assign pc_gen_itlb_o[12] = pc_gen_icache_o[12];
  assign pc_gen_itlb_o[11] = pc_gen_icache_o[11];
  assign pc_gen_itlb_o[10] = pc_gen_icache_o[10];
  assign pc_gen_itlb_o[9] = pc_gen_icache_o[9];
  assign pc_gen_itlb_o[8] = pc_gen_icache_o[8];
  assign pc_gen_itlb_o[7] = pc_gen_icache_o[7];
  assign pc_gen_itlb_o[6] = pc_gen_icache_o[6];
  assign pc_gen_itlb_o[5] = pc_gen_icache_o[5];
  assign pc_gen_itlb_o[4] = pc_gen_icache_o[4];
  assign pc_gen_itlb_o[3] = pc_gen_icache_o[3];
  assign pc_gen_itlb_o[2] = pc_gen_icache_o[2];
  assign pc_gen_itlb_o[1] = pc_gen_icache_o[1];
  assign pc_gen_itlb_o[0] = pc_gen_icache_o[0];
  assign N442 = icache_pc_gen_i[63:0] != pc_redirect;
  assign N443 = icache_pc_gen_i[63:0] == pc_redirect;

  instr_scan_eaddr_width_p64_instr_width_p32
  instr_scan_1
  (
    .instr_i(icache_pc_gen_i[95:64]),
    .scan_o({ scan_instr_is_compressed_, scan_instr_instr_scan_class__3_, scan_instr_instr_scan_class__2_, scan_instr_instr_scan_class__1_, scan_instr_instr_scan_class__0_, scan_instr_imm__63_, scan_instr_imm__62_, scan_instr_imm__61_, scan_instr_imm__60_, scan_instr_imm__59_, scan_instr_imm__58_, scan_instr_imm__57_, scan_instr_imm__56_, scan_instr_imm__55_, scan_instr_imm__54_, scan_instr_imm__53_, scan_instr_imm__52_, scan_instr_imm__51_, scan_instr_imm__50_, scan_instr_imm__49_, scan_instr_imm__48_, scan_instr_imm__47_, scan_instr_imm__46_, scan_instr_imm__45_, scan_instr_imm__44_, scan_instr_imm__43_, scan_instr_imm__42_, scan_instr_imm__41_, scan_instr_imm__40_, scan_instr_imm__39_, scan_instr_imm__38_, scan_instr_imm__37_, scan_instr_imm__36_, scan_instr_imm__35_, scan_instr_imm__34_, scan_instr_imm__33_, scan_instr_imm__32_, scan_instr_imm__31_, scan_instr_imm__30_, scan_instr_imm__29_, scan_instr_imm__28_, scan_instr_imm__27_, scan_instr_imm__26_, scan_instr_imm__25_, scan_instr_imm__24_, scan_instr_imm__23_, scan_instr_imm__22_, scan_instr_imm__21_, scan_instr_imm__20_, scan_instr_imm__19_, scan_instr_imm__18_, scan_instr_imm__17_, scan_instr_imm__16_, scan_instr_imm__15_, scan_instr_imm__14_, scan_instr_imm__13_, scan_instr_imm__12_, scan_instr_imm__11_, scan_instr_imm__10_, scan_instr_imm__9_, scan_instr_imm__8_, scan_instr_imm__7_, scan_instr_imm__6_, scan_instr_imm__5_, scan_instr_imm__4_, scan_instr_imm__3_, scan_instr_imm__2_, scan_instr_imm__1_, scan_instr_imm__0_ })
  );


  bp_fe_branch_predictor_eaddr_width_p64_btb_indx_width_p9_bht_indx_width_p5_ras_addr_width_p22
  genblk1_branch_prediction_1
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .attaboy_i(fe_pc_gen_i[0]),
    .r_v_i(bht_r_v_branch_jalr_inst),
    .w_v_i(fe_pc_gen_v_i),
    .pc_queue_i(last_pc),
    .pc_cmd_i(fe_pc_gen_i[101:38]),
    .pc_fwd_i(icache_pc_gen_i[63:0]),
    .branch_metadata_fwd_i(fe_pc_gen_i[37:2]),
    .predict_o(predict),
    .pc_o(btb_target),
    .branch_metadata_fwd_o({ pc_gen_fetch_branch_metadata_fwd__35_, pc_gen_fetch_branch_metadata_fwd__34_, pc_gen_fetch_branch_metadata_fwd__33_, pc_gen_fetch_branch_metadata_fwd__32_, pc_gen_fetch_branch_metadata_fwd__31_, pc_gen_fetch_branch_metadata_fwd__30_, pc_gen_fetch_branch_metadata_fwd__29_, pc_gen_fetch_branch_metadata_fwd__28_, pc_gen_fetch_branch_metadata_fwd__27_, pc_gen_fetch_branch_metadata_fwd__26_, pc_gen_fetch_branch_metadata_fwd__25_, pc_gen_fetch_branch_metadata_fwd__24_, pc_gen_fetch_branch_metadata_fwd__23_, pc_gen_fetch_branch_metadata_fwd__22_, pc_gen_fetch_branch_metadata_fwd__21_, pc_gen_fetch_branch_metadata_fwd__20_, pc_gen_fetch_branch_metadata_fwd__19_, pc_gen_fetch_branch_metadata_fwd__18_, pc_gen_fetch_branch_metadata_fwd__17_, pc_gen_fetch_branch_metadata_fwd__16_, pc_gen_fetch_branch_metadata_fwd__15_, pc_gen_fetch_branch_metadata_fwd__14_, pc_gen_fetch_branch_metadata_fwd__13_, pc_gen_fetch_branch_metadata_fwd__12_, pc_gen_fetch_branch_metadata_fwd__11_, pc_gen_fetch_branch_metadata_fwd__10_, pc_gen_fetch_branch_metadata_fwd__9_, pc_gen_fetch_branch_metadata_fwd__8_, pc_gen_fetch_branch_metadata_fwd__7_, pc_gen_fetch_branch_metadata_fwd__6_, pc_gen_fetch_branch_metadata_fwd__5_, pc_gen_fetch_branch_metadata_fwd__4_, pc_gen_fetch_branch_metadata_fwd__3_, pc_gen_fetch_branch_metadata_fwd__2_, pc_gen_fetch_branch_metadata_fwd__1_, pc_gen_fetch_branch_metadata_fwd__0_ })
  );

  assign N447 = ~scan_instr_instr_scan_class__0_;
  assign N448 = scan_instr_instr_scan_class__2_ | scan_instr_instr_scan_class__3_;
  assign N449 = scan_instr_instr_scan_class__1_ | N448;
  assign N450 = N447 | N449;
  assign N451 = ~N450;
  assign N452 = scan_instr_instr_scan_class__2_ | scan_instr_instr_scan_class__3_;
  assign N453 = scan_instr_instr_scan_class__1_ | N452;
  assign N454 = scan_instr_instr_scan_class__0_ | N453;
  assign N455 = ~N454;
  assign N456 = ~pc_gen_fe_o[202];
  assign N457 = N9 | N8;
  assign N458 = N10 | N457;
  assign N459 = N11 | N458;
  assign N460 = ~N459;
  assign N461 = ~N9;
  assign N462 = N461 | N8;
  assign N463 = N10 | N462;
  assign N464 = N11 | N463;
  assign N465 = ~N464;
  assign N466 = ~N8;
  assign N467 = N9 | N466;
  assign N468 = N10 | N467;
  assign N469 = N11 | N468;
  assign N470 = ~N469;
  assign N471 = N461 | N466;
  assign N472 = N10 | N471;
  assign N473 = N11 | N472;
  assign N474 = ~N473;
  assign N475 = ~scan_instr_instr_scan_class__1_;
  assign N476 = scan_instr_instr_scan_class__2_ | scan_instr_instr_scan_class__3_;
  assign N477 = N475 | N476;
  assign N478 = scan_instr_instr_scan_class__0_ | N477;
  assign N479 = ~N478;
  assign N480 = scan_instr_instr_scan_class__2_ | scan_instr_instr_scan_class__3_;
  assign N481 = scan_instr_instr_scan_class__1_ | N480;
  assign N482 = scan_instr_instr_scan_class__0_ | N481;
  assign N483 = ~N482;
  assign N484 = scan_instr_instr_scan_class__2_ | scan_instr_instr_scan_class__3_;
  assign N485 = scan_instr_instr_scan_class__1_ | N484;
  assign N486 = N447 | N485;
  assign N487 = ~N486;
  assign { N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156 } = pc_gen_icache_o + { 1'b1, 1'b0, 1'b0 };
  assign { N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27 } = icache_pc_gen_i[63:0] + { scan_instr_imm__63_, scan_instr_imm__62_, scan_instr_imm__61_, scan_instr_imm__60_, scan_instr_imm__59_, scan_instr_imm__58_, scan_instr_imm__57_, scan_instr_imm__56_, scan_instr_imm__55_, scan_instr_imm__54_, scan_instr_imm__53_, scan_instr_imm__52_, scan_instr_imm__51_, scan_instr_imm__50_, scan_instr_imm__49_, scan_instr_imm__48_, scan_instr_imm__47_, scan_instr_imm__46_, scan_instr_imm__45_, scan_instr_imm__44_, scan_instr_imm__43_, scan_instr_imm__42_, scan_instr_imm__41_, scan_instr_imm__40_, scan_instr_imm__39_, scan_instr_imm__38_, scan_instr_imm__37_, scan_instr_imm__36_, scan_instr_imm__35_, scan_instr_imm__34_, scan_instr_imm__33_, scan_instr_imm__32_, scan_instr_imm__31_, scan_instr_imm__30_, scan_instr_imm__29_, scan_instr_imm__28_, scan_instr_imm__27_, scan_instr_imm__26_, scan_instr_imm__25_, scan_instr_imm__24_, scan_instr_imm__23_, scan_instr_imm__22_, scan_instr_imm__21_, scan_instr_imm__20_, scan_instr_imm__19_, scan_instr_imm__18_, scan_instr_imm__17_, scan_instr_imm__16_, scan_instr_imm__15_, scan_instr_imm__14_, scan_instr_imm__13_, scan_instr_imm__12_, scan_instr_imm__11_, scan_instr_imm__10_, scan_instr_imm__9_, scan_instr_imm__8_, scan_instr_imm__7_, scan_instr_imm__6_, scan_instr_imm__5_, scan_instr_imm__4_, scan_instr_imm__3_, scan_instr_imm__2_, scan_instr_imm__1_, scan_instr_imm__0_ };
  assign { N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92 } = icache_pc_gen_i[63:0] + { scan_instr_imm__63_, scan_instr_imm__62_, scan_instr_imm__61_, scan_instr_imm__60_, scan_instr_imm__59_, scan_instr_imm__58_, scan_instr_imm__57_, scan_instr_imm__56_, scan_instr_imm__55_, scan_instr_imm__54_, scan_instr_imm__53_, scan_instr_imm__52_, scan_instr_imm__51_, scan_instr_imm__50_, scan_instr_imm__49_, scan_instr_imm__48_, scan_instr_imm__47_, scan_instr_imm__46_, scan_instr_imm__45_, scan_instr_imm__44_, scan_instr_imm__43_, scan_instr_imm__42_, scan_instr_imm__41_, scan_instr_imm__40_, scan_instr_imm__39_, scan_instr_imm__38_, scan_instr_imm__37_, scan_instr_imm__36_, scan_instr_imm__35_, scan_instr_imm__34_, scan_instr_imm__33_, scan_instr_imm__32_, scan_instr_imm__31_, scan_instr_imm__30_, scan_instr_imm__29_, scan_instr_imm__28_, scan_instr_imm__27_, scan_instr_imm__26_, scan_instr_imm__25_, scan_instr_imm__24_, scan_instr_imm__23_, scan_instr_imm__22_, scan_instr_imm__21_, scan_instr_imm__20_, scan_instr_imm__19_, scan_instr_imm__18_, scan_instr_imm__17_, scan_instr_imm__16_, scan_instr_imm__15_, scan_instr_imm__14_, scan_instr_imm__13_, scan_instr_imm__12_, scan_instr_imm__11_, scan_instr_imm__10_, scan_instr_imm__9_, scan_instr_imm__8_, scan_instr_imm__7_, scan_instr_imm__6_, scan_instr_imm__5_, scan_instr_imm__4_, scan_instr_imm__3_, scan_instr_imm__2_, scan_instr_imm__1_, scan_instr_imm__0_ };
  assign pc_gen_fe_o[132:1] = (N0)? { icache_pc_gen_i[63:0], icache_pc_gen_i[95:64], pc_gen_fetch_branch_metadata_fwd__35_, pc_gen_fetch_branch_metadata_fwd__34_, pc_gen_fetch_branch_metadata_fwd__33_, pc_gen_fetch_branch_metadata_fwd__32_, pc_gen_fetch_branch_metadata_fwd__31_, pc_gen_fetch_branch_metadata_fwd__30_, pc_gen_fetch_branch_metadata_fwd__29_, pc_gen_fetch_branch_metadata_fwd__28_, pc_gen_fetch_branch_metadata_fwd__27_, pc_gen_fetch_branch_metadata_fwd__26_, pc_gen_fetch_branch_metadata_fwd__25_, pc_gen_fetch_branch_metadata_fwd__24_, pc_gen_fetch_branch_metadata_fwd__23_, pc_gen_fetch_branch_metadata_fwd__22_, pc_gen_fetch_branch_metadata_fwd__21_, pc_gen_fetch_branch_metadata_fwd__20_, pc_gen_fetch_branch_metadata_fwd__19_, pc_gen_fetch_branch_metadata_fwd__18_, pc_gen_fetch_branch_metadata_fwd__17_, pc_gen_fetch_branch_metadata_fwd__16_, pc_gen_fetch_branch_metadata_fwd__15_, pc_gen_fetch_branch_metadata_fwd__14_, pc_gen_fetch_branch_metadata_fwd__13_, pc_gen_fetch_branch_metadata_fwd__12_, pc_gen_fetch_branch_metadata_fwd__11_, pc_gen_fetch_branch_metadata_fwd__10_, pc_gen_fetch_branch_metadata_fwd__9_, pc_gen_fetch_branch_metadata_fwd__8_, pc_gen_fetch_branch_metadata_fwd__7_, pc_gen_fetch_branch_metadata_fwd__6_, pc_gen_fetch_branch_metadata_fwd__5_, pc_gen_fetch_branch_metadata_fwd__4_, pc_gen_fetch_branch_metadata_fwd__3_, pc_gen_fetch_branch_metadata_fwd__2_, pc_gen_fetch_branch_metadata_fwd__1_, pc_gen_fetch_branch_metadata_fwd__0_ } : 
                              (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, pc_gen_exception_exception_code__1_, pc_gen_exception_exception_code__1_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N456;
  assign N1 = pc_gen_fe_o[202];
  assign pc_gen_fe_v_o = (N2)? 1'b0 : 
                         (N3)? N15 : 1'b0;
  assign N2 = N14;
  assign N3 = N13;
  assign fe_pc_gen_ready_o = (N2)? 1'b0 : 
                             (N3)? fe_pc_gen_v_i : 1'b0;
  assign pc_gen_icache_v_o = (N2)? 1'b0 : 
                             (N3)? N16 : 1'b0;
  assign next_pc = (N4)? icache_miss_pc : 
                   (N221)? fe_pc_gen_i[101:38] : 
                   (N224)? btb_target : 
                   (N227)? { N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27 } : 
                   (N230)? { N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92 } : 
                   (N25)? { N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156 } : 1'b0;
  assign N4 = icache_miss_i;
  assign { N241, N239 } = (N5)? { 1'b1, 1'b1 } : 
                          (N434)? { 1'b1, 1'b1 } : 
                          (N437)? { 1'b1, 1'b1 } : 
                          (N440)? { 1'b1, 1'b1 } : 
                          (N238)? { 1'b0, 1'b0 } : 1'b0;
  assign N5 = N234;
  assign { N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N240 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N434)? pc_redirect : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N437)? next_pc : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N440)? icache_miss_pc : 1'b0;
  assign { N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N434)? pc_gen_icache_o : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N437)? pc_gen_icache_o : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N440)? pc_gen_icache_o : 1'b0;
  assign { N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N434)? last_pc : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N437)? last_pc : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N440)? last_pc : 1'b0;
  assign N446 = (N6)? 1'b0 : 
                (N7)? stalled_pc_redirect_n : 1'b0;
  assign N6 = N445;
  assign N7 = N444;
  assign N8 = ~fe_pc_gen_i[41];
  assign N9 = ~fe_pc_gen_i[40];
  assign N10 = ~fe_pc_gen_i[39];
  assign N11 = ~fe_pc_gen_i[38];
  assign misalignment = N491 & N474;
  assign N491 = N490 & N470;
  assign N490 = N489 & N465;
  assign N489 = N488 & N460;
  assign N488 = fe_pc_gen_v_i & fe_pc_gen_i[1];
  assign pc_gen_fe_o[202] = misalignment;
  assign N12 = ~misalignment;
  assign pc_gen_exception_exception_code__1_ = N12;
  assign N13 = ~reset_i;
  assign N14 = reset_i;
  assign N15 = N492 & N493;
  assign N492 = pc_gen_fe_ready_i & icache_pc_gen_v_i;
  assign N493 = ~icache_miss_i;
  assign N16 = pc_gen_fe_ready_i & N493;
  assign N17 = fe_pc_gen_i[1] & fe_pc_gen_v_i;
  assign N18 = N494 & N487;
  assign N494 = predict & icache_pc_gen_v_i;
  assign N19 = N495 & N483;
  assign N495 = predict & icache_pc_gen_v_i;
  assign N20 = icache_pc_gen_v_i & N479;
  assign N21 = N17 | icache_miss_i;
  assign N22 = N18 | N21;
  assign N23 = N19 | N22;
  assign N24 = N20 | N23;
  assign N25 = ~N24;
  assign N26 = N227;
  assign N91 = N230;
  assign N220 = ~icache_miss_i;
  assign N221 = N17 & N220;
  assign N222 = ~N17;
  assign N223 = N220 & N222;
  assign N224 = N18 & N223;
  assign N225 = ~N18;
  assign N226 = N223 & N225;
  assign N227 = N19 & N226;
  assign N228 = ~N19;
  assign N229 = N226 & N228;
  assign N230 = N20 & N229;
  assign N231 = stalled_pc_redirect & icache_miss_i;
  assign N232 = pc_gen_icache_ready_i & pc_gen_fe_ready_i;
  assign N233 = icache_miss_i & N496;
  assign N496 = ~pc_gen_icache_ready_i;
  assign N234 = reset_i;
  assign N235 = N231 | N234;
  assign N236 = N232 | N235;
  assign N237 = N233 | N236;
  assign N238 = ~N237;
  assign N433 = ~N234;
  assign N434 = N231 & N433;
  assign N435 = ~N231;
  assign N436 = N433 & N435;
  assign N437 = N232 & N436;
  assign N438 = ~N232;
  assign N439 = N436 & N438;
  assign N440 = N233 & N439;
  assign N441 = fe_pc_gen_v_i & fe_pc_gen_i[1];
  assign stalled_pc_redirect_n = N499 | N502;
  assign N499 = N497 | N498;
  assign N497 = fe_pc_gen_v_i & fe_pc_gen_i[1];
  assign N498 = stalled_pc_redirect & N442;
  assign N502 = N500 & N501;
  assign N500 = stalled_pc_redirect & N443;
  assign N501 = ~pc_gen_fe_v_o;
  assign N444 = ~reset_i;
  assign N445 = reset_i;
  assign bht_r_v_branch_jalr_inst = icache_pc_gen_v_i & N503;
  assign N503 = N451 | N455;

  always @(posedge clk_i) begin
    if(N239) begin
      { icache_miss_pc[63:0] } <= { N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369 };
      { pc_gen_icache_o[0:0] } <= { N240 };
      { last_pc[63:29] } <= { N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334 };
    end 
    if(N241) begin
      { pc_gen_icache_o[63:1] } <= { N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242 };
      { last_pc[28:0] } <= { N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305 };
    end 
    if(N441) begin
      { pc_redirect[63:0] } <= { fe_pc_gen_i[101:38] };
    end 
    if(1'b1) begin
      stalled_pc_redirect <= N446;
    end 
  end


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p96_els_p64
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [95:0] data_i;
  input [5:0] addr_i;
  input [95:0] w_mask_i;
  output [95:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [95:0] data_o;

  hard_mem_1rw_bit_mask_d64_w96_wrapper
  macro_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  addr_i,
  data_i,
  write_mask_i,
  data_o
);

  input [8:0] addr_i;
  input [63:0] data_i;
  input [7:0] write_mask_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [63:0] data_o;

  hard_mem_1rw_byte_mask_d512_w64_wrapper
  macro_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .w_i(w_i),
    .addr_i(addr_i),
    .data_i(data_i),
    .write_mask_i(write_mask_i),
    .data_o(data_o)
  );


endmodule



module bsg_scan_width_p8_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [7:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__7_,t_1__6_,
  t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__7_ = i[0] | 1'b0;
  assign t_1__6_ = i[1] | i[0];
  assign t_1__5_ = i[2] | i[1];
  assign t_1__4_ = i[3] | i[2];
  assign t_1__3_ = i[4] | i[3];
  assign t_1__2_ = i[5] | i[4];
  assign t_1__1_ = i[6] | i[5];
  assign t_1__0_ = i[7] | i[6];
  assign t_2__7_ = t_1__7_ | 1'b0;
  assign t_2__6_ = t_1__6_ | 1'b0;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign o[0] = t_2__7_ | 1'b0;
  assign o[1] = t_2__6_ | 1'b0;
  assign o[2] = t_2__5_ | 1'b0;
  assign o[3] = t_2__4_ | 1'b0;
  assign o[4] = t_2__3_ | t_2__7_;
  assign o[5] = t_2__2_ | t_2__6_;
  assign o[6] = t_2__1_ | t_2__5_;
  assign o[7] = t_2__0_ | t_2__4_;

endmodule



module bsg_priority_encode_one_hot_out_width_p8_lo_to_hi_p1
(
  i,
  o
);

  input [7:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire N0,N1,N2,N3,N4,N5,N6;
  wire [7:1] scan_lo;

  bsg_scan_width_p8_or_p1_lo_to_hi_p1
  scan
  (
    .i(i),
    .o({ scan_lo, o[0:0] })
  );

  assign o[7] = scan_lo[7] & N0;
  assign N0 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N1;
  assign N1 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N2;
  assign N2 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N3;
  assign N3 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N4;
  assign N4 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N5;
  assign N5 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N6;
  assign N6 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p1
(
  i,
  addr_o,
  v_o
);

  input [0:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign v_o = i[0];
  assign addr_o[0] = 1'b0;

endmodule



module bsg_encode_one_hot_width_p2
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o,aligned_vs;
  wire v_o;
  wire [1:0] aligned_addrs;

  bsg_encode_one_hot_width_p1
  aligned_left
  (
    .i(i[0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p1
  aligned_right
  (
    .i(i[1]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[0])
  );

  assign v_o = addr_o[0] | aligned_vs[0];

endmodule



module bsg_encode_one_hot_width_p4
(
  i,
  addr_o,
  v_o
);

  input [3:0] i;
  output [1:0] addr_o;
  output v_o;
  wire [1:0] addr_o,aligned_addrs;
  wire v_o;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p2
  aligned_left
  (
    .i(i[1:0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p2
  aligned_right
  (
    .i(i[3:2]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[1])
  );

  assign v_o = addr_o[1] | aligned_vs[0];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[1];

endmodule



module bsg_encode_one_hot_width_p8_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [3:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p4
  aligned_left
  (
    .i(i[3:0]),
    .addr_o(aligned_addrs[1:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p4
  aligned_right
  (
    .i(i[7:4]),
    .addr_o(aligned_addrs[3:2]),
    .v_o(addr_o[2])
  );

  assign v_o = addr_o[2] | aligned_vs[0];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[3];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[2];

endmodule



module bsg_priority_encode_width_p8_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [7:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p8_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo)
  );


  bsg_encode_one_hot_width_p8_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o),
    .v_o(v_o)
  );


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p7_els_p64
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [6:0] data_i;
  input [5:0] addr_i;
  input [6:0] w_mask_i;
  output [6:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [6:0] data_o;

  hard_mem_1rw_bit_mask_d64_w7_wrapper
  macro_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bp_be_dcache_lru_encode_ways_p8
(
  lru_i,
  way_id_o
);

  input [6:0] lru_i;
  output [2:0] way_id_o;
  wire [2:0] way_id_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30;
  assign N11 = N8 & N9;
  assign N12 = N11 & N10;
  assign N13 = lru_i[3] & N9;
  assign N14 = N13 & N10;
  assign N16 = N15 & lru_i[1];
  assign N17 = N16 & N10;
  assign N18 = lru_i[4] & lru_i[1];
  assign N19 = N18 & N10;
  assign N22 = N20 & N21;
  assign N23 = N22 & lru_i[0];
  assign N24 = lru_i[5] & N21;
  assign N25 = N24 & lru_i[0];
  assign N27 = N26 & lru_i[2];
  assign N28 = N27 & lru_i[0];
  assign N29 = lru_i[6] & lru_i[2];
  assign N30 = N29 & lru_i[0];
  assign way_id_o = (N0)? { 1'b0, 1'b0, 1'b0 } : 
                    (N1)? { 1'b0, 1'b0, 1'b1 } : 
                    (N2)? { 1'b0, 1'b1, 1'b0 } : 
                    (N3)? { 1'b0, 1'b1, 1'b1 } : 
                    (N4)? { 1'b1, 1'b0, 1'b0 } : 
                    (N5)? { 1'b1, 1'b0, 1'b1 } : 
                    (N6)? { 1'b1, 1'b1, 1'b0 } : 
                    (N7)? { 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N0 = N12;
  assign N1 = N14;
  assign N2 = N17;
  assign N3 = N19;
  assign N4 = N23;
  assign N5 = N25;
  assign N6 = N28;
  assign N7 = N30;
  assign N8 = ~lru_i[3];
  assign N9 = ~lru_i[1];
  assign N10 = ~lru_i[0];
  assign N15 = ~lru_i[4];
  assign N20 = ~lru_i[5];
  assign N21 = ~lru_i[2];
  assign N26 = ~lru_i[6];

endmodule



module bp_fe_lce_req_data_width_p64_lce_addr_width_p22_num_cce_p1_num_lce_p2_lce_sets_p64_ways_p8_block_size_in_bytes_p8
(
  clk_i,
  reset_i,
  id_i,
  miss_i,
  miss_addr_i,
  lru_way_i,
  cache_miss_o,
  tr_received_i,
  cce_data_received_i,
  tag_set_i,
  tag_set_wakeup_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_yumi_i
);

  input [0:0] id_i;
  input [21:0] miss_addr_i;
  input [2:0] lru_way_i;
  output [29:0] lce_req_o;
  output [25:0] lce_resp_o;
  input clk_i;
  input reset_i;
  input miss_i;
  input tr_received_i;
  input cce_data_received_i;
  input tag_set_i;
  input tag_set_wakeup_i;
  input lce_req_ready_i;
  input lce_resp_yumi_i;
  output cache_miss_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  wire cache_miss_o,lce_req_v_o,lce_resp_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,tr_received_n,
  cce_data_received_n,tag_set_n,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,
  N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112;
  wire [2:0] state_n,lru_way_n;
  wire [21:0] miss_addr_n;
  reg [25:0] lce_resp_o;
  reg [29:0] lce_req_o;
  reg [2:0] state_r;
  reg tr_received_r,cce_data_received_r,tag_set_r;
  assign lce_resp_o[23] = 1'b1;
  assign lce_req_o[29] = lce_resp_o[25];
  assign lce_req_o[25] = lce_resp_o[21];
  assign lce_req_o[24] = lce_resp_o[20];
  assign lce_req_o[23] = lce_resp_o[19];
  assign lce_req_o[22] = lce_resp_o[18];
  assign lce_req_o[21] = lce_resp_o[17];
  assign lce_req_o[20] = lce_resp_o[16];
  assign lce_req_o[19] = lce_resp_o[15];
  assign lce_req_o[18] = lce_resp_o[14];
  assign lce_req_o[17] = lce_resp_o[13];
  assign lce_req_o[16] = lce_resp_o[12];
  assign lce_req_o[15] = lce_resp_o[11];
  assign lce_req_o[14] = lce_resp_o[10];
  assign lce_req_o[13] = lce_resp_o[9];
  assign lce_req_o[12] = lce_resp_o[8];
  assign lce_req_o[11] = lce_resp_o[7];
  assign lce_req_o[10] = lce_resp_o[6];
  assign lce_req_o[9] = lce_resp_o[5];
  assign lce_req_o[8] = lce_resp_o[4];
  assign lce_req_o[7] = lce_resp_o[3];
  assign lce_req_o[6] = lce_resp_o[2];
  assign lce_req_o[5] = lce_resp_o[1];
  assign lce_req_o[4] = lce_resp_o[0];
  assign lce_req_o[0] = 1'b0;
  assign lce_req_o[26] = 1'b0;
  assign lce_req_o[27] = 1'b0;
  assign lce_req_o[28] = id_i[0];
  assign lce_resp_o[24] = id_i[0];
  assign N15 = N12 & N13;
  assign N16 = N15 & N14;
  assign N17 = state_r[2] | state_r[1];
  assign N18 = N17 | N14;
  assign N20 = N12 | state_r[1];
  assign N21 = N20 | state_r[0];
  assign N23 = state_r[2] | N13;
  assign N24 = N23 | state_r[0];
  assign N26 = state_r[2] | N13;
  assign N27 = N26 | N14;
  assign { N40, N39, N38 } = (N0)? { 1'b0, 1'b1, 1'b0 } : 
                             (N53)? { 1'b0, 1'b1, 1'b1 } : 
                             (N37)? { 1'b1, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N9;
  assign { N43, N42, N41 } = (N1)? { 1'b0, 1'b0, 1'b0 } : 
                             (N51)? { N40, N39, N38 } : 
                             (N35)? { 1'b1, 1'b0, 1'b0 } : 1'b0;
  assign N1 = tag_set_wakeup_i;
  assign cache_miss_o = (N2)? miss_i : 
                        (N3)? 1'b1 : 
                        (N4)? 1'b1 : 
                        (N5)? 1'b1 : 
                        (N6)? 1'b1 : 
                        (N49)? 1'b0 : 1'b0;
  assign N2 = N16;
  assign N3 = N19;
  assign N4 = N22;
  assign N5 = N25;
  assign N6 = N28;
  assign state_n = (N2)? { 1'b0, 1'b0, 1'b1 } : 
                   (N3)? { lce_req_ready_i, 1'b0, N30 } : 
                   (N4)? { N43, N42, N41 } : 
                   (N5)? { 1'b0, N44, 1'b0 } : 
                   (N6)? { 1'b0, N44, N44 } : 
                   (N49)? state_r : 1'b0;
  assign miss_addr_n = (N2)? miss_addr_i : 
                       (N49)? lce_resp_o[21:0] : 1'b0;
  assign lru_way_n = (N2)? lru_way_i : 
                     (N49)? lce_req_o[3:1] : 1'b0;
  assign tr_received_n = (N2)? 1'b0 : 
                         (N4)? 1'b1 : 
                         (N49)? tr_received_r : 1'b0;
  assign cce_data_received_n = (N2)? 1'b0 : 
                               (N4)? 1'b1 : 
                               (N49)? cce_data_received_r : 1'b0;
  assign tag_set_n = (N2)? 1'b0 : 
                     (N4)? 1'b1 : 
                     (N49)? tag_set_r : 1'b0;
  assign lce_req_v_o = (N2)? 1'b0 : 
                       (N3)? 1'b1 : 
                       (N4)? 1'b0 : 
                       (N5)? 1'b0 : 
                       (N6)? 1'b0 : 
                       (N49)? 1'b0 : 1'b0;
  assign lce_resp_v_o = (N2)? 1'b0 : 
                        (N3)? 1'b0 : 
                        (N4)? 1'b0 : 
                        (N5)? 1'b1 : 
                        (N6)? 1'b1 : 
                        (N49)? 1'b0 : 1'b0;
  assign lce_resp_o[22] = (N2)? 1'b0 : 
                          (N3)? 1'b0 : 
                          (N4)? 1'b0 : 
                          (N5)? 1'b0 : 
                          (N6)? 1'b1 : 
                          (N49)? 1'b0 : 1'b0;
  assign { N57, N56, N55 } = (N7)? { 1'b0, 1'b0, 1'b0 } : 
                             (N8)? state_n : 1'b0;
  assign N7 = reset_i;
  assign N8 = N54;
  assign { N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58 } = (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                            (N8)? miss_addr_n : 1'b0;
  assign N80 = (N7)? 1'b0 : 
               (N8)? tr_received_n : 1'b0;
  assign N81 = (N7)? 1'b0 : 
               (N8)? cce_data_received_n : 1'b0;
  assign N82 = (N7)? 1'b0 : 
               (N8)? tag_set_n : 1'b0;
  assign { N85, N84, N83 } = (N7)? { 1'b0, 1'b0, 1'b0 } : 
                             (N8)? lru_way_n : 1'b0;
  assign N9 = tr_received_r | tr_received_i;
  assign N10 = cce_data_received_r | cce_data_received_i;
  assign N11 = tag_set_r | tag_set_i;
  assign N12 = ~state_r[2];
  assign N13 = ~state_r[1];
  assign N14 = ~state_r[0];
  assign N19 = ~N18;
  assign N22 = ~N21;
  assign N25 = ~N24;
  assign N28 = ~N27;
  assign N29 = ~miss_i;
  assign N30 = ~lce_req_ready_i;
  assign N31 = ~tr_received_i;
  assign N32 = ~cce_data_received_i;
  assign N33 = ~tag_set_i;
  assign N34 = N11 | tag_set_wakeup_i;
  assign N35 = ~N34;
  assign N36 = N10 | N9;
  assign N37 = ~N36;
  assign N44 = ~lce_resp_yumi_i;
  assign N45 = N19 | N16;
  assign N46 = N22 | N45;
  assign N47 = N25 | N46;
  assign N48 = N28 | N47;
  assign N49 = ~N48;
  assign N50 = ~tag_set_wakeup_i;
  assign N51 = N11 & N50;
  assign N52 = ~N9;
  assign N53 = N10 & N52;
  assign N54 = ~reset_i;
  assign N86 = N16 & N54;
  assign N87 = N29 & N86;
  assign N88 = N19 & N54;
  assign N89 = N87 | N88;
  assign N90 = N22 & N54;
  assign N91 = N89 | N90;
  assign N92 = N25 & N54;
  assign N93 = N91 | N92;
  assign N94 = N28 & N54;
  assign N95 = N93 | N94;
  assign N96 = ~N95;
  assign N97 = ~N87;
  assign N98 = N31 & N90;
  assign N99 = N89 | N98;
  assign N100 = N99 | N92;
  assign N101 = N100 | N94;
  assign N102 = ~N101;
  assign N103 = N32 & N90;
  assign N104 = N89 | N103;
  assign N105 = N104 | N92;
  assign N106 = N105 | N94;
  assign N107 = ~N106;
  assign N108 = N33 & N90;
  assign N109 = N89 | N108;
  assign N110 = N109 | N92;
  assign N111 = N110 | N94;
  assign N112 = ~N111;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { lce_resp_o[25:25] } <= { 1'b0 };
    end 
    if(N96) begin
      { lce_req_o[3:1] } <= { N85, N84, N83 };
      { lce_resp_o[21:0] } <= { N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58 };
    end 
    if(N97) begin
      { state_r[2:0] } <= { N57, N56, N55 };
    end 
    if(N102) begin
      tr_received_r <= N80;
    end 
    if(N107) begin
      cce_data_received_r <= N81;
    end 
    if(N112) begin
      tag_set_r <= N82;
    end 
  end


endmodule



// module bsg_mem_p36
// (
//   w_clk_i,
//   w_reset_i,
//   w_v_i,
//   w_addr_i,
//   w_data_i,
//   r_v_i,
//   r_addr_i,
//   r_data_o
// );

//   input [0:0] w_addr_i;
//   input [35:0] w_data_i;
//   input [0:0] r_addr_i;
//   output [35:0] r_data_o;
//   input w_clk_i;
//   input w_reset_i;
//   input w_v_i;
//   input r_v_i;
//   wire [35:0] r_data_o;
//   wire N0,N1,N2,N3,N4,N5,N7,N8;
//   reg [71:0] mem;
//   assign r_data_o[35] = (N3)? mem[35] : 
//                         (N0)? mem[71] : 1'b0;
//   assign N0 = r_addr_i[0];
//   assign r_data_o[34] = (N3)? mem[34] : 
//                         (N0)? mem[70] : 1'b0;
//   assign r_data_o[33] = (N3)? mem[33] : 
//                         (N0)? mem[69] : 1'b0;
//   assign r_data_o[32] = (N3)? mem[32] : 
//                         (N0)? mem[68] : 1'b0;
//   assign r_data_o[31] = (N3)? mem[31] : 
//                         (N0)? mem[67] : 1'b0;
//   assign r_data_o[30] = (N3)? mem[30] : 
//                         (N0)? mem[66] : 1'b0;
//   assign r_data_o[29] = (N3)? mem[29] : 
//                         (N0)? mem[65] : 1'b0;
//   assign r_data_o[28] = (N3)? mem[28] : 
//                         (N0)? mem[64] : 1'b0;
//   assign r_data_o[27] = (N3)? mem[27] : 
//                         (N0)? mem[63] : 1'b0;
//   assign r_data_o[26] = (N3)? mem[26] : 
//                         (N0)? mem[62] : 1'b0;
//   assign r_data_o[25] = (N3)? mem[25] : 
//                         (N0)? mem[61] : 1'b0;
//   assign r_data_o[24] = (N3)? mem[24] : 
//                         (N0)? mem[60] : 1'b0;
//   assign r_data_o[23] = (N3)? mem[23] : 
//                         (N0)? mem[59] : 1'b0;
//   assign r_data_o[22] = (N3)? mem[22] : 
//                         (N0)? mem[58] : 1'b0;
//   assign r_data_o[21] = (N3)? mem[21] : 
//                         (N0)? mem[57] : 1'b0;
//   assign r_data_o[20] = (N3)? mem[20] : 
//                         (N0)? mem[56] : 1'b0;
//   assign r_data_o[19] = (N3)? mem[19] : 
//                         (N0)? mem[55] : 1'b0;
//   assign r_data_o[18] = (N3)? mem[18] : 
//                         (N0)? mem[54] : 1'b0;
//   assign r_data_o[17] = (N3)? mem[17] : 
//                         (N0)? mem[53] : 1'b0;
//   assign r_data_o[16] = (N3)? mem[16] : 
//                         (N0)? mem[52] : 1'b0;
//   assign r_data_o[15] = (N3)? mem[15] : 
//                         (N0)? mem[51] : 1'b0;
//   assign r_data_o[14] = (N3)? mem[14] : 
//                         (N0)? mem[50] : 1'b0;
//   assign r_data_o[13] = (N3)? mem[13] : 
//                         (N0)? mem[49] : 1'b0;
//   assign r_data_o[12] = (N3)? mem[12] : 
//                         (N0)? mem[48] : 1'b0;
//   assign r_data_o[11] = (N3)? mem[11] : 
//                         (N0)? mem[47] : 1'b0;
//   assign r_data_o[10] = (N3)? mem[10] : 
//                         (N0)? mem[46] : 1'b0;
//   assign r_data_o[9] = (N3)? mem[9] : 
//                        (N0)? mem[45] : 1'b0;
//   assign r_data_o[8] = (N3)? mem[8] : 
//                        (N0)? mem[44] : 1'b0;
//   assign r_data_o[7] = (N3)? mem[7] : 
//                        (N0)? mem[43] : 1'b0;
//   assign r_data_o[6] = (N3)? mem[6] : 
//                        (N0)? mem[42] : 1'b0;
//   assign r_data_o[5] = (N3)? mem[5] : 
//                        (N0)? mem[41] : 1'b0;
//   assign r_data_o[4] = (N3)? mem[4] : 
//                        (N0)? mem[40] : 1'b0;
//   assign r_data_o[3] = (N3)? mem[3] : 
//                        (N0)? mem[39] : 1'b0;
//   assign r_data_o[2] = (N3)? mem[2] : 
//                        (N0)? mem[38] : 1'b0;
//   assign r_data_o[1] = (N3)? mem[1] : 
//                        (N0)? mem[37] : 1'b0;
//   assign r_data_o[0] = (N3)? mem[0] : 
//                        (N0)? mem[36] : 1'b0;
//   assign N5 = ~w_addr_i[0];
//   assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
//                       (N2)? { 1'b0, 1'b0 } : 1'b0;
//   assign N1 = w_v_i;
//   assign N2 = N4;
//   assign N3 = ~r_addr_i[0];
//   assign N4 = ~w_v_i;

//   always @(posedge w_clk_i) begin
//     if(N8) begin
//       { mem[71:36] } <= { w_data_i[35:0] };
//     end 
//     if(N7) begin
//       { mem[35:0] } <= { w_data_i[35:0] };
//     end 
//   end


// endmodule



module bsg_mem_1r1w_width_p36_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [35:0] w_data_i;
  input [0:0] r_addr_i;
  output [35:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [35:0] r_data_o;

  bsg_mem_p36
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p36
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [35:0] data_i;
  output [35:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [35:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p36_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 : 
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 : 
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 : 
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 : 
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 : 
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 : 
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end 
    if(N9) begin
      tail_r <= N10;
    end 
    if(N11) begin
      head_r <= N12;
    end 
  end


endmodule



module bp_fe_lce_cmd_data_width_p64_lce_data_width_p512_lce_addr_width_p22_lce_sets_p64_ways_p8_tag_width_p10_num_cce_p1_num_lce_p2_block_size_in_bytes_p8
(
  clk_i,
  reset_i,
  id_i,
  lce_ready_o,
  tag_set_o,
  tag_set_wakeup_o,
  data_mem_data_i,
  data_mem_pkt_o,
  data_mem_pkt_v_o,
  data_mem_pkt_yumi_i,
  tag_mem_pkt_o,
  tag_mem_pkt_v_o,
  tag_mem_pkt_yumi_i,
  metadata_mem_pkt_v_o,
  metadata_mem_pkt_o,
  metadata_mem_pkt_yumi_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_yumi_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_yumi_o,
  lce_tr_resp_o,
  lce_tr_resp_v_o,
  lce_tr_resp_ready_i
);

  input [0:0] id_i;
  input [511:0] data_mem_data_i;
  output [521:0] data_mem_pkt_o;
  output [22:0] tag_mem_pkt_o;
  output [9:0] metadata_mem_pkt_o;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  input [35:0] lce_cmd_i;
  output [538:0] lce_tr_resp_o;
  input clk_i;
  input reset_i;
  input data_mem_pkt_yumi_i;
  input tag_mem_pkt_yumi_i;
  input metadata_mem_pkt_yumi_i;
  input lce_resp_yumi_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_tr_resp_ready_i;
  output lce_ready_o;
  output tag_set_o;
  output tag_set_wakeup_o;
  output data_mem_pkt_v_o;
  output tag_mem_pkt_v_o;
  output metadata_mem_pkt_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_yumi_o;
  output lce_tr_resp_v_o;
  wire [521:0] data_mem_pkt_o;
  wire [22:0] tag_mem_pkt_o;
  wire [9:0] metadata_mem_pkt_o;
  wire [25:0] lce_resp_o;
  wire [536:0] lce_data_resp_o;
  wire [538:0] lce_tr_resp_o;
  wire lce_ready_o,tag_set_o,tag_set_wakeup_o,data_mem_pkt_v_o,tag_mem_pkt_v_o,
  metadata_mem_pkt_v_o,lce_resp_v_o,lce_data_resp_v_o,lce_cmd_yumi_o,lce_tr_resp_v_o,N0,
  N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,
  N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,
  N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,
  N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,
  N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,
  N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,
  N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,
  N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,
  N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,
  N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,
  N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,
  N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,
  N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,
  N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,
  N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,
  N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,
  N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,
  N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,
  N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,
  N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,
  N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,
  N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,
  N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,
  N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,
  N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,
  N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,
  N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,
  N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,
  N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,
  N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,
  N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,
  N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,
  N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,
  N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,
  N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,
  N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,
  N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,
  N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,
  N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,
  N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,
  N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,
  N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,
  N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,
  N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,
  N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
  N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,
  N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,N774,
  N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,N790,
  N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,N806,
  N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,N822,
  N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,N838,
  N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,N854,
  N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,N870,
  N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,N886,
  N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,N902,
  N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,N918,
  N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,N934,
  N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,N950,
  N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,N966,
  N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,N982,
  N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,N998,
  N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1011,
  N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038,
  N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,N1051,
  N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,
  N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091,
  N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118,
  N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,N1131,
  N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,
  N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,N1171,
  N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,N1198,
  N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,N1211,
  N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,N1238,
  N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,N1251,
  N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,N1278,
  N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,N1291,
  N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,
  N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,N1318,
  N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,N1331,
  N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,
  N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,N1358,
  N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,N1371,
  N1372,N1373,N1374,N1375,N1376,N1378,N1379,N1380,N1381,N1382,N1383,N1384,N1385,
  N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,
  N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407;
  wire [1:0] state_n;
  reg flag_updated_lru_r,flag_data_buffered_r,flag_invalidate_r;
  reg [1:0] state_r;
  reg [5:0] syn_ack_cnt_r;
  reg [511:0] data_r;
  assign data_mem_pkt_o[0] = 1'b0;
  assign data_mem_pkt_o[1] = 1'b0;
  assign data_mem_pkt_o[2] = 1'b0;
  assign data_mem_pkt_o[3] = 1'b0;
  assign data_mem_pkt_o[4] = 1'b0;
  assign data_mem_pkt_o[5] = 1'b0;
  assign data_mem_pkt_o[6] = 1'b0;
  assign data_mem_pkt_o[7] = 1'b0;
  assign data_mem_pkt_o[8] = 1'b0;
  assign data_mem_pkt_o[9] = 1'b0;
  assign data_mem_pkt_o[10] = 1'b0;
  assign data_mem_pkt_o[11] = 1'b0;
  assign data_mem_pkt_o[12] = 1'b0;
  assign data_mem_pkt_o[13] = 1'b0;
  assign data_mem_pkt_o[14] = 1'b0;
  assign data_mem_pkt_o[15] = 1'b0;
  assign data_mem_pkt_o[16] = 1'b0;
  assign data_mem_pkt_o[17] = 1'b0;
  assign data_mem_pkt_o[18] = 1'b0;
  assign data_mem_pkt_o[19] = 1'b0;
  assign data_mem_pkt_o[20] = 1'b0;
  assign data_mem_pkt_o[21] = 1'b0;
  assign data_mem_pkt_o[22] = 1'b0;
  assign data_mem_pkt_o[23] = 1'b0;
  assign data_mem_pkt_o[24] = 1'b0;
  assign data_mem_pkt_o[25] = 1'b0;
  assign data_mem_pkt_o[26] = 1'b0;
  assign data_mem_pkt_o[27] = 1'b0;
  assign data_mem_pkt_o[28] = 1'b0;
  assign data_mem_pkt_o[29] = 1'b0;
  assign data_mem_pkt_o[30] = 1'b0;
  assign data_mem_pkt_o[31] = 1'b0;
  assign data_mem_pkt_o[32] = 1'b0;
  assign data_mem_pkt_o[33] = 1'b0;
  assign data_mem_pkt_o[34] = 1'b0;
  assign data_mem_pkt_o[35] = 1'b0;
  assign data_mem_pkt_o[36] = 1'b0;
  assign data_mem_pkt_o[37] = 1'b0;
  assign data_mem_pkt_o[38] = 1'b0;
  assign data_mem_pkt_o[39] = 1'b0;
  assign data_mem_pkt_o[40] = 1'b0;
  assign data_mem_pkt_o[41] = 1'b0;
  assign data_mem_pkt_o[42] = 1'b0;
  assign data_mem_pkt_o[43] = 1'b0;
  assign data_mem_pkt_o[44] = 1'b0;
  assign data_mem_pkt_o[45] = 1'b0;
  assign data_mem_pkt_o[46] = 1'b0;
  assign data_mem_pkt_o[47] = 1'b0;
  assign data_mem_pkt_o[48] = 1'b0;
  assign data_mem_pkt_o[49] = 1'b0;
  assign data_mem_pkt_o[50] = 1'b0;
  assign data_mem_pkt_o[51] = 1'b0;
  assign data_mem_pkt_o[52] = 1'b0;
  assign data_mem_pkt_o[53] = 1'b0;
  assign data_mem_pkt_o[54] = 1'b0;
  assign data_mem_pkt_o[55] = 1'b0;
  assign data_mem_pkt_o[56] = 1'b0;
  assign data_mem_pkt_o[57] = 1'b0;
  assign data_mem_pkt_o[58] = 1'b0;
  assign data_mem_pkt_o[59] = 1'b0;
  assign data_mem_pkt_o[60] = 1'b0;
  assign data_mem_pkt_o[61] = 1'b0;
  assign data_mem_pkt_o[62] = 1'b0;
  assign data_mem_pkt_o[63] = 1'b0;
  assign data_mem_pkt_o[64] = 1'b0;
  assign data_mem_pkt_o[74] = 1'b0;
  assign data_mem_pkt_o[75] = 1'b0;
  assign data_mem_pkt_o[76] = 1'b0;
  assign data_mem_pkt_o[77] = 1'b0;
  assign data_mem_pkt_o[78] = 1'b0;
  assign data_mem_pkt_o[79] = 1'b0;
  assign data_mem_pkt_o[80] = 1'b0;
  assign data_mem_pkt_o[81] = 1'b0;
  assign data_mem_pkt_o[82] = 1'b0;
  assign data_mem_pkt_o[83] = 1'b0;
  assign data_mem_pkt_o[84] = 1'b0;
  assign data_mem_pkt_o[85] = 1'b0;
  assign data_mem_pkt_o[86] = 1'b0;
  assign data_mem_pkt_o[87] = 1'b0;
  assign data_mem_pkt_o[88] = 1'b0;
  assign data_mem_pkt_o[89] = 1'b0;
  assign data_mem_pkt_o[90] = 1'b0;
  assign data_mem_pkt_o[91] = 1'b0;
  assign data_mem_pkt_o[92] = 1'b0;
  assign data_mem_pkt_o[93] = 1'b0;
  assign data_mem_pkt_o[94] = 1'b0;
  assign data_mem_pkt_o[95] = 1'b0;
  assign data_mem_pkt_o[96] = 1'b0;
  assign data_mem_pkt_o[97] = 1'b0;
  assign data_mem_pkt_o[98] = 1'b0;
  assign data_mem_pkt_o[99] = 1'b0;
  assign data_mem_pkt_o[100] = 1'b0;
  assign data_mem_pkt_o[101] = 1'b0;
  assign data_mem_pkt_o[102] = 1'b0;
  assign data_mem_pkt_o[103] = 1'b0;
  assign data_mem_pkt_o[104] = 1'b0;
  assign data_mem_pkt_o[105] = 1'b0;
  assign data_mem_pkt_o[106] = 1'b0;
  assign data_mem_pkt_o[107] = 1'b0;
  assign data_mem_pkt_o[108] = 1'b0;
  assign data_mem_pkt_o[109] = 1'b0;
  assign data_mem_pkt_o[110] = 1'b0;
  assign data_mem_pkt_o[111] = 1'b0;
  assign data_mem_pkt_o[112] = 1'b0;
  assign data_mem_pkt_o[113] = 1'b0;
  assign data_mem_pkt_o[114] = 1'b0;
  assign data_mem_pkt_o[115] = 1'b0;
  assign data_mem_pkt_o[116] = 1'b0;
  assign data_mem_pkt_o[117] = 1'b0;
  assign data_mem_pkt_o[118] = 1'b0;
  assign data_mem_pkt_o[119] = 1'b0;
  assign data_mem_pkt_o[120] = 1'b0;
  assign data_mem_pkt_o[121] = 1'b0;
  assign data_mem_pkt_o[122] = 1'b0;
  assign data_mem_pkt_o[123] = 1'b0;
  assign data_mem_pkt_o[124] = 1'b0;
  assign data_mem_pkt_o[125] = 1'b0;
  assign data_mem_pkt_o[126] = 1'b0;
  assign data_mem_pkt_o[127] = 1'b0;
  assign data_mem_pkt_o[128] = 1'b0;
  assign data_mem_pkt_o[129] = 1'b0;
  assign data_mem_pkt_o[130] = 1'b0;
  assign data_mem_pkt_o[131] = 1'b0;
  assign data_mem_pkt_o[132] = 1'b0;
  assign data_mem_pkt_o[133] = 1'b0;
  assign data_mem_pkt_o[134] = 1'b0;
  assign data_mem_pkt_o[135] = 1'b0;
  assign data_mem_pkt_o[136] = 1'b0;
  assign data_mem_pkt_o[137] = 1'b0;
  assign data_mem_pkt_o[138] = 1'b0;
  assign data_mem_pkt_o[139] = 1'b0;
  assign data_mem_pkt_o[140] = 1'b0;
  assign data_mem_pkt_o[141] = 1'b0;
  assign data_mem_pkt_o[142] = 1'b0;
  assign data_mem_pkt_o[143] = 1'b0;
  assign data_mem_pkt_o[144] = 1'b0;
  assign data_mem_pkt_o[145] = 1'b0;
  assign data_mem_pkt_o[146] = 1'b0;
  assign data_mem_pkt_o[147] = 1'b0;
  assign data_mem_pkt_o[148] = 1'b0;
  assign data_mem_pkt_o[149] = 1'b0;
  assign data_mem_pkt_o[150] = 1'b0;
  assign data_mem_pkt_o[151] = 1'b0;
  assign data_mem_pkt_o[152] = 1'b0;
  assign data_mem_pkt_o[153] = 1'b0;
  assign data_mem_pkt_o[154] = 1'b0;
  assign data_mem_pkt_o[155] = 1'b0;
  assign data_mem_pkt_o[156] = 1'b0;
  assign data_mem_pkt_o[157] = 1'b0;
  assign data_mem_pkt_o[158] = 1'b0;
  assign data_mem_pkt_o[159] = 1'b0;
  assign data_mem_pkt_o[160] = 1'b0;
  assign data_mem_pkt_o[161] = 1'b0;
  assign data_mem_pkt_o[162] = 1'b0;
  assign data_mem_pkt_o[163] = 1'b0;
  assign data_mem_pkt_o[164] = 1'b0;
  assign data_mem_pkt_o[165] = 1'b0;
  assign data_mem_pkt_o[166] = 1'b0;
  assign data_mem_pkt_o[167] = 1'b0;
  assign data_mem_pkt_o[168] = 1'b0;
  assign data_mem_pkt_o[169] = 1'b0;
  assign data_mem_pkt_o[170] = 1'b0;
  assign data_mem_pkt_o[171] = 1'b0;
  assign data_mem_pkt_o[172] = 1'b0;
  assign data_mem_pkt_o[173] = 1'b0;
  assign data_mem_pkt_o[174] = 1'b0;
  assign data_mem_pkt_o[175] = 1'b0;
  assign data_mem_pkt_o[176] = 1'b0;
  assign data_mem_pkt_o[177] = 1'b0;
  assign data_mem_pkt_o[178] = 1'b0;
  assign data_mem_pkt_o[179] = 1'b0;
  assign data_mem_pkt_o[180] = 1'b0;
  assign data_mem_pkt_o[181] = 1'b0;
  assign data_mem_pkt_o[182] = 1'b0;
  assign data_mem_pkt_o[183] = 1'b0;
  assign data_mem_pkt_o[184] = 1'b0;
  assign data_mem_pkt_o[185] = 1'b0;
  assign data_mem_pkt_o[186] = 1'b0;
  assign data_mem_pkt_o[187] = 1'b0;
  assign data_mem_pkt_o[188] = 1'b0;
  assign data_mem_pkt_o[189] = 1'b0;
  assign data_mem_pkt_o[190] = 1'b0;
  assign data_mem_pkt_o[191] = 1'b0;
  assign data_mem_pkt_o[192] = 1'b0;
  assign data_mem_pkt_o[193] = 1'b0;
  assign data_mem_pkt_o[194] = 1'b0;
  assign data_mem_pkt_o[195] = 1'b0;
  assign data_mem_pkt_o[196] = 1'b0;
  assign data_mem_pkt_o[197] = 1'b0;
  assign data_mem_pkt_o[198] = 1'b0;
  assign data_mem_pkt_o[199] = 1'b0;
  assign data_mem_pkt_o[200] = 1'b0;
  assign data_mem_pkt_o[201] = 1'b0;
  assign data_mem_pkt_o[202] = 1'b0;
  assign data_mem_pkt_o[203] = 1'b0;
  assign data_mem_pkt_o[204] = 1'b0;
  assign data_mem_pkt_o[205] = 1'b0;
  assign data_mem_pkt_o[206] = 1'b0;
  assign data_mem_pkt_o[207] = 1'b0;
  assign data_mem_pkt_o[208] = 1'b0;
  assign data_mem_pkt_o[209] = 1'b0;
  assign data_mem_pkt_o[210] = 1'b0;
  assign data_mem_pkt_o[211] = 1'b0;
  assign data_mem_pkt_o[212] = 1'b0;
  assign data_mem_pkt_o[213] = 1'b0;
  assign data_mem_pkt_o[214] = 1'b0;
  assign data_mem_pkt_o[215] = 1'b0;
  assign data_mem_pkt_o[216] = 1'b0;
  assign data_mem_pkt_o[217] = 1'b0;
  assign data_mem_pkt_o[218] = 1'b0;
  assign data_mem_pkt_o[219] = 1'b0;
  assign data_mem_pkt_o[220] = 1'b0;
  assign data_mem_pkt_o[221] = 1'b0;
  assign data_mem_pkt_o[222] = 1'b0;
  assign data_mem_pkt_o[223] = 1'b0;
  assign data_mem_pkt_o[224] = 1'b0;
  assign data_mem_pkt_o[225] = 1'b0;
  assign data_mem_pkt_o[226] = 1'b0;
  assign data_mem_pkt_o[227] = 1'b0;
  assign data_mem_pkt_o[228] = 1'b0;
  assign data_mem_pkt_o[229] = 1'b0;
  assign data_mem_pkt_o[230] = 1'b0;
  assign data_mem_pkt_o[231] = 1'b0;
  assign data_mem_pkt_o[232] = 1'b0;
  assign data_mem_pkt_o[233] = 1'b0;
  assign data_mem_pkt_o[234] = 1'b0;
  assign data_mem_pkt_o[235] = 1'b0;
  assign data_mem_pkt_o[236] = 1'b0;
  assign data_mem_pkt_o[237] = 1'b0;
  assign data_mem_pkt_o[238] = 1'b0;
  assign data_mem_pkt_o[239] = 1'b0;
  assign data_mem_pkt_o[240] = 1'b0;
  assign data_mem_pkt_o[241] = 1'b0;
  assign data_mem_pkt_o[242] = 1'b0;
  assign data_mem_pkt_o[243] = 1'b0;
  assign data_mem_pkt_o[244] = 1'b0;
  assign data_mem_pkt_o[245] = 1'b0;
  assign data_mem_pkt_o[246] = 1'b0;
  assign data_mem_pkt_o[247] = 1'b0;
  assign data_mem_pkt_o[248] = 1'b0;
  assign data_mem_pkt_o[249] = 1'b0;
  assign data_mem_pkt_o[250] = 1'b0;
  assign data_mem_pkt_o[251] = 1'b0;
  assign data_mem_pkt_o[252] = 1'b0;
  assign data_mem_pkt_o[253] = 1'b0;
  assign data_mem_pkt_o[254] = 1'b0;
  assign data_mem_pkt_o[255] = 1'b0;
  assign data_mem_pkt_o[256] = 1'b0;
  assign data_mem_pkt_o[257] = 1'b0;
  assign data_mem_pkt_o[258] = 1'b0;
  assign data_mem_pkt_o[259] = 1'b0;
  assign data_mem_pkt_o[260] = 1'b0;
  assign data_mem_pkt_o[261] = 1'b0;
  assign data_mem_pkt_o[262] = 1'b0;
  assign data_mem_pkt_o[263] = 1'b0;
  assign data_mem_pkt_o[264] = 1'b0;
  assign data_mem_pkt_o[265] = 1'b0;
  assign data_mem_pkt_o[266] = 1'b0;
  assign data_mem_pkt_o[267] = 1'b0;
  assign data_mem_pkt_o[268] = 1'b0;
  assign data_mem_pkt_o[269] = 1'b0;
  assign data_mem_pkt_o[270] = 1'b0;
  assign data_mem_pkt_o[271] = 1'b0;
  assign data_mem_pkt_o[272] = 1'b0;
  assign data_mem_pkt_o[273] = 1'b0;
  assign data_mem_pkt_o[274] = 1'b0;
  assign data_mem_pkt_o[275] = 1'b0;
  assign data_mem_pkt_o[276] = 1'b0;
  assign data_mem_pkt_o[277] = 1'b0;
  assign data_mem_pkt_o[278] = 1'b0;
  assign data_mem_pkt_o[279] = 1'b0;
  assign data_mem_pkt_o[280] = 1'b0;
  assign data_mem_pkt_o[281] = 1'b0;
  assign data_mem_pkt_o[282] = 1'b0;
  assign data_mem_pkt_o[283] = 1'b0;
  assign data_mem_pkt_o[284] = 1'b0;
  assign data_mem_pkt_o[285] = 1'b0;
  assign data_mem_pkt_o[286] = 1'b0;
  assign data_mem_pkt_o[287] = 1'b0;
  assign data_mem_pkt_o[288] = 1'b0;
  assign data_mem_pkt_o[289] = 1'b0;
  assign data_mem_pkt_o[290] = 1'b0;
  assign data_mem_pkt_o[291] = 1'b0;
  assign data_mem_pkt_o[292] = 1'b0;
  assign data_mem_pkt_o[293] = 1'b0;
  assign data_mem_pkt_o[294] = 1'b0;
  assign data_mem_pkt_o[295] = 1'b0;
  assign data_mem_pkt_o[296] = 1'b0;
  assign data_mem_pkt_o[297] = 1'b0;
  assign data_mem_pkt_o[298] = 1'b0;
  assign data_mem_pkt_o[299] = 1'b0;
  assign data_mem_pkt_o[300] = 1'b0;
  assign data_mem_pkt_o[301] = 1'b0;
  assign data_mem_pkt_o[302] = 1'b0;
  assign data_mem_pkt_o[303] = 1'b0;
  assign data_mem_pkt_o[304] = 1'b0;
  assign data_mem_pkt_o[305] = 1'b0;
  assign data_mem_pkt_o[306] = 1'b0;
  assign data_mem_pkt_o[307] = 1'b0;
  assign data_mem_pkt_o[308] = 1'b0;
  assign data_mem_pkt_o[309] = 1'b0;
  assign data_mem_pkt_o[310] = 1'b0;
  assign data_mem_pkt_o[311] = 1'b0;
  assign data_mem_pkt_o[312] = 1'b0;
  assign data_mem_pkt_o[313] = 1'b0;
  assign data_mem_pkt_o[314] = 1'b0;
  assign data_mem_pkt_o[315] = 1'b0;
  assign data_mem_pkt_o[316] = 1'b0;
  assign data_mem_pkt_o[317] = 1'b0;
  assign data_mem_pkt_o[318] = 1'b0;
  assign data_mem_pkt_o[319] = 1'b0;
  assign data_mem_pkt_o[320] = 1'b0;
  assign data_mem_pkt_o[321] = 1'b0;
  assign data_mem_pkt_o[322] = 1'b0;
  assign data_mem_pkt_o[323] = 1'b0;
  assign data_mem_pkt_o[324] = 1'b0;
  assign data_mem_pkt_o[325] = 1'b0;
  assign data_mem_pkt_o[326] = 1'b0;
  assign data_mem_pkt_o[327] = 1'b0;
  assign data_mem_pkt_o[328] = 1'b0;
  assign data_mem_pkt_o[329] = 1'b0;
  assign data_mem_pkt_o[330] = 1'b0;
  assign data_mem_pkt_o[331] = 1'b0;
  assign data_mem_pkt_o[332] = 1'b0;
  assign data_mem_pkt_o[333] = 1'b0;
  assign data_mem_pkt_o[334] = 1'b0;
  assign data_mem_pkt_o[335] = 1'b0;
  assign data_mem_pkt_o[336] = 1'b0;
  assign data_mem_pkt_o[337] = 1'b0;
  assign data_mem_pkt_o[338] = 1'b0;
  assign data_mem_pkt_o[339] = 1'b0;
  assign data_mem_pkt_o[340] = 1'b0;
  assign data_mem_pkt_o[341] = 1'b0;
  assign data_mem_pkt_o[342] = 1'b0;
  assign data_mem_pkt_o[343] = 1'b0;
  assign data_mem_pkt_o[344] = 1'b0;
  assign data_mem_pkt_o[345] = 1'b0;
  assign data_mem_pkt_o[346] = 1'b0;
  assign data_mem_pkt_o[347] = 1'b0;
  assign data_mem_pkt_o[348] = 1'b0;
  assign data_mem_pkt_o[349] = 1'b0;
  assign data_mem_pkt_o[350] = 1'b0;
  assign data_mem_pkt_o[351] = 1'b0;
  assign data_mem_pkt_o[352] = 1'b0;
  assign data_mem_pkt_o[353] = 1'b0;
  assign data_mem_pkt_o[354] = 1'b0;
  assign data_mem_pkt_o[355] = 1'b0;
  assign data_mem_pkt_o[356] = 1'b0;
  assign data_mem_pkt_o[357] = 1'b0;
  assign data_mem_pkt_o[358] = 1'b0;
  assign data_mem_pkt_o[359] = 1'b0;
  assign data_mem_pkt_o[360] = 1'b0;
  assign data_mem_pkt_o[361] = 1'b0;
  assign data_mem_pkt_o[362] = 1'b0;
  assign data_mem_pkt_o[363] = 1'b0;
  assign data_mem_pkt_o[364] = 1'b0;
  assign data_mem_pkt_o[365] = 1'b0;
  assign data_mem_pkt_o[366] = 1'b0;
  assign data_mem_pkt_o[367] = 1'b0;
  assign data_mem_pkt_o[368] = 1'b0;
  assign data_mem_pkt_o[369] = 1'b0;
  assign data_mem_pkt_o[370] = 1'b0;
  assign data_mem_pkt_o[371] = 1'b0;
  assign data_mem_pkt_o[372] = 1'b0;
  assign data_mem_pkt_o[373] = 1'b0;
  assign data_mem_pkt_o[374] = 1'b0;
  assign data_mem_pkt_o[375] = 1'b0;
  assign data_mem_pkt_o[376] = 1'b0;
  assign data_mem_pkt_o[377] = 1'b0;
  assign data_mem_pkt_o[378] = 1'b0;
  assign data_mem_pkt_o[379] = 1'b0;
  assign data_mem_pkt_o[380] = 1'b0;
  assign data_mem_pkt_o[381] = 1'b0;
  assign data_mem_pkt_o[382] = 1'b0;
  assign data_mem_pkt_o[383] = 1'b0;
  assign data_mem_pkt_o[384] = 1'b0;
  assign data_mem_pkt_o[385] = 1'b0;
  assign data_mem_pkt_o[386] = 1'b0;
  assign data_mem_pkt_o[387] = 1'b0;
  assign data_mem_pkt_o[388] = 1'b0;
  assign data_mem_pkt_o[389] = 1'b0;
  assign data_mem_pkt_o[390] = 1'b0;
  assign data_mem_pkt_o[391] = 1'b0;
  assign data_mem_pkt_o[392] = 1'b0;
  assign data_mem_pkt_o[393] = 1'b0;
  assign data_mem_pkt_o[394] = 1'b0;
  assign data_mem_pkt_o[395] = 1'b0;
  assign data_mem_pkt_o[396] = 1'b0;
  assign data_mem_pkt_o[397] = 1'b0;
  assign data_mem_pkt_o[398] = 1'b0;
  assign data_mem_pkt_o[399] = 1'b0;
  assign data_mem_pkt_o[400] = 1'b0;
  assign data_mem_pkt_o[401] = 1'b0;
  assign data_mem_pkt_o[402] = 1'b0;
  assign data_mem_pkt_o[403] = 1'b0;
  assign data_mem_pkt_o[404] = 1'b0;
  assign data_mem_pkt_o[405] = 1'b0;
  assign data_mem_pkt_o[406] = 1'b0;
  assign data_mem_pkt_o[407] = 1'b0;
  assign data_mem_pkt_o[408] = 1'b0;
  assign data_mem_pkt_o[409] = 1'b0;
  assign data_mem_pkt_o[410] = 1'b0;
  assign data_mem_pkt_o[411] = 1'b0;
  assign data_mem_pkt_o[412] = 1'b0;
  assign data_mem_pkt_o[413] = 1'b0;
  assign data_mem_pkt_o[414] = 1'b0;
  assign data_mem_pkt_o[415] = 1'b0;
  assign data_mem_pkt_o[416] = 1'b0;
  assign data_mem_pkt_o[417] = 1'b0;
  assign data_mem_pkt_o[418] = 1'b0;
  assign data_mem_pkt_o[419] = 1'b0;
  assign data_mem_pkt_o[420] = 1'b0;
  assign data_mem_pkt_o[421] = 1'b0;
  assign data_mem_pkt_o[422] = 1'b0;
  assign data_mem_pkt_o[423] = 1'b0;
  assign data_mem_pkt_o[424] = 1'b0;
  assign data_mem_pkt_o[425] = 1'b0;
  assign data_mem_pkt_o[426] = 1'b0;
  assign data_mem_pkt_o[427] = 1'b0;
  assign data_mem_pkt_o[428] = 1'b0;
  assign data_mem_pkt_o[429] = 1'b0;
  assign data_mem_pkt_o[430] = 1'b0;
  assign data_mem_pkt_o[431] = 1'b0;
  assign data_mem_pkt_o[432] = 1'b0;
  assign data_mem_pkt_o[433] = 1'b0;
  assign data_mem_pkt_o[434] = 1'b0;
  assign data_mem_pkt_o[435] = 1'b0;
  assign data_mem_pkt_o[436] = 1'b0;
  assign data_mem_pkt_o[437] = 1'b0;
  assign data_mem_pkt_o[438] = 1'b0;
  assign data_mem_pkt_o[439] = 1'b0;
  assign data_mem_pkt_o[440] = 1'b0;
  assign data_mem_pkt_o[441] = 1'b0;
  assign data_mem_pkt_o[442] = 1'b0;
  assign data_mem_pkt_o[443] = 1'b0;
  assign data_mem_pkt_o[444] = 1'b0;
  assign data_mem_pkt_o[445] = 1'b0;
  assign data_mem_pkt_o[446] = 1'b0;
  assign data_mem_pkt_o[447] = 1'b0;
  assign data_mem_pkt_o[448] = 1'b0;
  assign data_mem_pkt_o[449] = 1'b0;
  assign data_mem_pkt_o[450] = 1'b0;
  assign data_mem_pkt_o[451] = 1'b0;
  assign data_mem_pkt_o[452] = 1'b0;
  assign data_mem_pkt_o[453] = 1'b0;
  assign data_mem_pkt_o[454] = 1'b0;
  assign data_mem_pkt_o[455] = 1'b0;
  assign data_mem_pkt_o[456] = 1'b0;
  assign data_mem_pkt_o[457] = 1'b0;
  assign data_mem_pkt_o[458] = 1'b0;
  assign data_mem_pkt_o[459] = 1'b0;
  assign data_mem_pkt_o[460] = 1'b0;
  assign data_mem_pkt_o[461] = 1'b0;
  assign data_mem_pkt_o[462] = 1'b0;
  assign data_mem_pkt_o[463] = 1'b0;
  assign data_mem_pkt_o[464] = 1'b0;
  assign data_mem_pkt_o[465] = 1'b0;
  assign data_mem_pkt_o[466] = 1'b0;
  assign data_mem_pkt_o[467] = 1'b0;
  assign data_mem_pkt_o[468] = 1'b0;
  assign data_mem_pkt_o[469] = 1'b0;
  assign data_mem_pkt_o[470] = 1'b0;
  assign data_mem_pkt_o[471] = 1'b0;
  assign data_mem_pkt_o[472] = 1'b0;
  assign data_mem_pkt_o[473] = 1'b0;
  assign data_mem_pkt_o[474] = 1'b0;
  assign data_mem_pkt_o[475] = 1'b0;
  assign data_mem_pkt_o[476] = 1'b0;
  assign data_mem_pkt_o[477] = 1'b0;
  assign data_mem_pkt_o[478] = 1'b0;
  assign data_mem_pkt_o[479] = 1'b0;
  assign data_mem_pkt_o[480] = 1'b0;
  assign data_mem_pkt_o[481] = 1'b0;
  assign data_mem_pkt_o[482] = 1'b0;
  assign data_mem_pkt_o[483] = 1'b0;
  assign data_mem_pkt_o[484] = 1'b0;
  assign data_mem_pkt_o[485] = 1'b0;
  assign data_mem_pkt_o[486] = 1'b0;
  assign data_mem_pkt_o[487] = 1'b0;
  assign data_mem_pkt_o[488] = 1'b0;
  assign data_mem_pkt_o[489] = 1'b0;
  assign data_mem_pkt_o[490] = 1'b0;
  assign data_mem_pkt_o[491] = 1'b0;
  assign data_mem_pkt_o[492] = 1'b0;
  assign data_mem_pkt_o[493] = 1'b0;
  assign data_mem_pkt_o[494] = 1'b0;
  assign data_mem_pkt_o[495] = 1'b0;
  assign data_mem_pkt_o[496] = 1'b0;
  assign data_mem_pkt_o[497] = 1'b0;
  assign data_mem_pkt_o[498] = 1'b0;
  assign data_mem_pkt_o[499] = 1'b0;
  assign data_mem_pkt_o[500] = 1'b0;
  assign data_mem_pkt_o[501] = 1'b0;
  assign data_mem_pkt_o[502] = 1'b0;
  assign data_mem_pkt_o[503] = 1'b0;
  assign data_mem_pkt_o[504] = 1'b0;
  assign data_mem_pkt_o[505] = 1'b0;
  assign data_mem_pkt_o[506] = 1'b0;
  assign data_mem_pkt_o[507] = 1'b0;
  assign data_mem_pkt_o[508] = 1'b0;
  assign data_mem_pkt_o[509] = 1'b0;
  assign data_mem_pkt_o[510] = 1'b0;
  assign data_mem_pkt_o[511] = 1'b0;
  assign data_mem_pkt_o[512] = 1'b0;
  assign data_mem_pkt_o[513] = 1'b0;
  assign data_mem_pkt_o[514] = 1'b0;
  assign data_mem_pkt_o[515] = 1'b0;
  assign data_mem_pkt_o[516] = 1'b0;
  assign data_mem_pkt_o[517] = 1'b0;
  assign data_mem_pkt_o[518] = 1'b0;
  assign data_mem_pkt_o[519] = 1'b0;
  assign data_mem_pkt_o[520] = 1'b0;
  assign data_mem_pkt_o[521] = 1'b0;
  assign lce_data_resp_o[0] = 1'b0;
  assign lce_data_resp_o[1] = 1'b0;
  assign lce_data_resp_o[2] = 1'b0;
  assign lce_data_resp_o[3] = 1'b0;
  assign lce_data_resp_o[4] = 1'b0;
  assign lce_data_resp_o[5] = 1'b0;
  assign lce_data_resp_o[6] = 1'b0;
  assign lce_data_resp_o[7] = 1'b0;
  assign lce_data_resp_o[8] = 1'b0;
  assign lce_data_resp_o[9] = 1'b0;
  assign lce_data_resp_o[10] = 1'b0;
  assign lce_data_resp_o[11] = 1'b0;
  assign lce_data_resp_o[12] = 1'b0;
  assign lce_data_resp_o[13] = 1'b0;
  assign lce_data_resp_o[14] = 1'b0;
  assign lce_data_resp_o[15] = 1'b0;
  assign lce_data_resp_o[16] = 1'b0;
  assign lce_data_resp_o[17] = 1'b0;
  assign lce_data_resp_o[18] = 1'b0;
  assign lce_data_resp_o[19] = 1'b0;
  assign lce_data_resp_o[20] = 1'b0;
  assign lce_data_resp_o[21] = 1'b0;
  assign lce_data_resp_o[22] = 1'b0;
  assign lce_data_resp_o[23] = 1'b0;
  assign lce_data_resp_o[24] = 1'b0;
  assign lce_data_resp_o[25] = 1'b0;
  assign lce_data_resp_o[26] = 1'b0;
  assign lce_data_resp_o[27] = 1'b0;
  assign lce_data_resp_o[28] = 1'b0;
  assign lce_data_resp_o[29] = 1'b0;
  assign lce_data_resp_o[30] = 1'b0;
  assign lce_data_resp_o[31] = 1'b0;
  assign lce_data_resp_o[32] = 1'b0;
  assign lce_data_resp_o[33] = 1'b0;
  assign lce_data_resp_o[34] = 1'b0;
  assign lce_data_resp_o[35] = 1'b0;
  assign lce_data_resp_o[36] = 1'b0;
  assign lce_data_resp_o[37] = 1'b0;
  assign lce_data_resp_o[38] = 1'b0;
  assign lce_data_resp_o[39] = 1'b0;
  assign lce_data_resp_o[40] = 1'b0;
  assign lce_data_resp_o[41] = 1'b0;
  assign lce_data_resp_o[42] = 1'b0;
  assign lce_data_resp_o[43] = 1'b0;
  assign lce_data_resp_o[44] = 1'b0;
  assign lce_data_resp_o[45] = 1'b0;
  assign lce_data_resp_o[46] = 1'b0;
  assign lce_data_resp_o[47] = 1'b0;
  assign lce_data_resp_o[48] = 1'b0;
  assign lce_data_resp_o[49] = 1'b0;
  assign lce_data_resp_o[50] = 1'b0;
  assign lce_data_resp_o[51] = 1'b0;
  assign lce_data_resp_o[52] = 1'b0;
  assign lce_data_resp_o[53] = 1'b0;
  assign lce_data_resp_o[54] = 1'b0;
  assign lce_data_resp_o[55] = 1'b0;
  assign lce_data_resp_o[56] = 1'b0;
  assign lce_data_resp_o[57] = 1'b0;
  assign lce_data_resp_o[58] = 1'b0;
  assign lce_data_resp_o[59] = 1'b0;
  assign lce_data_resp_o[60] = 1'b0;
  assign lce_data_resp_o[61] = 1'b0;
  assign lce_data_resp_o[62] = 1'b0;
  assign lce_data_resp_o[63] = 1'b0;
  assign lce_data_resp_o[64] = 1'b0;
  assign lce_data_resp_o[65] = 1'b0;
  assign lce_data_resp_o[66] = 1'b0;
  assign lce_data_resp_o[67] = 1'b0;
  assign lce_data_resp_o[68] = 1'b0;
  assign lce_data_resp_o[69] = 1'b0;
  assign lce_data_resp_o[70] = 1'b0;
  assign lce_data_resp_o[71] = 1'b0;
  assign lce_data_resp_o[72] = 1'b0;
  assign lce_data_resp_o[73] = 1'b0;
  assign lce_data_resp_o[74] = 1'b0;
  assign lce_data_resp_o[75] = 1'b0;
  assign lce_data_resp_o[76] = 1'b0;
  assign lce_data_resp_o[77] = 1'b0;
  assign lce_data_resp_o[78] = 1'b0;
  assign lce_data_resp_o[79] = 1'b0;
  assign lce_data_resp_o[80] = 1'b0;
  assign lce_data_resp_o[81] = 1'b0;
  assign lce_data_resp_o[82] = 1'b0;
  assign lce_data_resp_o[83] = 1'b0;
  assign lce_data_resp_o[84] = 1'b0;
  assign lce_data_resp_o[85] = 1'b0;
  assign lce_data_resp_o[86] = 1'b0;
  assign lce_data_resp_o[87] = 1'b0;
  assign lce_data_resp_o[88] = 1'b0;
  assign lce_data_resp_o[89] = 1'b0;
  assign lce_data_resp_o[90] = 1'b0;
  assign lce_data_resp_o[91] = 1'b0;
  assign lce_data_resp_o[92] = 1'b0;
  assign lce_data_resp_o[93] = 1'b0;
  assign lce_data_resp_o[94] = 1'b0;
  assign lce_data_resp_o[95] = 1'b0;
  assign lce_data_resp_o[96] = 1'b0;
  assign lce_data_resp_o[97] = 1'b0;
  assign lce_data_resp_o[98] = 1'b0;
  assign lce_data_resp_o[99] = 1'b0;
  assign lce_data_resp_o[100] = 1'b0;
  assign lce_data_resp_o[101] = 1'b0;
  assign lce_data_resp_o[102] = 1'b0;
  assign lce_data_resp_o[103] = 1'b0;
  assign lce_data_resp_o[104] = 1'b0;
  assign lce_data_resp_o[105] = 1'b0;
  assign lce_data_resp_o[106] = 1'b0;
  assign lce_data_resp_o[107] = 1'b0;
  assign lce_data_resp_o[108] = 1'b0;
  assign lce_data_resp_o[109] = 1'b0;
  assign lce_data_resp_o[110] = 1'b0;
  assign lce_data_resp_o[111] = 1'b0;
  assign lce_data_resp_o[112] = 1'b0;
  assign lce_data_resp_o[113] = 1'b0;
  assign lce_data_resp_o[114] = 1'b0;
  assign lce_data_resp_o[115] = 1'b0;
  assign lce_data_resp_o[116] = 1'b0;
  assign lce_data_resp_o[117] = 1'b0;
  assign lce_data_resp_o[118] = 1'b0;
  assign lce_data_resp_o[119] = 1'b0;
  assign lce_data_resp_o[120] = 1'b0;
  assign lce_data_resp_o[121] = 1'b0;
  assign lce_data_resp_o[122] = 1'b0;
  assign lce_data_resp_o[123] = 1'b0;
  assign lce_data_resp_o[124] = 1'b0;
  assign lce_data_resp_o[125] = 1'b0;
  assign lce_data_resp_o[126] = 1'b0;
  assign lce_data_resp_o[127] = 1'b0;
  assign lce_data_resp_o[128] = 1'b0;
  assign lce_data_resp_o[129] = 1'b0;
  assign lce_data_resp_o[130] = 1'b0;
  assign lce_data_resp_o[131] = 1'b0;
  assign lce_data_resp_o[132] = 1'b0;
  assign lce_data_resp_o[133] = 1'b0;
  assign lce_data_resp_o[134] = 1'b0;
  assign lce_data_resp_o[135] = 1'b0;
  assign lce_data_resp_o[136] = 1'b0;
  assign lce_data_resp_o[137] = 1'b0;
  assign lce_data_resp_o[138] = 1'b0;
  assign lce_data_resp_o[139] = 1'b0;
  assign lce_data_resp_o[140] = 1'b0;
  assign lce_data_resp_o[141] = 1'b0;
  assign lce_data_resp_o[142] = 1'b0;
  assign lce_data_resp_o[143] = 1'b0;
  assign lce_data_resp_o[144] = 1'b0;
  assign lce_data_resp_o[145] = 1'b0;
  assign lce_data_resp_o[146] = 1'b0;
  assign lce_data_resp_o[147] = 1'b0;
  assign lce_data_resp_o[148] = 1'b0;
  assign lce_data_resp_o[149] = 1'b0;
  assign lce_data_resp_o[150] = 1'b0;
  assign lce_data_resp_o[151] = 1'b0;
  assign lce_data_resp_o[152] = 1'b0;
  assign lce_data_resp_o[153] = 1'b0;
  assign lce_data_resp_o[154] = 1'b0;
  assign lce_data_resp_o[155] = 1'b0;
  assign lce_data_resp_o[156] = 1'b0;
  assign lce_data_resp_o[157] = 1'b0;
  assign lce_data_resp_o[158] = 1'b0;
  assign lce_data_resp_o[159] = 1'b0;
  assign lce_data_resp_o[160] = 1'b0;
  assign lce_data_resp_o[161] = 1'b0;
  assign lce_data_resp_o[162] = 1'b0;
  assign lce_data_resp_o[163] = 1'b0;
  assign lce_data_resp_o[164] = 1'b0;
  assign lce_data_resp_o[165] = 1'b0;
  assign lce_data_resp_o[166] = 1'b0;
  assign lce_data_resp_o[167] = 1'b0;
  assign lce_data_resp_o[168] = 1'b0;
  assign lce_data_resp_o[169] = 1'b0;
  assign lce_data_resp_o[170] = 1'b0;
  assign lce_data_resp_o[171] = 1'b0;
  assign lce_data_resp_o[172] = 1'b0;
  assign lce_data_resp_o[173] = 1'b0;
  assign lce_data_resp_o[174] = 1'b0;
  assign lce_data_resp_o[175] = 1'b0;
  assign lce_data_resp_o[176] = 1'b0;
  assign lce_data_resp_o[177] = 1'b0;
  assign lce_data_resp_o[178] = 1'b0;
  assign lce_data_resp_o[179] = 1'b0;
  assign lce_data_resp_o[180] = 1'b0;
  assign lce_data_resp_o[181] = 1'b0;
  assign lce_data_resp_o[182] = 1'b0;
  assign lce_data_resp_o[183] = 1'b0;
  assign lce_data_resp_o[184] = 1'b0;
  assign lce_data_resp_o[185] = 1'b0;
  assign lce_data_resp_o[186] = 1'b0;
  assign lce_data_resp_o[187] = 1'b0;
  assign lce_data_resp_o[188] = 1'b0;
  assign lce_data_resp_o[189] = 1'b0;
  assign lce_data_resp_o[190] = 1'b0;
  assign lce_data_resp_o[191] = 1'b0;
  assign lce_data_resp_o[192] = 1'b0;
  assign lce_data_resp_o[193] = 1'b0;
  assign lce_data_resp_o[194] = 1'b0;
  assign lce_data_resp_o[195] = 1'b0;
  assign lce_data_resp_o[196] = 1'b0;
  assign lce_data_resp_o[197] = 1'b0;
  assign lce_data_resp_o[198] = 1'b0;
  assign lce_data_resp_o[199] = 1'b0;
  assign lce_data_resp_o[200] = 1'b0;
  assign lce_data_resp_o[201] = 1'b0;
  assign lce_data_resp_o[202] = 1'b0;
  assign lce_data_resp_o[203] = 1'b0;
  assign lce_data_resp_o[204] = 1'b0;
  assign lce_data_resp_o[205] = 1'b0;
  assign lce_data_resp_o[206] = 1'b0;
  assign lce_data_resp_o[207] = 1'b0;
  assign lce_data_resp_o[208] = 1'b0;
  assign lce_data_resp_o[209] = 1'b0;
  assign lce_data_resp_o[210] = 1'b0;
  assign lce_data_resp_o[211] = 1'b0;
  assign lce_data_resp_o[212] = 1'b0;
  assign lce_data_resp_o[213] = 1'b0;
  assign lce_data_resp_o[214] = 1'b0;
  assign lce_data_resp_o[215] = 1'b0;
  assign lce_data_resp_o[216] = 1'b0;
  assign lce_data_resp_o[217] = 1'b0;
  assign lce_data_resp_o[218] = 1'b0;
  assign lce_data_resp_o[219] = 1'b0;
  assign lce_data_resp_o[220] = 1'b0;
  assign lce_data_resp_o[221] = 1'b0;
  assign lce_data_resp_o[222] = 1'b0;
  assign lce_data_resp_o[223] = 1'b0;
  assign lce_data_resp_o[224] = 1'b0;
  assign lce_data_resp_o[225] = 1'b0;
  assign lce_data_resp_o[226] = 1'b0;
  assign lce_data_resp_o[227] = 1'b0;
  assign lce_data_resp_o[228] = 1'b0;
  assign lce_data_resp_o[229] = 1'b0;
  assign lce_data_resp_o[230] = 1'b0;
  assign lce_data_resp_o[231] = 1'b0;
  assign lce_data_resp_o[232] = 1'b0;
  assign lce_data_resp_o[233] = 1'b0;
  assign lce_data_resp_o[234] = 1'b0;
  assign lce_data_resp_o[235] = 1'b0;
  assign lce_data_resp_o[236] = 1'b0;
  assign lce_data_resp_o[237] = 1'b0;
  assign lce_data_resp_o[238] = 1'b0;
  assign lce_data_resp_o[239] = 1'b0;
  assign lce_data_resp_o[240] = 1'b0;
  assign lce_data_resp_o[241] = 1'b0;
  assign lce_data_resp_o[242] = 1'b0;
  assign lce_data_resp_o[243] = 1'b0;
  assign lce_data_resp_o[244] = 1'b0;
  assign lce_data_resp_o[245] = 1'b0;
  assign lce_data_resp_o[246] = 1'b0;
  assign lce_data_resp_o[247] = 1'b0;
  assign lce_data_resp_o[248] = 1'b0;
  assign lce_data_resp_o[249] = 1'b0;
  assign lce_data_resp_o[250] = 1'b0;
  assign lce_data_resp_o[251] = 1'b0;
  assign lce_data_resp_o[252] = 1'b0;
  assign lce_data_resp_o[253] = 1'b0;
  assign lce_data_resp_o[254] = 1'b0;
  assign lce_data_resp_o[255] = 1'b0;
  assign lce_data_resp_o[256] = 1'b0;
  assign lce_data_resp_o[257] = 1'b0;
  assign lce_data_resp_o[258] = 1'b0;
  assign lce_data_resp_o[259] = 1'b0;
  assign lce_data_resp_o[260] = 1'b0;
  assign lce_data_resp_o[261] = 1'b0;
  assign lce_data_resp_o[262] = 1'b0;
  assign lce_data_resp_o[263] = 1'b0;
  assign lce_data_resp_o[264] = 1'b0;
  assign lce_data_resp_o[265] = 1'b0;
  assign lce_data_resp_o[266] = 1'b0;
  assign lce_data_resp_o[267] = 1'b0;
  assign lce_data_resp_o[268] = 1'b0;
  assign lce_data_resp_o[269] = 1'b0;
  assign lce_data_resp_o[270] = 1'b0;
  assign lce_data_resp_o[271] = 1'b0;
  assign lce_data_resp_o[272] = 1'b0;
  assign lce_data_resp_o[273] = 1'b0;
  assign lce_data_resp_o[274] = 1'b0;
  assign lce_data_resp_o[275] = 1'b0;
  assign lce_data_resp_o[276] = 1'b0;
  assign lce_data_resp_o[277] = 1'b0;
  assign lce_data_resp_o[278] = 1'b0;
  assign lce_data_resp_o[279] = 1'b0;
  assign lce_data_resp_o[280] = 1'b0;
  assign lce_data_resp_o[281] = 1'b0;
  assign lce_data_resp_o[282] = 1'b0;
  assign lce_data_resp_o[283] = 1'b0;
  assign lce_data_resp_o[284] = 1'b0;
  assign lce_data_resp_o[285] = 1'b0;
  assign lce_data_resp_o[286] = 1'b0;
  assign lce_data_resp_o[287] = 1'b0;
  assign lce_data_resp_o[288] = 1'b0;
  assign lce_data_resp_o[289] = 1'b0;
  assign lce_data_resp_o[290] = 1'b0;
  assign lce_data_resp_o[291] = 1'b0;
  assign lce_data_resp_o[292] = 1'b0;
  assign lce_data_resp_o[293] = 1'b0;
  assign lce_data_resp_o[294] = 1'b0;
  assign lce_data_resp_o[295] = 1'b0;
  assign lce_data_resp_o[296] = 1'b0;
  assign lce_data_resp_o[297] = 1'b0;
  assign lce_data_resp_o[298] = 1'b0;
  assign lce_data_resp_o[299] = 1'b0;
  assign lce_data_resp_o[300] = 1'b0;
  assign lce_data_resp_o[301] = 1'b0;
  assign lce_data_resp_o[302] = 1'b0;
  assign lce_data_resp_o[303] = 1'b0;
  assign lce_data_resp_o[304] = 1'b0;
  assign lce_data_resp_o[305] = 1'b0;
  assign lce_data_resp_o[306] = 1'b0;
  assign lce_data_resp_o[307] = 1'b0;
  assign lce_data_resp_o[308] = 1'b0;
  assign lce_data_resp_o[309] = 1'b0;
  assign lce_data_resp_o[310] = 1'b0;
  assign lce_data_resp_o[311] = 1'b0;
  assign lce_data_resp_o[312] = 1'b0;
  assign lce_data_resp_o[313] = 1'b0;
  assign lce_data_resp_o[314] = 1'b0;
  assign lce_data_resp_o[315] = 1'b0;
  assign lce_data_resp_o[316] = 1'b0;
  assign lce_data_resp_o[317] = 1'b0;
  assign lce_data_resp_o[318] = 1'b0;
  assign lce_data_resp_o[319] = 1'b0;
  assign lce_data_resp_o[320] = 1'b0;
  assign lce_data_resp_o[321] = 1'b0;
  assign lce_data_resp_o[322] = 1'b0;
  assign lce_data_resp_o[323] = 1'b0;
  assign lce_data_resp_o[324] = 1'b0;
  assign lce_data_resp_o[325] = 1'b0;
  assign lce_data_resp_o[326] = 1'b0;
  assign lce_data_resp_o[327] = 1'b0;
  assign lce_data_resp_o[328] = 1'b0;
  assign lce_data_resp_o[329] = 1'b0;
  assign lce_data_resp_o[330] = 1'b0;
  assign lce_data_resp_o[331] = 1'b0;
  assign lce_data_resp_o[332] = 1'b0;
  assign lce_data_resp_o[333] = 1'b0;
  assign lce_data_resp_o[334] = 1'b0;
  assign lce_data_resp_o[335] = 1'b0;
  assign lce_data_resp_o[336] = 1'b0;
  assign lce_data_resp_o[337] = 1'b0;
  assign lce_data_resp_o[338] = 1'b0;
  assign lce_data_resp_o[339] = 1'b0;
  assign lce_data_resp_o[340] = 1'b0;
  assign lce_data_resp_o[341] = 1'b0;
  assign lce_data_resp_o[342] = 1'b0;
  assign lce_data_resp_o[343] = 1'b0;
  assign lce_data_resp_o[344] = 1'b0;
  assign lce_data_resp_o[345] = 1'b0;
  assign lce_data_resp_o[346] = 1'b0;
  assign lce_data_resp_o[347] = 1'b0;
  assign lce_data_resp_o[348] = 1'b0;
  assign lce_data_resp_o[349] = 1'b0;
  assign lce_data_resp_o[350] = 1'b0;
  assign lce_data_resp_o[351] = 1'b0;
  assign lce_data_resp_o[352] = 1'b0;
  assign lce_data_resp_o[353] = 1'b0;
  assign lce_data_resp_o[354] = 1'b0;
  assign lce_data_resp_o[355] = 1'b0;
  assign lce_data_resp_o[356] = 1'b0;
  assign lce_data_resp_o[357] = 1'b0;
  assign lce_data_resp_o[358] = 1'b0;
  assign lce_data_resp_o[359] = 1'b0;
  assign lce_data_resp_o[360] = 1'b0;
  assign lce_data_resp_o[361] = 1'b0;
  assign lce_data_resp_o[362] = 1'b0;
  assign lce_data_resp_o[363] = 1'b0;
  assign lce_data_resp_o[364] = 1'b0;
  assign lce_data_resp_o[365] = 1'b0;
  assign lce_data_resp_o[366] = 1'b0;
  assign lce_data_resp_o[367] = 1'b0;
  assign lce_data_resp_o[368] = 1'b0;
  assign lce_data_resp_o[369] = 1'b0;
  assign lce_data_resp_o[370] = 1'b0;
  assign lce_data_resp_o[371] = 1'b0;
  assign lce_data_resp_o[372] = 1'b0;
  assign lce_data_resp_o[373] = 1'b0;
  assign lce_data_resp_o[374] = 1'b0;
  assign lce_data_resp_o[375] = 1'b0;
  assign lce_data_resp_o[376] = 1'b0;
  assign lce_data_resp_o[377] = 1'b0;
  assign lce_data_resp_o[378] = 1'b0;
  assign lce_data_resp_o[379] = 1'b0;
  assign lce_data_resp_o[380] = 1'b0;
  assign lce_data_resp_o[381] = 1'b0;
  assign lce_data_resp_o[382] = 1'b0;
  assign lce_data_resp_o[383] = 1'b0;
  assign lce_data_resp_o[384] = 1'b0;
  assign lce_data_resp_o[385] = 1'b0;
  assign lce_data_resp_o[386] = 1'b0;
  assign lce_data_resp_o[387] = 1'b0;
  assign lce_data_resp_o[388] = 1'b0;
  assign lce_data_resp_o[389] = 1'b0;
  assign lce_data_resp_o[390] = 1'b0;
  assign lce_data_resp_o[391] = 1'b0;
  assign lce_data_resp_o[392] = 1'b0;
  assign lce_data_resp_o[393] = 1'b0;
  assign lce_data_resp_o[394] = 1'b0;
  assign lce_data_resp_o[395] = 1'b0;
  assign lce_data_resp_o[396] = 1'b0;
  assign lce_data_resp_o[397] = 1'b0;
  assign lce_data_resp_o[398] = 1'b0;
  assign lce_data_resp_o[399] = 1'b0;
  assign lce_data_resp_o[400] = 1'b0;
  assign lce_data_resp_o[401] = 1'b0;
  assign lce_data_resp_o[402] = 1'b0;
  assign lce_data_resp_o[403] = 1'b0;
  assign lce_data_resp_o[404] = 1'b0;
  assign lce_data_resp_o[405] = 1'b0;
  assign lce_data_resp_o[406] = 1'b0;
  assign lce_data_resp_o[407] = 1'b0;
  assign lce_data_resp_o[408] = 1'b0;
  assign lce_data_resp_o[409] = 1'b0;
  assign lce_data_resp_o[410] = 1'b0;
  assign lce_data_resp_o[411] = 1'b0;
  assign lce_data_resp_o[412] = 1'b0;
  assign lce_data_resp_o[413] = 1'b0;
  assign lce_data_resp_o[414] = 1'b0;
  assign lce_data_resp_o[415] = 1'b0;
  assign lce_data_resp_o[416] = 1'b0;
  assign lce_data_resp_o[417] = 1'b0;
  assign lce_data_resp_o[418] = 1'b0;
  assign lce_data_resp_o[419] = 1'b0;
  assign lce_data_resp_o[420] = 1'b0;
  assign lce_data_resp_o[421] = 1'b0;
  assign lce_data_resp_o[422] = 1'b0;
  assign lce_data_resp_o[423] = 1'b0;
  assign lce_data_resp_o[424] = 1'b0;
  assign lce_data_resp_o[425] = 1'b0;
  assign lce_data_resp_o[426] = 1'b0;
  assign lce_data_resp_o[427] = 1'b0;
  assign lce_data_resp_o[428] = 1'b0;
  assign lce_data_resp_o[429] = 1'b0;
  assign lce_data_resp_o[430] = 1'b0;
  assign lce_data_resp_o[431] = 1'b0;
  assign lce_data_resp_o[432] = 1'b0;
  assign lce_data_resp_o[433] = 1'b0;
  assign lce_data_resp_o[434] = 1'b0;
  assign lce_data_resp_o[435] = 1'b0;
  assign lce_data_resp_o[436] = 1'b0;
  assign lce_data_resp_o[437] = 1'b0;
  assign lce_data_resp_o[438] = 1'b0;
  assign lce_data_resp_o[439] = 1'b0;
  assign lce_data_resp_o[440] = 1'b0;
  assign lce_data_resp_o[441] = 1'b0;
  assign lce_data_resp_o[442] = 1'b0;
  assign lce_data_resp_o[443] = 1'b0;
  assign lce_data_resp_o[444] = 1'b0;
  assign lce_data_resp_o[445] = 1'b0;
  assign lce_data_resp_o[446] = 1'b0;
  assign lce_data_resp_o[447] = 1'b0;
  assign lce_data_resp_o[448] = 1'b0;
  assign lce_data_resp_o[449] = 1'b0;
  assign lce_data_resp_o[450] = 1'b0;
  assign lce_data_resp_o[451] = 1'b0;
  assign lce_data_resp_o[452] = 1'b0;
  assign lce_data_resp_o[453] = 1'b0;
  assign lce_data_resp_o[454] = 1'b0;
  assign lce_data_resp_o[455] = 1'b0;
  assign lce_data_resp_o[456] = 1'b0;
  assign lce_data_resp_o[457] = 1'b0;
  assign lce_data_resp_o[458] = 1'b0;
  assign lce_data_resp_o[459] = 1'b0;
  assign lce_data_resp_o[460] = 1'b0;
  assign lce_data_resp_o[461] = 1'b0;
  assign lce_data_resp_o[462] = 1'b0;
  assign lce_data_resp_o[463] = 1'b0;
  assign lce_data_resp_o[464] = 1'b0;
  assign lce_data_resp_o[465] = 1'b0;
  assign lce_data_resp_o[466] = 1'b0;
  assign lce_data_resp_o[467] = 1'b0;
  assign lce_data_resp_o[468] = 1'b0;
  assign lce_data_resp_o[469] = 1'b0;
  assign lce_data_resp_o[470] = 1'b0;
  assign lce_data_resp_o[471] = 1'b0;
  assign lce_data_resp_o[472] = 1'b0;
  assign lce_data_resp_o[473] = 1'b0;
  assign lce_data_resp_o[474] = 1'b0;
  assign lce_data_resp_o[475] = 1'b0;
  assign lce_data_resp_o[476] = 1'b0;
  assign lce_data_resp_o[477] = 1'b0;
  assign lce_data_resp_o[478] = 1'b0;
  assign lce_data_resp_o[479] = 1'b0;
  assign lce_data_resp_o[480] = 1'b0;
  assign lce_data_resp_o[481] = 1'b0;
  assign lce_data_resp_o[482] = 1'b0;
  assign lce_data_resp_o[483] = 1'b0;
  assign lce_data_resp_o[484] = 1'b0;
  assign lce_data_resp_o[485] = 1'b0;
  assign lce_data_resp_o[486] = 1'b0;
  assign lce_data_resp_o[487] = 1'b0;
  assign lce_data_resp_o[488] = 1'b0;
  assign lce_data_resp_o[489] = 1'b0;
  assign lce_data_resp_o[490] = 1'b0;
  assign lce_data_resp_o[491] = 1'b0;
  assign lce_data_resp_o[492] = 1'b0;
  assign lce_data_resp_o[493] = 1'b0;
  assign lce_data_resp_o[494] = 1'b0;
  assign lce_data_resp_o[495] = 1'b0;
  assign lce_data_resp_o[496] = 1'b0;
  assign lce_data_resp_o[497] = 1'b0;
  assign lce_data_resp_o[498] = 1'b0;
  assign lce_data_resp_o[499] = 1'b0;
  assign lce_data_resp_o[500] = 1'b0;
  assign lce_data_resp_o[501] = 1'b0;
  assign lce_data_resp_o[502] = 1'b0;
  assign lce_data_resp_o[503] = 1'b0;
  assign lce_data_resp_o[504] = 1'b0;
  assign lce_data_resp_o[505] = 1'b0;
  assign lce_data_resp_o[506] = 1'b0;
  assign lce_data_resp_o[507] = 1'b0;
  assign lce_data_resp_o[508] = 1'b0;
  assign lce_data_resp_o[509] = 1'b0;
  assign lce_data_resp_o[510] = 1'b0;
  assign lce_data_resp_o[511] = 1'b0;
  assign lce_resp_o[23] = 1'b0;
  assign N24 = state_r[1] | N23;
  assign N27 = N26 | state_r[0];
  assign N29 = N26 & N23;
  assign lce_ready_o = state_r[0] | state_r[1];
  assign N1378 = ~lce_cmd_i[31];
  assign N1379 = lce_cmd_i[32] | lce_cmd_i[33];
  assign N1380 = N1378 | N1379;
  assign N1381 = ~N1380;
  assign N1382 = ~lce_cmd_i[33];
  assign N1383 = ~lce_cmd_i[32];
  assign N1384 = N1383 | N1382;
  assign N1385 = lce_cmd_i[31] | N1384;
  assign N1386 = ~N1385;
  assign N1387 = syn_ack_cnt_r[4] | syn_ack_cnt_r[5];
  assign N1388 = syn_ack_cnt_r[3] | N1387;
  assign N1389 = syn_ack_cnt_r[2] | N1388;
  assign N1390 = syn_ack_cnt_r[1] | N1389;
  assign N1391 = syn_ack_cnt_r[0] | N1390;
  assign N1392 = ~N1391;
  assign N1393 = lce_cmd_i[32] | N1382;
  assign N1394 = N1378 | N1393;
  assign N1395 = ~N1394;
  assign N1396 = lce_cmd_i[31] | N1393;
  assign N1397 = ~N1396;
  assign N1398 = N1378 | N1400;
  assign N1399 = ~N1398;
  assign N1400 = N1383 | lce_cmd_i[33];
  assign N1401 = lce_cmd_i[31] | N1400;
  assign N1402 = ~N1401;
  assign N1403 = lce_cmd_i[31] | N1379;
  assign N1404 = ~N1403;
  assign { N673, N672, N671, N670, N669, N668 } = syn_ack_cnt_r + 1'b1;
  assign N38 = (N0)? 1'b0 : 
               (N1)? lce_cmd_v_i : 1'b0;
  assign N0 = flag_invalidate_r;
  assign N1 = N37;
  assign N41 = (N2)? 1'b0 : 
               (N700)? 1'b1 : 
               (N40)? tag_mem_pkt_yumi_i : 1'b0;
  assign N2 = lce_resp_yumi_i;
  assign N44 = (N3)? 1'b0 : 
               (N4)? N43 : 1'b0;
  assign N3 = flag_updated_lru_r;
  assign N4 = N42;
  assign N47 = (N2)? 1'b0 : 
               (N702)? 1'b1 : 
               (N46)? metadata_mem_pkt_yumi_i : 1'b0;
  assign { N57, N56, N55, N54, N53, N52, N51, N50, N49 } = (N5)? { lce_cmd_i[20:15], lce_cmd_i[8:6] } : 
                                                           (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                           (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                           (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                           (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                           (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N5 = N1402;
  assign N6 = N1401;
  assign N7 = 1'b0;
  assign N58 = (N5)? lce_cmd_v_i : 
               (N6)? 1'b0 : 
               (N7)? 1'b0 : 
               (N7)? 1'b0 : 
               (N7)? 1'b0 : 
               (N7)? 1'b0 : 1'b0;
  assign { N60, N59 } = (N5)? { data_mem_pkt_yumi_i, N35 } : 
                        (N6)? state_r : 1'b0;
  assign { N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                           (N8)? { lce_cmd_i[34:34], id_i[0:0], 1'b1, lce_cmd_i[30:9] } : 
                                                                                                                                           (N61)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                           (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                           (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                           (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = N1399;
  assign N87 = (N5)? 1'b0 : 
               (N8)? lce_cmd_v_i : 
               (N61)? 1'b0 : 
               (N7)? 1'b0 : 
               (N7)? 1'b0 : 
               (N7)? 1'b0 : 1'b0;
  assign N88 = (N5)? 1'b0 : 
               (N8)? N36 : 
               (N9)? tag_mem_pkt_yumi_i : 
               (N10)? tag_mem_pkt_yumi_i : 
               (N11)? lce_resp_yumi_i : 
               (N34)? 1'b0 : 1'b0;
  assign N9 = N1397;
  assign N10 = N1395;
  assign N11 = N1386;
  assign { N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                  (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                  (N9)? { lce_cmd_i[5:4], lce_cmd_i[30:21], 1'b1 } : 
                                                                                  (N10)? { lce_cmd_i[5:4], lce_cmd_i[30:21], 1'b1 } : 
                                                                                  (N89)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                  (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N111, N110, N109, N108, N107, N106, N105, N104, N103 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                    (N9)? { lce_cmd_i[20:15], lce_cmd_i[8:6] } : 
                                                                    (N10)? { lce_cmd_i[20:15], lce_cmd_i[8:6] } : 
                                                                    (N11)? { lce_cmd_i[20:15], lce_cmd_i[8:6] } : 
                                                                    (N34)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N112 = (N5)? 1'b0 : 
                (N8)? 1'b0 : 
                (N9)? lce_cmd_v_i : 
                (N10)? lce_cmd_v_i : 
                (N11)? N38 : 
                (N34)? 1'b0 : 1'b0;
  assign N114 = (N5)? 1'b0 : 
                (N8)? 1'b0 : 
                (N9)? tag_mem_pkt_yumi_i : 
                (N113)? 1'b0 : 
                (N7)? 1'b0 : 
                (N7)? 1'b0 : 1'b0;
  assign N115 = (N5)? 1'b0 : 
                (N8)? 1'b0 : 
                (N9)? 1'b0 : 
                (N10)? tag_mem_pkt_yumi_i : 
                (N89)? 1'b0 : 
                (N7)? 1'b0 : 1'b0;
  assign N116 = (N11)? N41 : 
                (N34)? flag_invalidate_r : 1'b0;
  assign { N126, N125, N124, N123, N122, N121, N120, N119, N118, N117 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N11)? { lce_cmd_i[20:15], lce_cmd_i[8:6], 1'b1 } : 
                                                                          (N34)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N127 = (N5)? 1'b0 : 
                (N8)? 1'b0 : 
                (N9)? 1'b0 : 
                (N10)? 1'b0 : 
                (N11)? N44 : 
                (N34)? 1'b0 : 1'b0;
  assign N128 = (N11)? N47 : 
                (N34)? flag_updated_lru_r : 1'b0;
  assign { N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                          (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                          (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                          (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                          (N11)? { lce_cmd_i[34:34], id_i[0:0], lce_cmd_i[30:21], lce_cmd_i[14:9] } : 
                                                                                                                          (N34)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N147 = (N5)? 1'b0 : 
                (N8)? 1'b0 : 
                (N9)? 1'b0 : 
                (N10)? 1'b0 : 
                (N11)? N48 : 
                (N34)? 1'b0 : 1'b0;
  assign { N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150 } = (N12)? data_r : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N13)? data_mem_data_i : 1'b0;
  assign N12 = flag_data_buffered_r;
  assign N13 = N149;
  assign { N677, N676 } = (N14)? { 1'b0, 1'b1 } : 
                          (N675)? state_r : 1'b0;
  assign N14 = N674;
  assign { N683, N682, N681, N680, N679, N678 } = (N15)? lce_cmd_i[20:15] : 
                                                  (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                  (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = N1381;
  assign N16 = N1380;
  assign N684 = (N15)? lce_cmd_v_i : 
                (N16)? 1'b0 : 
                (N7)? 1'b0 : 1'b0;
  assign N685 = (N15)? tag_mem_pkt_yumi_i : 
                (N17)? lce_resp_yumi_i : 
                (N664)? 1'b0 : 1'b0;
  assign N17 = N1404;
  assign { N687, N686 } = (N15)? { 1'b0, 1'b0 } : 
                          (N17)? { lce_cmd_i[34:34], id_i[0:0] } : 
                          (N664)? { 1'b0, 1'b0 } : 1'b0;
  assign N688 = (N15)? 1'b0 : 
                (N17)? lce_cmd_v_i : 
                (N664)? 1'b0 : 1'b0;
  assign { N694, N693, N692, N691, N690, N689 } = (N17)? { N673, N672, N671, N670, N669, N668 } : 
                                                  (N664)? syn_ack_cnt_r : 1'b0;
  assign { N696, N695 } = (N17)? { N677, N676 } : 
                          (N664)? state_r : 1'b0;
  assign lce_resp_v_o = (N18)? N147 : 
                        (N19)? 1'b0 : 
                        (N20)? N688 : 
                        (N699)? 1'b0 : 1'b0;
  assign N18 = N25;
  assign N19 = N28;
  assign N20 = N29;
  assign data_mem_pkt_o[73:65] = (N18)? { N57, N56, N55, N54, N53, N52, N51, N50, N49 } : 
                                 (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                 (N699)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign data_mem_pkt_v_o = (N18)? N58 : 
                            (N19)? 1'b0 : 
                            (N20)? 1'b0 : 
                            (N699)? 1'b0 : 1'b0;
  assign state_n = (N18)? { N60, N59 } : 
                   (N19)? { N148, lce_tr_resp_ready_i } : 
                   (N20)? { N696, N695 } : 1'b0;
  assign lce_data_resp_o[536:512] = (N18)? { N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62 } : 
                                    (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                    (N699)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_data_resp_v_o = (N18)? N87 : 
                             (N19)? 1'b0 : 
                             (N20)? 1'b0 : 
                             (N699)? 1'b0 : 1'b0;
  assign lce_cmd_yumi_o = (N18)? N88 : 
                          (N19)? lce_tr_resp_ready_i : 
                          (N20)? N685 : 
                          (N699)? 1'b0 : 1'b0;
  assign tag_mem_pkt_o = (N18)? { N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N1386 } : 
                         (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N20)? { N683, N682, N681, N680, N679, N678, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N699)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_mem_pkt_v_o = (N18)? N112 : 
                           (N19)? 1'b0 : 
                           (N20)? N684 : 
                           (N699)? 1'b0 : 1'b0;
  assign tag_set_o = (N18)? N114 : 
                     (N19)? 1'b0 : 
                     (N20)? 1'b0 : 
                     (N699)? 1'b0 : 1'b0;
  assign tag_set_wakeup_o = (N18)? N115 : 
                            (N19)? 1'b0 : 
                            (N20)? 1'b0 : 
                            (N699)? 1'b0 : 1'b0;
  assign metadata_mem_pkt_o = (N18)? { N126, N125, N124, N123, N122, N121, N120, N119, N118, N117 } : 
                              (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N20)? { N683, N682, N681, N680, N679, N678, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N699)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign metadata_mem_pkt_v_o = (N18)? N127 : 
                                (N19)? 1'b0 : 
                                (N20)? N684 : 
                                (N699)? 1'b0 : 1'b0;
  assign { lce_resp_o[25:24], lce_resp_o[22:0] } = (N18)? { N146, N145, N117, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N126, N125, N124, N123, N122, N121, N134, N133, N132, N131, N130, N129 } : 
                                                   (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                   (N20)? { N687, N686, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                   (N699)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_tr_resp_o = (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N19)? { lce_cmd_i[3:3], id_i[0:0], lce_cmd_i[2:0], lce_cmd_i[30:9], N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150 } : 
                         (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                         (N699)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_tr_resp_v_o = (N18)? 1'b0 : 
                           (N19)? 1'b1 : 
                           (N20)? 1'b0 : 
                           (N699)? 1'b0 : 1'b0;
  assign { N705, N704 } = (N21)? { 1'b0, 1'b0 } : 
                          (N22)? state_n : 1'b0;
  assign N21 = reset_i;
  assign N22 = N703;
  assign { N711, N710, N709, N708, N707, N706 } = (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                  (N22)? { N694, N693, N692, N691, N690, N689 } : 1'b0;
  assign { N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712 } = (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N22)? data_mem_data_i : 1'b0;
  assign N1224 = (N21)? 1'b0 : 
                 (N22)? N148 : 1'b0;
  assign N1225 = (N21)? 1'b0 : 
                 (N22)? N116 : 1'b0;
  assign N1226 = (N21)? 1'b0 : 
                 (N22)? N128 : 1'b0;
  assign N23 = ~state_r[0];
  assign N25 = ~N24;
  assign N26 = ~state_r[1];
  assign N28 = ~N27;
  assign N30 = N1399 | N1402;
  assign N31 = N1397 | N30;
  assign N32 = N1395 | N31;
  assign N33 = N1386 | N32;
  assign N34 = ~N33;
  assign N35 = ~data_mem_pkt_yumi_i;
  assign N36 = lce_data_resp_ready_i & lce_cmd_v_i;
  assign N37 = ~flag_invalidate_r;
  assign N39 = flag_invalidate_r | lce_resp_yumi_i;
  assign N40 = ~N39;
  assign N42 = ~flag_updated_lru_r;
  assign N43 = flag_invalidate_r | tag_mem_pkt_yumi_i;
  assign N45 = flag_updated_lru_r | lce_resp_yumi_i;
  assign N46 = ~N45;
  assign N48 = N1405 & N1406;
  assign N1405 = flag_invalidate_r | tag_mem_pkt_yumi_i;
  assign N1406 = flag_updated_lru_r | metadata_mem_pkt_yumi_i;
  assign N61 = ~N30;
  assign N89 = ~N32;
  assign N113 = ~N31;
  assign N148 = ~lce_tr_resp_ready_i;
  assign N149 = ~flag_data_buffered_r;
  assign N662 = N29;
  assign N663 = N1404 | N1381;
  assign N664 = ~N663;
  assign N665 = N662 & N1404;
  assign N666 = lce_cmd_v_i & lce_resp_yumi_i;
  assign N667 = ~N666;
  assign N674 = N1407 & lce_resp_yumi_i;
  assign N1407 = N1392 & lce_cmd_v_i;
  assign N675 = ~N674;
  assign N697 = N28 | N25;
  assign N698 = N29 | N697;
  assign N699 = ~N698;
  assign N700 = flag_invalidate_r & N701;
  assign N701 = ~lce_resp_yumi_i;
  assign N702 = flag_updated_lru_r & N701;
  assign N703 = ~reset_i;
  assign N1227 = N25 & N703;
  assign N1228 = N1402 & N1227;
  assign N1229 = N25 & N703;
  assign N1230 = N1399 & N1229;
  assign N1231 = N1228 | N1230;
  assign N1232 = N25 & N703;
  assign N1233 = N1397 & N1232;
  assign N1234 = N1231 | N1233;
  assign N1235 = N25 & N703;
  assign N1236 = N1395 & N1235;
  assign N1237 = N1234 | N1236;
  assign N1238 = N28 & N703;
  assign N1239 = N1237 | N1238;
  assign N1240 = N29 & N703;
  assign N1241 = N1239 | N1240;
  assign N1242 = N699 & N703;
  assign N1243 = N1241 | N1242;
  assign N1244 = ~N1243;
  assign N1245 = N29 & N703;
  assign N1246 = N1381 & N1245;
  assign N1247 = N699 & N703;
  assign N1248 = N1246 | N1247;
  assign N1249 = ~N1248;
  assign N1250 = N29 & N703;
  assign N1251 = N1381 & N1250;
  assign N1252 = N699 & N703;
  assign N1253 = N1251 | N1252;
  assign N1254 = ~N1253;
  assign N1255 = N25 & N703;
  assign N1256 = N28 & N703;
  assign N1257 = N1255 | N1256;
  assign N1258 = N29 & N703;
  assign N1259 = N1381 & N1258;
  assign N1260 = N1257 | N1259;
  assign N1261 = N29 & N703;
  assign N1262 = N1404 & N1261;
  assign N1263 = N667 & N1262;
  assign N1264 = N1260 | N1263;
  assign N1265 = N699 & N703;
  assign N1266 = N1264 | N1265;
  assign N1267 = ~N1266;
  assign N1268 = N25 & N703;
  assign N1269 = N28 & N703;
  assign N1270 = N1268 | N1269;
  assign N1271 = N29 & N703;
  assign N1272 = N1381 & N1271;
  assign N1273 = N1270 | N1272;
  assign N1274 = N1404 & N1271;
  assign N1275 = N667 & N1274;
  assign N1276 = N1273 | N1275;
  assign N1277 = N699 & N703;
  assign N1278 = N1276 | N1277;
  assign N1279 = ~N1278;
  assign N1280 = N28 & N703;
  assign N1281 = N1268 | N1280;
  assign N1282 = N1281 | N1272;
  assign N1283 = N1282 | N1275;
  assign N1284 = N699 & N703;
  assign N1285 = N1283 | N1284;
  assign N1286 = ~N1285;
  assign N1287 = N28 & N703;
  assign N1288 = N1268 | N1287;
  assign N1289 = N1288 | N1272;
  assign N1290 = N1289 | N1275;
  assign N1291 = N1290 | N1284;
  assign N1292 = ~N1291;
  assign N1293 = N28 & N703;
  assign N1294 = N1268 | N1293;
  assign N1295 = N1294 | N1272;
  assign N1296 = N1295 | N1275;
  assign N1297 = N1296 | N1284;
  assign N1298 = ~N1297;
  assign N1299 = flag_data_buffered_r & N1293;
  assign N1300 = N1268 | N1299;
  assign N1301 = N1300 | N1271;
  assign N1302 = N1301 | N1284;
  assign N1303 = ~N1302;
  assign N1304 = flag_data_buffered_r & N1287;
  assign N1305 = N1268 | N1304;
  assign N1306 = N1305 | N1271;
  assign N1307 = N1306 | N1284;
  assign N1308 = ~N1307;
  assign N1309 = N1305 | N1261;
  assign N1310 = N1309 | N1277;
  assign N1311 = ~N1310;
  assign N1312 = N1255 | N1304;
  assign N1313 = N1312 | N1261;
  assign N1314 = N1313 | N1277;
  assign N1315 = ~N1314;
  assign N1316 = flag_data_buffered_r & N1280;
  assign N1317 = N1255 | N1316;
  assign N1318 = N1317 | N1261;
  assign N1319 = N1318 | N1277;
  assign N1320 = ~N1319;
  assign N1321 = N1317 | N1258;
  assign N1322 = N1321 | N1265;
  assign N1323 = ~N1322;
  assign N1324 = N1235 | N1316;
  assign N1325 = N1324 | N1258;
  assign N1326 = N1325 | N1265;
  assign N1327 = ~N1326;
  assign N1328 = flag_data_buffered_r & N1269;
  assign N1329 = N1235 | N1328;
  assign N1330 = N1329 | N1258;
  assign N1331 = N1330 | N1265;
  assign N1332 = ~N1331;
  assign N1333 = N1329 | N1250;
  assign N1334 = N1333 | N1252;
  assign N1335 = ~N1334;
  assign N1336 = N1232 | N1328;
  assign N1337 = N1336 | N1250;
  assign N1338 = N1337 | N1252;
  assign N1339 = ~N1338;
  assign N1340 = flag_data_buffered_r & N1256;
  assign N1341 = N1232 | N1340;
  assign N1342 = N1341 | N1250;
  assign N1343 = N1342 | N1252;
  assign N1344 = ~N1343;
  assign N1345 = N1341 | N1245;
  assign N1346 = N1345 | N1247;
  assign N1347 = ~N1346;
  assign N1348 = N1229 | N1340;
  assign N1349 = N1348 | N1245;
  assign N1350 = N1349 | N1247;
  assign N1351 = ~N1350;
  assign N1352 = flag_data_buffered_r & N1238;
  assign N1353 = N1229 | N1352;
  assign N1354 = N1353 | N1245;
  assign N1355 = N1354 | N1247;
  assign N1356 = ~N1355;
  assign N1357 = N1353 | N1240;
  assign N1358 = N1357 | N1242;
  assign N1359 = ~N1358;
  assign N1360 = N1227 | N1352;
  assign N1361 = N1360 | N1240;
  assign N1362 = N1361 | N1242;
  assign N1363 = ~N1362;
  assign N1364 = N1227 | N1240;
  assign N1365 = N1364 | N1242;
  assign N1366 = ~N1365;
  assign N1367 = N1399 & N1227;
  assign N1368 = N1228 | N1367;
  assign N1369 = N1397 & N1227;
  assign N1370 = N1368 | N1369;
  assign N1371 = N1395 & N1227;
  assign N1372 = N1370 | N1371;
  assign N1373 = N1372 | N1238;
  assign N1374 = N1373 | N1240;
  assign N1375 = N1374 | N1242;
  assign N1376 = ~N1375;

  always @(posedge clk_i) begin
    if(N1244) begin
      flag_updated_lru_r <= N1226;
    end 
    if(N1249) begin
      { state_r[1:1] } <= { N705 };
    end 
    if(N1254) begin
      { state_r[0:0] } <= { N704 };
    end 
    if(N1267) begin
      { syn_ack_cnt_r[5:5] } <= { N711 };
    end 
    if(N1279) begin
      { syn_ack_cnt_r[4:4] } <= { N710 };
    end 
    if(N1286) begin
      { syn_ack_cnt_r[3:3] } <= { N709 };
    end 
    if(N1292) begin
      { syn_ack_cnt_r[2:2] } <= { N708 };
    end 
    if(N1298) begin
      { syn_ack_cnt_r[1:0] } <= { N707, N706 };
    end 
    if(N1303) begin
      { data_r[511:494] } <= { N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206 };
    end 
    if(N1308) begin
      { data_r[493:493] } <= { N1205 };
    end 
    if(N1311) begin
      { data_r[492:490] } <= { N1204, N1203, N1202 };
    end 
    if(N1315) begin
      { data_r[489:395] } <= { N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107 };
    end 
    if(N1320) begin
      { data_r[394:394] } <= { N1106 };
    end 
    if(N1323) begin
      { data_r[393:391] } <= { N1105, N1104, N1103 };
    end 
    if(N1327) begin
      { data_r[390:296] } <= { N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008 };
    end 
    if(N1332) begin
      { data_r[295:295] } <= { N1007 };
    end 
    if(N1335) begin
      { data_r[294:292] } <= { N1006, N1005, N1004 };
    end 
    if(N1339) begin
      { data_r[291:197] } <= { N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909 };
    end 
    if(N1344) begin
      { data_r[196:196] } <= { N908 };
    end 
    if(N1347) begin
      { data_r[195:193] } <= { N907, N906, N905 };
    end 
    if(N1351) begin
      { data_r[192:98] } <= { N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810 };
    end 
    if(N1356) begin
      { data_r[97:97] } <= { N809 };
    end 
    if(N1359) begin
      { data_r[96:94] } <= { N808, N807, N806 };
    end 
    if(N1363) begin
      { data_r[93:0] } <= { N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712 };
    end 
    if(N1366) begin
      flag_data_buffered_r <= N1224;
    end 
    if(N1376) begin
      flag_invalidate_r <= N1225;
    end 
  end


endmodule



// module bsg_mem_p540
// (
//   w_clk_i,
//   w_reset_i,
//   w_v_i,
//   w_addr_i,
//   w_data_i,
//   r_v_i,
//   r_addr_i,
//   r_data_o
// );

//   input [0:0] w_addr_i;
//   input [539:0] w_data_i;
//   input [0:0] r_addr_i;
//   output [539:0] r_data_o;
//   input w_clk_i;
//   input w_reset_i;
//   input w_v_i;
//   input r_v_i;
//   wire [539:0] r_data_o;
//   wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;
//   reg [1079:0] mem;
//   assign r_data_o[539] = (N3)? mem[539] : 
//                          (N0)? mem[1079] : 1'b0;
//   assign N0 = r_addr_i[0];
//   assign r_data_o[538] = (N3)? mem[538] : 
//                          (N0)? mem[1078] : 1'b0;
//   assign r_data_o[537] = (N3)? mem[537] : 
//                          (N0)? mem[1077] : 1'b0;
//   assign r_data_o[536] = (N3)? mem[536] : 
//                          (N0)? mem[1076] : 1'b0;
//   assign r_data_o[535] = (N3)? mem[535] : 
//                          (N0)? mem[1075] : 1'b0;
//   assign r_data_o[534] = (N3)? mem[534] : 
//                          (N0)? mem[1074] : 1'b0;
//   assign r_data_o[533] = (N3)? mem[533] : 
//                          (N0)? mem[1073] : 1'b0;
//   assign r_data_o[532] = (N3)? mem[532] : 
//                          (N0)? mem[1072] : 1'b0;
//   assign r_data_o[531] = (N3)? mem[531] : 
//                          (N0)? mem[1071] : 1'b0;
//   assign r_data_o[530] = (N3)? mem[530] : 
//                          (N0)? mem[1070] : 1'b0;
//   assign r_data_o[529] = (N3)? mem[529] : 
//                          (N0)? mem[1069] : 1'b0;
//   assign r_data_o[528] = (N3)? mem[528] : 
//                          (N0)? mem[1068] : 1'b0;
//   assign r_data_o[527] = (N3)? mem[527] : 
//                          (N0)? mem[1067] : 1'b0;
//   assign r_data_o[526] = (N3)? mem[526] : 
//                          (N0)? mem[1066] : 1'b0;
//   assign r_data_o[525] = (N3)? mem[525] : 
//                          (N0)? mem[1065] : 1'b0;
//   assign r_data_o[524] = (N3)? mem[524] : 
//                          (N0)? mem[1064] : 1'b0;
//   assign r_data_o[523] = (N3)? mem[523] : 
//                          (N0)? mem[1063] : 1'b0;
//   assign r_data_o[522] = (N3)? mem[522] : 
//                          (N0)? mem[1062] : 1'b0;
//   assign r_data_o[521] = (N3)? mem[521] : 
//                          (N0)? mem[1061] : 1'b0;
//   assign r_data_o[520] = (N3)? mem[520] : 
//                          (N0)? mem[1060] : 1'b0;
//   assign r_data_o[519] = (N3)? mem[519] : 
//                          (N0)? mem[1059] : 1'b0;
//   assign r_data_o[518] = (N3)? mem[518] : 
//                          (N0)? mem[1058] : 1'b0;
//   assign r_data_o[517] = (N3)? mem[517] : 
//                          (N0)? mem[1057] : 1'b0;
//   assign r_data_o[516] = (N3)? mem[516] : 
//                          (N0)? mem[1056] : 1'b0;
//   assign r_data_o[515] = (N3)? mem[515] : 
//                          (N0)? mem[1055] : 1'b0;
//   assign r_data_o[514] = (N3)? mem[514] : 
//                          (N0)? mem[1054] : 1'b0;
//   assign r_data_o[513] = (N3)? mem[513] : 
//                          (N0)? mem[1053] : 1'b0;
//   assign r_data_o[512] = (N3)? mem[512] : 
//                          (N0)? mem[1052] : 1'b0;
//   assign r_data_o[511] = (N3)? mem[511] : 
//                          (N0)? mem[1051] : 1'b0;
//   assign r_data_o[510] = (N3)? mem[510] : 
//                          (N0)? mem[1050] : 1'b0;
//   assign r_data_o[509] = (N3)? mem[509] : 
//                          (N0)? mem[1049] : 1'b0;
//   assign r_data_o[508] = (N3)? mem[508] : 
//                          (N0)? mem[1048] : 1'b0;
//   assign r_data_o[507] = (N3)? mem[507] : 
//                          (N0)? mem[1047] : 1'b0;
//   assign r_data_o[506] = (N3)? mem[506] : 
//                          (N0)? mem[1046] : 1'b0;
//   assign r_data_o[505] = (N3)? mem[505] : 
//                          (N0)? mem[1045] : 1'b0;
//   assign r_data_o[504] = (N3)? mem[504] : 
//                          (N0)? mem[1044] : 1'b0;
//   assign r_data_o[503] = (N3)? mem[503] : 
//                          (N0)? mem[1043] : 1'b0;
//   assign r_data_o[502] = (N3)? mem[502] : 
//                          (N0)? mem[1042] : 1'b0;
//   assign r_data_o[501] = (N3)? mem[501] : 
//                          (N0)? mem[1041] : 1'b0;
//   assign r_data_o[500] = (N3)? mem[500] : 
//                          (N0)? mem[1040] : 1'b0;
//   assign r_data_o[499] = (N3)? mem[499] : 
//                          (N0)? mem[1039] : 1'b0;
//   assign r_data_o[498] = (N3)? mem[498] : 
//                          (N0)? mem[1038] : 1'b0;
//   assign r_data_o[497] = (N3)? mem[497] : 
//                          (N0)? mem[1037] : 1'b0;
//   assign r_data_o[496] = (N3)? mem[496] : 
//                          (N0)? mem[1036] : 1'b0;
//   assign r_data_o[495] = (N3)? mem[495] : 
//                          (N0)? mem[1035] : 1'b0;
//   assign r_data_o[494] = (N3)? mem[494] : 
//                          (N0)? mem[1034] : 1'b0;
//   assign r_data_o[493] = (N3)? mem[493] : 
//                          (N0)? mem[1033] : 1'b0;
//   assign r_data_o[492] = (N3)? mem[492] : 
//                          (N0)? mem[1032] : 1'b0;
//   assign r_data_o[491] = (N3)? mem[491] : 
//                          (N0)? mem[1031] : 1'b0;
//   assign r_data_o[490] = (N3)? mem[490] : 
//                          (N0)? mem[1030] : 1'b0;
//   assign r_data_o[489] = (N3)? mem[489] : 
//                          (N0)? mem[1029] : 1'b0;
//   assign r_data_o[488] = (N3)? mem[488] : 
//                          (N0)? mem[1028] : 1'b0;
//   assign r_data_o[487] = (N3)? mem[487] : 
//                          (N0)? mem[1027] : 1'b0;
//   assign r_data_o[486] = (N3)? mem[486] : 
//                          (N0)? mem[1026] : 1'b0;
//   assign r_data_o[485] = (N3)? mem[485] : 
//                          (N0)? mem[1025] : 1'b0;
//   assign r_data_o[484] = (N3)? mem[484] : 
//                          (N0)? mem[1024] : 1'b0;
//   assign r_data_o[483] = (N3)? mem[483] : 
//                          (N0)? mem[1023] : 1'b0;
//   assign r_data_o[482] = (N3)? mem[482] : 
//                          (N0)? mem[1022] : 1'b0;
//   assign r_data_o[481] = (N3)? mem[481] : 
//                          (N0)? mem[1021] : 1'b0;
//   assign r_data_o[480] = (N3)? mem[480] : 
//                          (N0)? mem[1020] : 1'b0;
//   assign r_data_o[479] = (N3)? mem[479] : 
//                          (N0)? mem[1019] : 1'b0;
//   assign r_data_o[478] = (N3)? mem[478] : 
//                          (N0)? mem[1018] : 1'b0;
//   assign r_data_o[477] = (N3)? mem[477] : 
//                          (N0)? mem[1017] : 1'b0;
//   assign r_data_o[476] = (N3)? mem[476] : 
//                          (N0)? mem[1016] : 1'b0;
//   assign r_data_o[475] = (N3)? mem[475] : 
//                          (N0)? mem[1015] : 1'b0;
//   assign r_data_o[474] = (N3)? mem[474] : 
//                          (N0)? mem[1014] : 1'b0;
//   assign r_data_o[473] = (N3)? mem[473] : 
//                          (N0)? mem[1013] : 1'b0;
//   assign r_data_o[472] = (N3)? mem[472] : 
//                          (N0)? mem[1012] : 1'b0;
//   assign r_data_o[471] = (N3)? mem[471] : 
//                          (N0)? mem[1011] : 1'b0;
//   assign r_data_o[470] = (N3)? mem[470] : 
//                          (N0)? mem[1010] : 1'b0;
//   assign r_data_o[469] = (N3)? mem[469] : 
//                          (N0)? mem[1009] : 1'b0;
//   assign r_data_o[468] = (N3)? mem[468] : 
//                          (N0)? mem[1008] : 1'b0;
//   assign r_data_o[467] = (N3)? mem[467] : 
//                          (N0)? mem[1007] : 1'b0;
//   assign r_data_o[466] = (N3)? mem[466] : 
//                          (N0)? mem[1006] : 1'b0;
//   assign r_data_o[465] = (N3)? mem[465] : 
//                          (N0)? mem[1005] : 1'b0;
//   assign r_data_o[464] = (N3)? mem[464] : 
//                          (N0)? mem[1004] : 1'b0;
//   assign r_data_o[463] = (N3)? mem[463] : 
//                          (N0)? mem[1003] : 1'b0;
//   assign r_data_o[462] = (N3)? mem[462] : 
//                          (N0)? mem[1002] : 1'b0;
//   assign r_data_o[461] = (N3)? mem[461] : 
//                          (N0)? mem[1001] : 1'b0;
//   assign r_data_o[460] = (N3)? mem[460] : 
//                          (N0)? mem[1000] : 1'b0;
//   assign r_data_o[459] = (N3)? mem[459] : 
//                          (N0)? mem[999] : 1'b0;
//   assign r_data_o[458] = (N3)? mem[458] : 
//                          (N0)? mem[998] : 1'b0;
//   assign r_data_o[457] = (N3)? mem[457] : 
//                          (N0)? mem[997] : 1'b0;
//   assign r_data_o[456] = (N3)? mem[456] : 
//                          (N0)? mem[996] : 1'b0;
//   assign r_data_o[455] = (N3)? mem[455] : 
//                          (N0)? mem[995] : 1'b0;
//   assign r_data_o[454] = (N3)? mem[454] : 
//                          (N0)? mem[994] : 1'b0;
//   assign r_data_o[453] = (N3)? mem[453] : 
//                          (N0)? mem[993] : 1'b0;
//   assign r_data_o[452] = (N3)? mem[452] : 
//                          (N0)? mem[992] : 1'b0;
//   assign r_data_o[451] = (N3)? mem[451] : 
//                          (N0)? mem[991] : 1'b0;
//   assign r_data_o[450] = (N3)? mem[450] : 
//                          (N0)? mem[990] : 1'b0;
//   assign r_data_o[449] = (N3)? mem[449] : 
//                          (N0)? mem[989] : 1'b0;
//   assign r_data_o[448] = (N3)? mem[448] : 
//                          (N0)? mem[988] : 1'b0;
//   assign r_data_o[447] = (N3)? mem[447] : 
//                          (N0)? mem[987] : 1'b0;
//   assign r_data_o[446] = (N3)? mem[446] : 
//                          (N0)? mem[986] : 1'b0;
//   assign r_data_o[445] = (N3)? mem[445] : 
//                          (N0)? mem[985] : 1'b0;
//   assign r_data_o[444] = (N3)? mem[444] : 
//                          (N0)? mem[984] : 1'b0;
//   assign r_data_o[443] = (N3)? mem[443] : 
//                          (N0)? mem[983] : 1'b0;
//   assign r_data_o[442] = (N3)? mem[442] : 
//                          (N0)? mem[982] : 1'b0;
//   assign r_data_o[441] = (N3)? mem[441] : 
//                          (N0)? mem[981] : 1'b0;
//   assign r_data_o[440] = (N3)? mem[440] : 
//                          (N0)? mem[980] : 1'b0;
//   assign r_data_o[439] = (N3)? mem[439] : 
//                          (N0)? mem[979] : 1'b0;
//   assign r_data_o[438] = (N3)? mem[438] : 
//                          (N0)? mem[978] : 1'b0;
//   assign r_data_o[437] = (N3)? mem[437] : 
//                          (N0)? mem[977] : 1'b0;
//   assign r_data_o[436] = (N3)? mem[436] : 
//                          (N0)? mem[976] : 1'b0;
//   assign r_data_o[435] = (N3)? mem[435] : 
//                          (N0)? mem[975] : 1'b0;
//   assign r_data_o[434] = (N3)? mem[434] : 
//                          (N0)? mem[974] : 1'b0;
//   assign r_data_o[433] = (N3)? mem[433] : 
//                          (N0)? mem[973] : 1'b0;
//   assign r_data_o[432] = (N3)? mem[432] : 
//                          (N0)? mem[972] : 1'b0;
//   assign r_data_o[431] = (N3)? mem[431] : 
//                          (N0)? mem[971] : 1'b0;
//   assign r_data_o[430] = (N3)? mem[430] : 
//                          (N0)? mem[970] : 1'b0;
//   assign r_data_o[429] = (N3)? mem[429] : 
//                          (N0)? mem[969] : 1'b0;
//   assign r_data_o[428] = (N3)? mem[428] : 
//                          (N0)? mem[968] : 1'b0;
//   assign r_data_o[427] = (N3)? mem[427] : 
//                          (N0)? mem[967] : 1'b0;
//   assign r_data_o[426] = (N3)? mem[426] : 
//                          (N0)? mem[966] : 1'b0;
//   assign r_data_o[425] = (N3)? mem[425] : 
//                          (N0)? mem[965] : 1'b0;
//   assign r_data_o[424] = (N3)? mem[424] : 
//                          (N0)? mem[964] : 1'b0;
//   assign r_data_o[423] = (N3)? mem[423] : 
//                          (N0)? mem[963] : 1'b0;
//   assign r_data_o[422] = (N3)? mem[422] : 
//                          (N0)? mem[962] : 1'b0;
//   assign r_data_o[421] = (N3)? mem[421] : 
//                          (N0)? mem[961] : 1'b0;
//   assign r_data_o[420] = (N3)? mem[420] : 
//                          (N0)? mem[960] : 1'b0;
//   assign r_data_o[419] = (N3)? mem[419] : 
//                          (N0)? mem[959] : 1'b0;
//   assign r_data_o[418] = (N3)? mem[418] : 
//                          (N0)? mem[958] : 1'b0;
//   assign r_data_o[417] = (N3)? mem[417] : 
//                          (N0)? mem[957] : 1'b0;
//   assign r_data_o[416] = (N3)? mem[416] : 
//                          (N0)? mem[956] : 1'b0;
//   assign r_data_o[415] = (N3)? mem[415] : 
//                          (N0)? mem[955] : 1'b0;
//   assign r_data_o[414] = (N3)? mem[414] : 
//                          (N0)? mem[954] : 1'b0;
//   assign r_data_o[413] = (N3)? mem[413] : 
//                          (N0)? mem[953] : 1'b0;
//   assign r_data_o[412] = (N3)? mem[412] : 
//                          (N0)? mem[952] : 1'b0;
//   assign r_data_o[411] = (N3)? mem[411] : 
//                          (N0)? mem[951] : 1'b0;
//   assign r_data_o[410] = (N3)? mem[410] : 
//                          (N0)? mem[950] : 1'b0;
//   assign r_data_o[409] = (N3)? mem[409] : 
//                          (N0)? mem[949] : 1'b0;
//   assign r_data_o[408] = (N3)? mem[408] : 
//                          (N0)? mem[948] : 1'b0;
//   assign r_data_o[407] = (N3)? mem[407] : 
//                          (N0)? mem[947] : 1'b0;
//   assign r_data_o[406] = (N3)? mem[406] : 
//                          (N0)? mem[946] : 1'b0;
//   assign r_data_o[405] = (N3)? mem[405] : 
//                          (N0)? mem[945] : 1'b0;
//   assign r_data_o[404] = (N3)? mem[404] : 
//                          (N0)? mem[944] : 1'b0;
//   assign r_data_o[403] = (N3)? mem[403] : 
//                          (N0)? mem[943] : 1'b0;
//   assign r_data_o[402] = (N3)? mem[402] : 
//                          (N0)? mem[942] : 1'b0;
//   assign r_data_o[401] = (N3)? mem[401] : 
//                          (N0)? mem[941] : 1'b0;
//   assign r_data_o[400] = (N3)? mem[400] : 
//                          (N0)? mem[940] : 1'b0;
//   assign r_data_o[399] = (N3)? mem[399] : 
//                          (N0)? mem[939] : 1'b0;
//   assign r_data_o[398] = (N3)? mem[398] : 
//                          (N0)? mem[938] : 1'b0;
//   assign r_data_o[397] = (N3)? mem[397] : 
//                          (N0)? mem[937] : 1'b0;
//   assign r_data_o[396] = (N3)? mem[396] : 
//                          (N0)? mem[936] : 1'b0;
//   assign r_data_o[395] = (N3)? mem[395] : 
//                          (N0)? mem[935] : 1'b0;
//   assign r_data_o[394] = (N3)? mem[394] : 
//                          (N0)? mem[934] : 1'b0;
//   assign r_data_o[393] = (N3)? mem[393] : 
//                          (N0)? mem[933] : 1'b0;
//   assign r_data_o[392] = (N3)? mem[392] : 
//                          (N0)? mem[932] : 1'b0;
//   assign r_data_o[391] = (N3)? mem[391] : 
//                          (N0)? mem[931] : 1'b0;
//   assign r_data_o[390] = (N3)? mem[390] : 
//                          (N0)? mem[930] : 1'b0;
//   assign r_data_o[389] = (N3)? mem[389] : 
//                          (N0)? mem[929] : 1'b0;
//   assign r_data_o[388] = (N3)? mem[388] : 
//                          (N0)? mem[928] : 1'b0;
//   assign r_data_o[387] = (N3)? mem[387] : 
//                          (N0)? mem[927] : 1'b0;
//   assign r_data_o[386] = (N3)? mem[386] : 
//                          (N0)? mem[926] : 1'b0;
//   assign r_data_o[385] = (N3)? mem[385] : 
//                          (N0)? mem[925] : 1'b0;
//   assign r_data_o[384] = (N3)? mem[384] : 
//                          (N0)? mem[924] : 1'b0;
//   assign r_data_o[383] = (N3)? mem[383] : 
//                          (N0)? mem[923] : 1'b0;
//   assign r_data_o[382] = (N3)? mem[382] : 
//                          (N0)? mem[922] : 1'b0;
//   assign r_data_o[381] = (N3)? mem[381] : 
//                          (N0)? mem[921] : 1'b0;
//   assign r_data_o[380] = (N3)? mem[380] : 
//                          (N0)? mem[920] : 1'b0;
//   assign r_data_o[379] = (N3)? mem[379] : 
//                          (N0)? mem[919] : 1'b0;
//   assign r_data_o[378] = (N3)? mem[378] : 
//                          (N0)? mem[918] : 1'b0;
//   assign r_data_o[377] = (N3)? mem[377] : 
//                          (N0)? mem[917] : 1'b0;
//   assign r_data_o[376] = (N3)? mem[376] : 
//                          (N0)? mem[916] : 1'b0;
//   assign r_data_o[375] = (N3)? mem[375] : 
//                          (N0)? mem[915] : 1'b0;
//   assign r_data_o[374] = (N3)? mem[374] : 
//                          (N0)? mem[914] : 1'b0;
//   assign r_data_o[373] = (N3)? mem[373] : 
//                          (N0)? mem[913] : 1'b0;
//   assign r_data_o[372] = (N3)? mem[372] : 
//                          (N0)? mem[912] : 1'b0;
//   assign r_data_o[371] = (N3)? mem[371] : 
//                          (N0)? mem[911] : 1'b0;
//   assign r_data_o[370] = (N3)? mem[370] : 
//                          (N0)? mem[910] : 1'b0;
//   assign r_data_o[369] = (N3)? mem[369] : 
//                          (N0)? mem[909] : 1'b0;
//   assign r_data_o[368] = (N3)? mem[368] : 
//                          (N0)? mem[908] : 1'b0;
//   assign r_data_o[367] = (N3)? mem[367] : 
//                          (N0)? mem[907] : 1'b0;
//   assign r_data_o[366] = (N3)? mem[366] : 
//                          (N0)? mem[906] : 1'b0;
//   assign r_data_o[365] = (N3)? mem[365] : 
//                          (N0)? mem[905] : 1'b0;
//   assign r_data_o[364] = (N3)? mem[364] : 
//                          (N0)? mem[904] : 1'b0;
//   assign r_data_o[363] = (N3)? mem[363] : 
//                          (N0)? mem[903] : 1'b0;
//   assign r_data_o[362] = (N3)? mem[362] : 
//                          (N0)? mem[902] : 1'b0;
//   assign r_data_o[361] = (N3)? mem[361] : 
//                          (N0)? mem[901] : 1'b0;
//   assign r_data_o[360] = (N3)? mem[360] : 
//                          (N0)? mem[900] : 1'b0;
//   assign r_data_o[359] = (N3)? mem[359] : 
//                          (N0)? mem[899] : 1'b0;
//   assign r_data_o[358] = (N3)? mem[358] : 
//                          (N0)? mem[898] : 1'b0;
//   assign r_data_o[357] = (N3)? mem[357] : 
//                          (N0)? mem[897] : 1'b0;
//   assign r_data_o[356] = (N3)? mem[356] : 
//                          (N0)? mem[896] : 1'b0;
//   assign r_data_o[355] = (N3)? mem[355] : 
//                          (N0)? mem[895] : 1'b0;
//   assign r_data_o[354] = (N3)? mem[354] : 
//                          (N0)? mem[894] : 1'b0;
//   assign r_data_o[353] = (N3)? mem[353] : 
//                          (N0)? mem[893] : 1'b0;
//   assign r_data_o[352] = (N3)? mem[352] : 
//                          (N0)? mem[892] : 1'b0;
//   assign r_data_o[351] = (N3)? mem[351] : 
//                          (N0)? mem[891] : 1'b0;
//   assign r_data_o[350] = (N3)? mem[350] : 
//                          (N0)? mem[890] : 1'b0;
//   assign r_data_o[349] = (N3)? mem[349] : 
//                          (N0)? mem[889] : 1'b0;
//   assign r_data_o[348] = (N3)? mem[348] : 
//                          (N0)? mem[888] : 1'b0;
//   assign r_data_o[347] = (N3)? mem[347] : 
//                          (N0)? mem[887] : 1'b0;
//   assign r_data_o[346] = (N3)? mem[346] : 
//                          (N0)? mem[886] : 1'b0;
//   assign r_data_o[345] = (N3)? mem[345] : 
//                          (N0)? mem[885] : 1'b0;
//   assign r_data_o[344] = (N3)? mem[344] : 
//                          (N0)? mem[884] : 1'b0;
//   assign r_data_o[343] = (N3)? mem[343] : 
//                          (N0)? mem[883] : 1'b0;
//   assign r_data_o[342] = (N3)? mem[342] : 
//                          (N0)? mem[882] : 1'b0;
//   assign r_data_o[341] = (N3)? mem[341] : 
//                          (N0)? mem[881] : 1'b0;
//   assign r_data_o[340] = (N3)? mem[340] : 
//                          (N0)? mem[880] : 1'b0;
//   assign r_data_o[339] = (N3)? mem[339] : 
//                          (N0)? mem[879] : 1'b0;
//   assign r_data_o[338] = (N3)? mem[338] : 
//                          (N0)? mem[878] : 1'b0;
//   assign r_data_o[337] = (N3)? mem[337] : 
//                          (N0)? mem[877] : 1'b0;
//   assign r_data_o[336] = (N3)? mem[336] : 
//                          (N0)? mem[876] : 1'b0;
//   assign r_data_o[335] = (N3)? mem[335] : 
//                          (N0)? mem[875] : 1'b0;
//   assign r_data_o[334] = (N3)? mem[334] : 
//                          (N0)? mem[874] : 1'b0;
//   assign r_data_o[333] = (N3)? mem[333] : 
//                          (N0)? mem[873] : 1'b0;
//   assign r_data_o[332] = (N3)? mem[332] : 
//                          (N0)? mem[872] : 1'b0;
//   assign r_data_o[331] = (N3)? mem[331] : 
//                          (N0)? mem[871] : 1'b0;
//   assign r_data_o[330] = (N3)? mem[330] : 
//                          (N0)? mem[870] : 1'b0;
//   assign r_data_o[329] = (N3)? mem[329] : 
//                          (N0)? mem[869] : 1'b0;
//   assign r_data_o[328] = (N3)? mem[328] : 
//                          (N0)? mem[868] : 1'b0;
//   assign r_data_o[327] = (N3)? mem[327] : 
//                          (N0)? mem[867] : 1'b0;
//   assign r_data_o[326] = (N3)? mem[326] : 
//                          (N0)? mem[866] : 1'b0;
//   assign r_data_o[325] = (N3)? mem[325] : 
//                          (N0)? mem[865] : 1'b0;
//   assign r_data_o[324] = (N3)? mem[324] : 
//                          (N0)? mem[864] : 1'b0;
//   assign r_data_o[323] = (N3)? mem[323] : 
//                          (N0)? mem[863] : 1'b0;
//   assign r_data_o[322] = (N3)? mem[322] : 
//                          (N0)? mem[862] : 1'b0;
//   assign r_data_o[321] = (N3)? mem[321] : 
//                          (N0)? mem[861] : 1'b0;
//   assign r_data_o[320] = (N3)? mem[320] : 
//                          (N0)? mem[860] : 1'b0;
//   assign r_data_o[319] = (N3)? mem[319] : 
//                          (N0)? mem[859] : 1'b0;
//   assign r_data_o[318] = (N3)? mem[318] : 
//                          (N0)? mem[858] : 1'b0;
//   assign r_data_o[317] = (N3)? mem[317] : 
//                          (N0)? mem[857] : 1'b0;
//   assign r_data_o[316] = (N3)? mem[316] : 
//                          (N0)? mem[856] : 1'b0;
//   assign r_data_o[315] = (N3)? mem[315] : 
//                          (N0)? mem[855] : 1'b0;
//   assign r_data_o[314] = (N3)? mem[314] : 
//                          (N0)? mem[854] : 1'b0;
//   assign r_data_o[313] = (N3)? mem[313] : 
//                          (N0)? mem[853] : 1'b0;
//   assign r_data_o[312] = (N3)? mem[312] : 
//                          (N0)? mem[852] : 1'b0;
//   assign r_data_o[311] = (N3)? mem[311] : 
//                          (N0)? mem[851] : 1'b0;
//   assign r_data_o[310] = (N3)? mem[310] : 
//                          (N0)? mem[850] : 1'b0;
//   assign r_data_o[309] = (N3)? mem[309] : 
//                          (N0)? mem[849] : 1'b0;
//   assign r_data_o[308] = (N3)? mem[308] : 
//                          (N0)? mem[848] : 1'b0;
//   assign r_data_o[307] = (N3)? mem[307] : 
//                          (N0)? mem[847] : 1'b0;
//   assign r_data_o[306] = (N3)? mem[306] : 
//                          (N0)? mem[846] : 1'b0;
//   assign r_data_o[305] = (N3)? mem[305] : 
//                          (N0)? mem[845] : 1'b0;
//   assign r_data_o[304] = (N3)? mem[304] : 
//                          (N0)? mem[844] : 1'b0;
//   assign r_data_o[303] = (N3)? mem[303] : 
//                          (N0)? mem[843] : 1'b0;
//   assign r_data_o[302] = (N3)? mem[302] : 
//                          (N0)? mem[842] : 1'b0;
//   assign r_data_o[301] = (N3)? mem[301] : 
//                          (N0)? mem[841] : 1'b0;
//   assign r_data_o[300] = (N3)? mem[300] : 
//                          (N0)? mem[840] : 1'b0;
//   assign r_data_o[299] = (N3)? mem[299] : 
//                          (N0)? mem[839] : 1'b0;
//   assign r_data_o[298] = (N3)? mem[298] : 
//                          (N0)? mem[838] : 1'b0;
//   assign r_data_o[297] = (N3)? mem[297] : 
//                          (N0)? mem[837] : 1'b0;
//   assign r_data_o[296] = (N3)? mem[296] : 
//                          (N0)? mem[836] : 1'b0;
//   assign r_data_o[295] = (N3)? mem[295] : 
//                          (N0)? mem[835] : 1'b0;
//   assign r_data_o[294] = (N3)? mem[294] : 
//                          (N0)? mem[834] : 1'b0;
//   assign r_data_o[293] = (N3)? mem[293] : 
//                          (N0)? mem[833] : 1'b0;
//   assign r_data_o[292] = (N3)? mem[292] : 
//                          (N0)? mem[832] : 1'b0;
//   assign r_data_o[291] = (N3)? mem[291] : 
//                          (N0)? mem[831] : 1'b0;
//   assign r_data_o[290] = (N3)? mem[290] : 
//                          (N0)? mem[830] : 1'b0;
//   assign r_data_o[289] = (N3)? mem[289] : 
//                          (N0)? mem[829] : 1'b0;
//   assign r_data_o[288] = (N3)? mem[288] : 
//                          (N0)? mem[828] : 1'b0;
//   assign r_data_o[287] = (N3)? mem[287] : 
//                          (N0)? mem[827] : 1'b0;
//   assign r_data_o[286] = (N3)? mem[286] : 
//                          (N0)? mem[826] : 1'b0;
//   assign r_data_o[285] = (N3)? mem[285] : 
//                          (N0)? mem[825] : 1'b0;
//   assign r_data_o[284] = (N3)? mem[284] : 
//                          (N0)? mem[824] : 1'b0;
//   assign r_data_o[283] = (N3)? mem[283] : 
//                          (N0)? mem[823] : 1'b0;
//   assign r_data_o[282] = (N3)? mem[282] : 
//                          (N0)? mem[822] : 1'b0;
//   assign r_data_o[281] = (N3)? mem[281] : 
//                          (N0)? mem[821] : 1'b0;
//   assign r_data_o[280] = (N3)? mem[280] : 
//                          (N0)? mem[820] : 1'b0;
//   assign r_data_o[279] = (N3)? mem[279] : 
//                          (N0)? mem[819] : 1'b0;
//   assign r_data_o[278] = (N3)? mem[278] : 
//                          (N0)? mem[818] : 1'b0;
//   assign r_data_o[277] = (N3)? mem[277] : 
//                          (N0)? mem[817] : 1'b0;
//   assign r_data_o[276] = (N3)? mem[276] : 
//                          (N0)? mem[816] : 1'b0;
//   assign r_data_o[275] = (N3)? mem[275] : 
//                          (N0)? mem[815] : 1'b0;
//   assign r_data_o[274] = (N3)? mem[274] : 
//                          (N0)? mem[814] : 1'b0;
//   assign r_data_o[273] = (N3)? mem[273] : 
//                          (N0)? mem[813] : 1'b0;
//   assign r_data_o[272] = (N3)? mem[272] : 
//                          (N0)? mem[812] : 1'b0;
//   assign r_data_o[271] = (N3)? mem[271] : 
//                          (N0)? mem[811] : 1'b0;
//   assign r_data_o[270] = (N3)? mem[270] : 
//                          (N0)? mem[810] : 1'b0;
//   assign r_data_o[269] = (N3)? mem[269] : 
//                          (N0)? mem[809] : 1'b0;
//   assign r_data_o[268] = (N3)? mem[268] : 
//                          (N0)? mem[808] : 1'b0;
//   assign r_data_o[267] = (N3)? mem[267] : 
//                          (N0)? mem[807] : 1'b0;
//   assign r_data_o[266] = (N3)? mem[266] : 
//                          (N0)? mem[806] : 1'b0;
//   assign r_data_o[265] = (N3)? mem[265] : 
//                          (N0)? mem[805] : 1'b0;
//   assign r_data_o[264] = (N3)? mem[264] : 
//                          (N0)? mem[804] : 1'b0;
//   assign r_data_o[263] = (N3)? mem[263] : 
//                          (N0)? mem[803] : 1'b0;
//   assign r_data_o[262] = (N3)? mem[262] : 
//                          (N0)? mem[802] : 1'b0;
//   assign r_data_o[261] = (N3)? mem[261] : 
//                          (N0)? mem[801] : 1'b0;
//   assign r_data_o[260] = (N3)? mem[260] : 
//                          (N0)? mem[800] : 1'b0;
//   assign r_data_o[259] = (N3)? mem[259] : 
//                          (N0)? mem[799] : 1'b0;
//   assign r_data_o[258] = (N3)? mem[258] : 
//                          (N0)? mem[798] : 1'b0;
//   assign r_data_o[257] = (N3)? mem[257] : 
//                          (N0)? mem[797] : 1'b0;
//   assign r_data_o[256] = (N3)? mem[256] : 
//                          (N0)? mem[796] : 1'b0;
//   assign r_data_o[255] = (N3)? mem[255] : 
//                          (N0)? mem[795] : 1'b0;
//   assign r_data_o[254] = (N3)? mem[254] : 
//                          (N0)? mem[794] : 1'b0;
//   assign r_data_o[253] = (N3)? mem[253] : 
//                          (N0)? mem[793] : 1'b0;
//   assign r_data_o[252] = (N3)? mem[252] : 
//                          (N0)? mem[792] : 1'b0;
//   assign r_data_o[251] = (N3)? mem[251] : 
//                          (N0)? mem[791] : 1'b0;
//   assign r_data_o[250] = (N3)? mem[250] : 
//                          (N0)? mem[790] : 1'b0;
//   assign r_data_o[249] = (N3)? mem[249] : 
//                          (N0)? mem[789] : 1'b0;
//   assign r_data_o[248] = (N3)? mem[248] : 
//                          (N0)? mem[788] : 1'b0;
//   assign r_data_o[247] = (N3)? mem[247] : 
//                          (N0)? mem[787] : 1'b0;
//   assign r_data_o[246] = (N3)? mem[246] : 
//                          (N0)? mem[786] : 1'b0;
//   assign r_data_o[245] = (N3)? mem[245] : 
//                          (N0)? mem[785] : 1'b0;
//   assign r_data_o[244] = (N3)? mem[244] : 
//                          (N0)? mem[784] : 1'b0;
//   assign r_data_o[243] = (N3)? mem[243] : 
//                          (N0)? mem[783] : 1'b0;
//   assign r_data_o[242] = (N3)? mem[242] : 
//                          (N0)? mem[782] : 1'b0;
//   assign r_data_o[241] = (N3)? mem[241] : 
//                          (N0)? mem[781] : 1'b0;
//   assign r_data_o[240] = (N3)? mem[240] : 
//                          (N0)? mem[780] : 1'b0;
//   assign r_data_o[239] = (N3)? mem[239] : 
//                          (N0)? mem[779] : 1'b0;
//   assign r_data_o[238] = (N3)? mem[238] : 
//                          (N0)? mem[778] : 1'b0;
//   assign r_data_o[237] = (N3)? mem[237] : 
//                          (N0)? mem[777] : 1'b0;
//   assign r_data_o[236] = (N3)? mem[236] : 
//                          (N0)? mem[776] : 1'b0;
//   assign r_data_o[235] = (N3)? mem[235] : 
//                          (N0)? mem[775] : 1'b0;
//   assign r_data_o[234] = (N3)? mem[234] : 
//                          (N0)? mem[774] : 1'b0;
//   assign r_data_o[233] = (N3)? mem[233] : 
//                          (N0)? mem[773] : 1'b0;
//   assign r_data_o[232] = (N3)? mem[232] : 
//                          (N0)? mem[772] : 1'b0;
//   assign r_data_o[231] = (N3)? mem[231] : 
//                          (N0)? mem[771] : 1'b0;
//   assign r_data_o[230] = (N3)? mem[230] : 
//                          (N0)? mem[770] : 1'b0;
//   assign r_data_o[229] = (N3)? mem[229] : 
//                          (N0)? mem[769] : 1'b0;
//   assign r_data_o[228] = (N3)? mem[228] : 
//                          (N0)? mem[768] : 1'b0;
//   assign r_data_o[227] = (N3)? mem[227] : 
//                          (N0)? mem[767] : 1'b0;
//   assign r_data_o[226] = (N3)? mem[226] : 
//                          (N0)? mem[766] : 1'b0;
//   assign r_data_o[225] = (N3)? mem[225] : 
//                          (N0)? mem[765] : 1'b0;
//   assign r_data_o[224] = (N3)? mem[224] : 
//                          (N0)? mem[764] : 1'b0;
//   assign r_data_o[223] = (N3)? mem[223] : 
//                          (N0)? mem[763] : 1'b0;
//   assign r_data_o[222] = (N3)? mem[222] : 
//                          (N0)? mem[762] : 1'b0;
//   assign r_data_o[221] = (N3)? mem[221] : 
//                          (N0)? mem[761] : 1'b0;
//   assign r_data_o[220] = (N3)? mem[220] : 
//                          (N0)? mem[760] : 1'b0;
//   assign r_data_o[219] = (N3)? mem[219] : 
//                          (N0)? mem[759] : 1'b0;
//   assign r_data_o[218] = (N3)? mem[218] : 
//                          (N0)? mem[758] : 1'b0;
//   assign r_data_o[217] = (N3)? mem[217] : 
//                          (N0)? mem[757] : 1'b0;
//   assign r_data_o[216] = (N3)? mem[216] : 
//                          (N0)? mem[756] : 1'b0;
//   assign r_data_o[215] = (N3)? mem[215] : 
//                          (N0)? mem[755] : 1'b0;
//   assign r_data_o[214] = (N3)? mem[214] : 
//                          (N0)? mem[754] : 1'b0;
//   assign r_data_o[213] = (N3)? mem[213] : 
//                          (N0)? mem[753] : 1'b0;
//   assign r_data_o[212] = (N3)? mem[212] : 
//                          (N0)? mem[752] : 1'b0;
//   assign r_data_o[211] = (N3)? mem[211] : 
//                          (N0)? mem[751] : 1'b0;
//   assign r_data_o[210] = (N3)? mem[210] : 
//                          (N0)? mem[750] : 1'b0;
//   assign r_data_o[209] = (N3)? mem[209] : 
//                          (N0)? mem[749] : 1'b0;
//   assign r_data_o[208] = (N3)? mem[208] : 
//                          (N0)? mem[748] : 1'b0;
//   assign r_data_o[207] = (N3)? mem[207] : 
//                          (N0)? mem[747] : 1'b0;
//   assign r_data_o[206] = (N3)? mem[206] : 
//                          (N0)? mem[746] : 1'b0;
//   assign r_data_o[205] = (N3)? mem[205] : 
//                          (N0)? mem[745] : 1'b0;
//   assign r_data_o[204] = (N3)? mem[204] : 
//                          (N0)? mem[744] : 1'b0;
//   assign r_data_o[203] = (N3)? mem[203] : 
//                          (N0)? mem[743] : 1'b0;
//   assign r_data_o[202] = (N3)? mem[202] : 
//                          (N0)? mem[742] : 1'b0;
//   assign r_data_o[201] = (N3)? mem[201] : 
//                          (N0)? mem[741] : 1'b0;
//   assign r_data_o[200] = (N3)? mem[200] : 
//                          (N0)? mem[740] : 1'b0;
//   assign r_data_o[199] = (N3)? mem[199] : 
//                          (N0)? mem[739] : 1'b0;
//   assign r_data_o[198] = (N3)? mem[198] : 
//                          (N0)? mem[738] : 1'b0;
//   assign r_data_o[197] = (N3)? mem[197] : 
//                          (N0)? mem[737] : 1'b0;
//   assign r_data_o[196] = (N3)? mem[196] : 
//                          (N0)? mem[736] : 1'b0;
//   assign r_data_o[195] = (N3)? mem[195] : 
//                          (N0)? mem[735] : 1'b0;
//   assign r_data_o[194] = (N3)? mem[194] : 
//                          (N0)? mem[734] : 1'b0;
//   assign r_data_o[193] = (N3)? mem[193] : 
//                          (N0)? mem[733] : 1'b0;
//   assign r_data_o[192] = (N3)? mem[192] : 
//                          (N0)? mem[732] : 1'b0;
//   assign r_data_o[191] = (N3)? mem[191] : 
//                          (N0)? mem[731] : 1'b0;
//   assign r_data_o[190] = (N3)? mem[190] : 
//                          (N0)? mem[730] : 1'b0;
//   assign r_data_o[189] = (N3)? mem[189] : 
//                          (N0)? mem[729] : 1'b0;
//   assign r_data_o[188] = (N3)? mem[188] : 
//                          (N0)? mem[728] : 1'b0;
//   assign r_data_o[187] = (N3)? mem[187] : 
//                          (N0)? mem[727] : 1'b0;
//   assign r_data_o[186] = (N3)? mem[186] : 
//                          (N0)? mem[726] : 1'b0;
//   assign r_data_o[185] = (N3)? mem[185] : 
//                          (N0)? mem[725] : 1'b0;
//   assign r_data_o[184] = (N3)? mem[184] : 
//                          (N0)? mem[724] : 1'b0;
//   assign r_data_o[183] = (N3)? mem[183] : 
//                          (N0)? mem[723] : 1'b0;
//   assign r_data_o[182] = (N3)? mem[182] : 
//                          (N0)? mem[722] : 1'b0;
//   assign r_data_o[181] = (N3)? mem[181] : 
//                          (N0)? mem[721] : 1'b0;
//   assign r_data_o[180] = (N3)? mem[180] : 
//                          (N0)? mem[720] : 1'b0;
//   assign r_data_o[179] = (N3)? mem[179] : 
//                          (N0)? mem[719] : 1'b0;
//   assign r_data_o[178] = (N3)? mem[178] : 
//                          (N0)? mem[718] : 1'b0;
//   assign r_data_o[177] = (N3)? mem[177] : 
//                          (N0)? mem[717] : 1'b0;
//   assign r_data_o[176] = (N3)? mem[176] : 
//                          (N0)? mem[716] : 1'b0;
//   assign r_data_o[175] = (N3)? mem[175] : 
//                          (N0)? mem[715] : 1'b0;
//   assign r_data_o[174] = (N3)? mem[174] : 
//                          (N0)? mem[714] : 1'b0;
//   assign r_data_o[173] = (N3)? mem[173] : 
//                          (N0)? mem[713] : 1'b0;
//   assign r_data_o[172] = (N3)? mem[172] : 
//                          (N0)? mem[712] : 1'b0;
//   assign r_data_o[171] = (N3)? mem[171] : 
//                          (N0)? mem[711] : 1'b0;
//   assign r_data_o[170] = (N3)? mem[170] : 
//                          (N0)? mem[710] : 1'b0;
//   assign r_data_o[169] = (N3)? mem[169] : 
//                          (N0)? mem[709] : 1'b0;
//   assign r_data_o[168] = (N3)? mem[168] : 
//                          (N0)? mem[708] : 1'b0;
//   assign r_data_o[167] = (N3)? mem[167] : 
//                          (N0)? mem[707] : 1'b0;
//   assign r_data_o[166] = (N3)? mem[166] : 
//                          (N0)? mem[706] : 1'b0;
//   assign r_data_o[165] = (N3)? mem[165] : 
//                          (N0)? mem[705] : 1'b0;
//   assign r_data_o[164] = (N3)? mem[164] : 
//                          (N0)? mem[704] : 1'b0;
//   assign r_data_o[163] = (N3)? mem[163] : 
//                          (N0)? mem[703] : 1'b0;
//   assign r_data_o[162] = (N3)? mem[162] : 
//                          (N0)? mem[702] : 1'b0;
//   assign r_data_o[161] = (N3)? mem[161] : 
//                          (N0)? mem[701] : 1'b0;
//   assign r_data_o[160] = (N3)? mem[160] : 
//                          (N0)? mem[700] : 1'b0;
//   assign r_data_o[159] = (N3)? mem[159] : 
//                          (N0)? mem[699] : 1'b0;
//   assign r_data_o[158] = (N3)? mem[158] : 
//                          (N0)? mem[698] : 1'b0;
//   assign r_data_o[157] = (N3)? mem[157] : 
//                          (N0)? mem[697] : 1'b0;
//   assign r_data_o[156] = (N3)? mem[156] : 
//                          (N0)? mem[696] : 1'b0;
//   assign r_data_o[155] = (N3)? mem[155] : 
//                          (N0)? mem[695] : 1'b0;
//   assign r_data_o[154] = (N3)? mem[154] : 
//                          (N0)? mem[694] : 1'b0;
//   assign r_data_o[153] = (N3)? mem[153] : 
//                          (N0)? mem[693] : 1'b0;
//   assign r_data_o[152] = (N3)? mem[152] : 
//                          (N0)? mem[692] : 1'b0;
//   assign r_data_o[151] = (N3)? mem[151] : 
//                          (N0)? mem[691] : 1'b0;
//   assign r_data_o[150] = (N3)? mem[150] : 
//                          (N0)? mem[690] : 1'b0;
//   assign r_data_o[149] = (N3)? mem[149] : 
//                          (N0)? mem[689] : 1'b0;
//   assign r_data_o[148] = (N3)? mem[148] : 
//                          (N0)? mem[688] : 1'b0;
//   assign r_data_o[147] = (N3)? mem[147] : 
//                          (N0)? mem[687] : 1'b0;
//   assign r_data_o[146] = (N3)? mem[146] : 
//                          (N0)? mem[686] : 1'b0;
//   assign r_data_o[145] = (N3)? mem[145] : 
//                          (N0)? mem[685] : 1'b0;
//   assign r_data_o[144] = (N3)? mem[144] : 
//                          (N0)? mem[684] : 1'b0;
//   assign r_data_o[143] = (N3)? mem[143] : 
//                          (N0)? mem[683] : 1'b0;
//   assign r_data_o[142] = (N3)? mem[142] : 
//                          (N0)? mem[682] : 1'b0;
//   assign r_data_o[141] = (N3)? mem[141] : 
//                          (N0)? mem[681] : 1'b0;
//   assign r_data_o[140] = (N3)? mem[140] : 
//                          (N0)? mem[680] : 1'b0;
//   assign r_data_o[139] = (N3)? mem[139] : 
//                          (N0)? mem[679] : 1'b0;
//   assign r_data_o[138] = (N3)? mem[138] : 
//                          (N0)? mem[678] : 1'b0;
//   assign r_data_o[137] = (N3)? mem[137] : 
//                          (N0)? mem[677] : 1'b0;
//   assign r_data_o[136] = (N3)? mem[136] : 
//                          (N0)? mem[676] : 1'b0;
//   assign r_data_o[135] = (N3)? mem[135] : 
//                          (N0)? mem[675] : 1'b0;
//   assign r_data_o[134] = (N3)? mem[134] : 
//                          (N0)? mem[674] : 1'b0;
//   assign r_data_o[133] = (N3)? mem[133] : 
//                          (N0)? mem[673] : 1'b0;
//   assign r_data_o[132] = (N3)? mem[132] : 
//                          (N0)? mem[672] : 1'b0;
//   assign r_data_o[131] = (N3)? mem[131] : 
//                          (N0)? mem[671] : 1'b0;
//   assign r_data_o[130] = (N3)? mem[130] : 
//                          (N0)? mem[670] : 1'b0;
//   assign r_data_o[129] = (N3)? mem[129] : 
//                          (N0)? mem[669] : 1'b0;
//   assign r_data_o[128] = (N3)? mem[128] : 
//                          (N0)? mem[668] : 1'b0;
//   assign r_data_o[127] = (N3)? mem[127] : 
//                          (N0)? mem[667] : 1'b0;
//   assign r_data_o[126] = (N3)? mem[126] : 
//                          (N0)? mem[666] : 1'b0;
//   assign r_data_o[125] = (N3)? mem[125] : 
//                          (N0)? mem[665] : 1'b0;
//   assign r_data_o[124] = (N3)? mem[124] : 
//                          (N0)? mem[664] : 1'b0;
//   assign r_data_o[123] = (N3)? mem[123] : 
//                          (N0)? mem[663] : 1'b0;
//   assign r_data_o[122] = (N3)? mem[122] : 
//                          (N0)? mem[662] : 1'b0;
//   assign r_data_o[121] = (N3)? mem[121] : 
//                          (N0)? mem[661] : 1'b0;
//   assign r_data_o[120] = (N3)? mem[120] : 
//                          (N0)? mem[660] : 1'b0;
//   assign r_data_o[119] = (N3)? mem[119] : 
//                          (N0)? mem[659] : 1'b0;
//   assign r_data_o[118] = (N3)? mem[118] : 
//                          (N0)? mem[658] : 1'b0;
//   assign r_data_o[117] = (N3)? mem[117] : 
//                          (N0)? mem[657] : 1'b0;
//   assign r_data_o[116] = (N3)? mem[116] : 
//                          (N0)? mem[656] : 1'b0;
//   assign r_data_o[115] = (N3)? mem[115] : 
//                          (N0)? mem[655] : 1'b0;
//   assign r_data_o[114] = (N3)? mem[114] : 
//                          (N0)? mem[654] : 1'b0;
//   assign r_data_o[113] = (N3)? mem[113] : 
//                          (N0)? mem[653] : 1'b0;
//   assign r_data_o[112] = (N3)? mem[112] : 
//                          (N0)? mem[652] : 1'b0;
//   assign r_data_o[111] = (N3)? mem[111] : 
//                          (N0)? mem[651] : 1'b0;
//   assign r_data_o[110] = (N3)? mem[110] : 
//                          (N0)? mem[650] : 1'b0;
//   assign r_data_o[109] = (N3)? mem[109] : 
//                          (N0)? mem[649] : 1'b0;
//   assign r_data_o[108] = (N3)? mem[108] : 
//                          (N0)? mem[648] : 1'b0;
//   assign r_data_o[107] = (N3)? mem[107] : 
//                          (N0)? mem[647] : 1'b0;
//   assign r_data_o[106] = (N3)? mem[106] : 
//                          (N0)? mem[646] : 1'b0;
//   assign r_data_o[105] = (N3)? mem[105] : 
//                          (N0)? mem[645] : 1'b0;
//   assign r_data_o[104] = (N3)? mem[104] : 
//                          (N0)? mem[644] : 1'b0;
//   assign r_data_o[103] = (N3)? mem[103] : 
//                          (N0)? mem[643] : 1'b0;
//   assign r_data_o[102] = (N3)? mem[102] : 
//                          (N0)? mem[642] : 1'b0;
//   assign r_data_o[101] = (N3)? mem[101] : 
//                          (N0)? mem[641] : 1'b0;
//   assign r_data_o[100] = (N3)? mem[100] : 
//                          (N0)? mem[640] : 1'b0;
//   assign r_data_o[99] = (N3)? mem[99] : 
//                         (N0)? mem[639] : 1'b0;
//   assign r_data_o[98] = (N3)? mem[98] : 
//                         (N0)? mem[638] : 1'b0;
//   assign r_data_o[97] = (N3)? mem[97] : 
//                         (N0)? mem[637] : 1'b0;
//   assign r_data_o[96] = (N3)? mem[96] : 
//                         (N0)? mem[636] : 1'b0;
//   assign r_data_o[95] = (N3)? mem[95] : 
//                         (N0)? mem[635] : 1'b0;
//   assign r_data_o[94] = (N3)? mem[94] : 
//                         (N0)? mem[634] : 1'b0;
//   assign r_data_o[93] = (N3)? mem[93] : 
//                         (N0)? mem[633] : 1'b0;
//   assign r_data_o[92] = (N3)? mem[92] : 
//                         (N0)? mem[632] : 1'b0;
//   assign r_data_o[91] = (N3)? mem[91] : 
//                         (N0)? mem[631] : 1'b0;
//   assign r_data_o[90] = (N3)? mem[90] : 
//                         (N0)? mem[630] : 1'b0;
//   assign r_data_o[89] = (N3)? mem[89] : 
//                         (N0)? mem[629] : 1'b0;
//   assign r_data_o[88] = (N3)? mem[88] : 
//                         (N0)? mem[628] : 1'b0;
//   assign r_data_o[87] = (N3)? mem[87] : 
//                         (N0)? mem[627] : 1'b0;
//   assign r_data_o[86] = (N3)? mem[86] : 
//                         (N0)? mem[626] : 1'b0;
//   assign r_data_o[85] = (N3)? mem[85] : 
//                         (N0)? mem[625] : 1'b0;
//   assign r_data_o[84] = (N3)? mem[84] : 
//                         (N0)? mem[624] : 1'b0;
//   assign r_data_o[83] = (N3)? mem[83] : 
//                         (N0)? mem[623] : 1'b0;
//   assign r_data_o[82] = (N3)? mem[82] : 
//                         (N0)? mem[622] : 1'b0;
//   assign r_data_o[81] = (N3)? mem[81] : 
//                         (N0)? mem[621] : 1'b0;
//   assign r_data_o[80] = (N3)? mem[80] : 
//                         (N0)? mem[620] : 1'b0;
//   assign r_data_o[79] = (N3)? mem[79] : 
//                         (N0)? mem[619] : 1'b0;
//   assign r_data_o[78] = (N3)? mem[78] : 
//                         (N0)? mem[618] : 1'b0;
//   assign r_data_o[77] = (N3)? mem[77] : 
//                         (N0)? mem[617] : 1'b0;
//   assign r_data_o[76] = (N3)? mem[76] : 
//                         (N0)? mem[616] : 1'b0;
//   assign r_data_o[75] = (N3)? mem[75] : 
//                         (N0)? mem[615] : 1'b0;
//   assign r_data_o[74] = (N3)? mem[74] : 
//                         (N0)? mem[614] : 1'b0;
//   assign r_data_o[73] = (N3)? mem[73] : 
//                         (N0)? mem[613] : 1'b0;
//   assign r_data_o[72] = (N3)? mem[72] : 
//                         (N0)? mem[612] : 1'b0;
//   assign r_data_o[71] = (N3)? mem[71] : 
//                         (N0)? mem[611] : 1'b0;
//   assign r_data_o[70] = (N3)? mem[70] : 
//                         (N0)? mem[610] : 1'b0;
//   assign r_data_o[69] = (N3)? mem[69] : 
//                         (N0)? mem[609] : 1'b0;
//   assign r_data_o[68] = (N3)? mem[68] : 
//                         (N0)? mem[608] : 1'b0;
//   assign r_data_o[67] = (N3)? mem[67] : 
//                         (N0)? mem[607] : 1'b0;
//   assign r_data_o[66] = (N3)? mem[66] : 
//                         (N0)? mem[606] : 1'b0;
//   assign r_data_o[65] = (N3)? mem[65] : 
//                         (N0)? mem[605] : 1'b0;
//   assign r_data_o[64] = (N3)? mem[64] : 
//                         (N0)? mem[604] : 1'b0;
//   assign r_data_o[63] = (N3)? mem[63] : 
//                         (N0)? mem[603] : 1'b0;
//   assign r_data_o[62] = (N3)? mem[62] : 
//                         (N0)? mem[602] : 1'b0;
//   assign r_data_o[61] = (N3)? mem[61] : 
//                         (N0)? mem[601] : 1'b0;
//   assign r_data_o[60] = (N3)? mem[60] : 
//                         (N0)? mem[600] : 1'b0;
//   assign r_data_o[59] = (N3)? mem[59] : 
//                         (N0)? mem[599] : 1'b0;
//   assign r_data_o[58] = (N3)? mem[58] : 
//                         (N0)? mem[598] : 1'b0;
//   assign r_data_o[57] = (N3)? mem[57] : 
//                         (N0)? mem[597] : 1'b0;
//   assign r_data_o[56] = (N3)? mem[56] : 
//                         (N0)? mem[596] : 1'b0;
//   assign r_data_o[55] = (N3)? mem[55] : 
//                         (N0)? mem[595] : 1'b0;
//   assign r_data_o[54] = (N3)? mem[54] : 
//                         (N0)? mem[594] : 1'b0;
//   assign r_data_o[53] = (N3)? mem[53] : 
//                         (N0)? mem[593] : 1'b0;
//   assign r_data_o[52] = (N3)? mem[52] : 
//                         (N0)? mem[592] : 1'b0;
//   assign r_data_o[51] = (N3)? mem[51] : 
//                         (N0)? mem[591] : 1'b0;
//   assign r_data_o[50] = (N3)? mem[50] : 
//                         (N0)? mem[590] : 1'b0;
//   assign r_data_o[49] = (N3)? mem[49] : 
//                         (N0)? mem[589] : 1'b0;
//   assign r_data_o[48] = (N3)? mem[48] : 
//                         (N0)? mem[588] : 1'b0;
//   assign r_data_o[47] = (N3)? mem[47] : 
//                         (N0)? mem[587] : 1'b0;
//   assign r_data_o[46] = (N3)? mem[46] : 
//                         (N0)? mem[586] : 1'b0;
//   assign r_data_o[45] = (N3)? mem[45] : 
//                         (N0)? mem[585] : 1'b0;
//   assign r_data_o[44] = (N3)? mem[44] : 
//                         (N0)? mem[584] : 1'b0;
//   assign r_data_o[43] = (N3)? mem[43] : 
//                         (N0)? mem[583] : 1'b0;
//   assign r_data_o[42] = (N3)? mem[42] : 
//                         (N0)? mem[582] : 1'b0;
//   assign r_data_o[41] = (N3)? mem[41] : 
//                         (N0)? mem[581] : 1'b0;
//   assign r_data_o[40] = (N3)? mem[40] : 
//                         (N0)? mem[580] : 1'b0;
//   assign r_data_o[39] = (N3)? mem[39] : 
//                         (N0)? mem[579] : 1'b0;
//   assign r_data_o[38] = (N3)? mem[38] : 
//                         (N0)? mem[578] : 1'b0;
//   assign r_data_o[37] = (N3)? mem[37] : 
//                         (N0)? mem[577] : 1'b0;
//   assign r_data_o[36] = (N3)? mem[36] : 
//                         (N0)? mem[576] : 1'b0;
//   assign r_data_o[35] = (N3)? mem[35] : 
//                         (N0)? mem[575] : 1'b0;
//   assign r_data_o[34] = (N3)? mem[34] : 
//                         (N0)? mem[574] : 1'b0;
//   assign r_data_o[33] = (N3)? mem[33] : 
//                         (N0)? mem[573] : 1'b0;
//   assign r_data_o[32] = (N3)? mem[32] : 
//                         (N0)? mem[572] : 1'b0;
//   assign r_data_o[31] = (N3)? mem[31] : 
//                         (N0)? mem[571] : 1'b0;
//   assign r_data_o[30] = (N3)? mem[30] : 
//                         (N0)? mem[570] : 1'b0;
//   assign r_data_o[29] = (N3)? mem[29] : 
//                         (N0)? mem[569] : 1'b0;
//   assign r_data_o[28] = (N3)? mem[28] : 
//                         (N0)? mem[568] : 1'b0;
//   assign r_data_o[27] = (N3)? mem[27] : 
//                         (N0)? mem[567] : 1'b0;
//   assign r_data_o[26] = (N3)? mem[26] : 
//                         (N0)? mem[566] : 1'b0;
//   assign r_data_o[25] = (N3)? mem[25] : 
//                         (N0)? mem[565] : 1'b0;
//   assign r_data_o[24] = (N3)? mem[24] : 
//                         (N0)? mem[564] : 1'b0;
//   assign r_data_o[23] = (N3)? mem[23] : 
//                         (N0)? mem[563] : 1'b0;
//   assign r_data_o[22] = (N3)? mem[22] : 
//                         (N0)? mem[562] : 1'b0;
//   assign r_data_o[21] = (N3)? mem[21] : 
//                         (N0)? mem[561] : 1'b0;
//   assign r_data_o[20] = (N3)? mem[20] : 
//                         (N0)? mem[560] : 1'b0;
//   assign r_data_o[19] = (N3)? mem[19] : 
//                         (N0)? mem[559] : 1'b0;
//   assign r_data_o[18] = (N3)? mem[18] : 
//                         (N0)? mem[558] : 1'b0;
//   assign r_data_o[17] = (N3)? mem[17] : 
//                         (N0)? mem[557] : 1'b0;
//   assign r_data_o[16] = (N3)? mem[16] : 
//                         (N0)? mem[556] : 1'b0;
//   assign r_data_o[15] = (N3)? mem[15] : 
//                         (N0)? mem[555] : 1'b0;
//   assign r_data_o[14] = (N3)? mem[14] : 
//                         (N0)? mem[554] : 1'b0;
//   assign r_data_o[13] = (N3)? mem[13] : 
//                         (N0)? mem[553] : 1'b0;
//   assign r_data_o[12] = (N3)? mem[12] : 
//                         (N0)? mem[552] : 1'b0;
//   assign r_data_o[11] = (N3)? mem[11] : 
//                         (N0)? mem[551] : 1'b0;
//   assign r_data_o[10] = (N3)? mem[10] : 
//                         (N0)? mem[550] : 1'b0;
//   assign r_data_o[9] = (N3)? mem[9] : 
//                        (N0)? mem[549] : 1'b0;
//   assign r_data_o[8] = (N3)? mem[8] : 
//                        (N0)? mem[548] : 1'b0;
//   assign r_data_o[7] = (N3)? mem[7] : 
//                        (N0)? mem[547] : 1'b0;
//   assign r_data_o[6] = (N3)? mem[6] : 
//                        (N0)? mem[546] : 1'b0;
//   assign r_data_o[5] = (N3)? mem[5] : 
//                        (N0)? mem[545] : 1'b0;
//   assign r_data_o[4] = (N3)? mem[4] : 
//                        (N0)? mem[544] : 1'b0;
//   assign r_data_o[3] = (N3)? mem[3] : 
//                        (N0)? mem[543] : 1'b0;
//   assign r_data_o[2] = (N3)? mem[2] : 
//                        (N0)? mem[542] : 1'b0;
//   assign r_data_o[1] = (N3)? mem[1] : 
//                        (N0)? mem[541] : 1'b0;
//   assign r_data_o[0] = (N3)? mem[0] : 
//                        (N0)? mem[540] : 1'b0;
//   assign N5 = ~w_addr_i[0];
//   assign { N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], N5, N5, N5, N5, N5, N5 } : 
//                                                                        (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
//   assign N1 = w_v_i;
//   assign N2 = N4;
//   assign N3 = ~r_addr_i[0];
//   assign N4 = ~w_v_i;

//   always @(posedge w_clk_i) begin
//     if(N13) begin
//       { mem[1079:981], mem[540:540] } <= { w_data_i[539:441], w_data_i[0:0] };
//     end 
//     if(N14) begin
//       { mem[980:882], mem[541:541] } <= { w_data_i[440:342], w_data_i[1:1] };
//     end 
//     if(N15) begin
//       { mem[881:783], mem[542:542] } <= { w_data_i[341:243], w_data_i[2:2] };
//     end 
//     if(N16) begin
//       { mem[782:684], mem[543:543] } <= { w_data_i[242:144], w_data_i[3:3] };
//     end 
//     if(N17) begin
//       { mem[683:585], mem[544:544] } <= { w_data_i[143:45], w_data_i[4:4] };
//     end 
//     if(N18) begin
//       { mem[584:545] } <= { w_data_i[44:5] };
//     end 
//     if(N7) begin
//       { mem[539:441], mem[0:0] } <= { w_data_i[539:441], w_data_i[0:0] };
//     end 
//     if(N8) begin
//       { mem[440:342], mem[1:1] } <= { w_data_i[440:342], w_data_i[1:1] };
//     end 
//     if(N9) begin
//       { mem[341:243], mem[2:2] } <= { w_data_i[341:243], w_data_i[2:2] };
//     end 
//     if(N10) begin
//       { mem[242:144], mem[3:3] } <= { w_data_i[242:144], w_data_i[3:3] };
//     end 
//     if(N11) begin
//       { mem[143:45], mem[4:4] } <= { w_data_i[143:45], w_data_i[4:4] };
//     end 
//     if(N12) begin
//       { mem[44:5] } <= { w_data_i[44:5] };
//     end 
//   end


// endmodule



module bsg_mem_1r1w_width_p540_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [539:0] w_data_i;
  input [0:0] r_addr_i;
  output [539:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [539:0] r_data_o;

  bsg_mem_p540
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p540
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [539:0] data_i;
  output [539:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [539:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p540_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 : 
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 : 
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 : 
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 : 
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 : 
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 : 
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end 
    if(N9) begin
      tail_r <= N10;
    end 
    if(N11) begin
      head_r <= N12;
    end 
  end


endmodule



module bp_fe_lce_data_cmd_data_width_p64_lce_addr_width_p22_lce_data_width_p512_num_cce_p1_num_lce_p2_lce_sets_p64_ways_p8_block_size_in_bytes_p8
(
  cce_data_received_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_yumi_o,
  data_mem_pkt_v_o,
  data_mem_pkt_o,
  data_mem_pkt_yumi_i
);

  input [539:0] lce_data_cmd_i;
  output [521:0] data_mem_pkt_o;
  input lce_data_cmd_v_i;
  input data_mem_pkt_yumi_i;
  output cce_data_received_o;
  output lce_data_cmd_yumi_o;
  output data_mem_pkt_v_o;
  wire [521:0] data_mem_pkt_o;
  wire cce_data_received_o,lce_data_cmd_yumi_o,data_mem_pkt_v_o,data_mem_pkt_yumi_i,
  lce_data_cmd_v_i;
  assign data_mem_pkt_o[512] = 1'b1;
  assign lce_data_cmd_yumi_o = data_mem_pkt_yumi_i;
  assign data_mem_pkt_v_o = lce_data_cmd_v_i;
  assign data_mem_pkt_o[521] = lce_data_cmd_i[523];
  assign data_mem_pkt_o[520] = lce_data_cmd_i[522];
  assign data_mem_pkt_o[519] = lce_data_cmd_i[521];
  assign data_mem_pkt_o[518] = lce_data_cmd_i[520];
  assign data_mem_pkt_o[517] = lce_data_cmd_i[519];
  assign data_mem_pkt_o[516] = lce_data_cmd_i[518];
  assign data_mem_pkt_o[515] = lce_data_cmd_i[536];
  assign data_mem_pkt_o[514] = lce_data_cmd_i[535];
  assign data_mem_pkt_o[513] = lce_data_cmd_i[534];
  assign data_mem_pkt_o[511] = lce_data_cmd_i[511];
  assign data_mem_pkt_o[510] = lce_data_cmd_i[510];
  assign data_mem_pkt_o[509] = lce_data_cmd_i[509];
  assign data_mem_pkt_o[508] = lce_data_cmd_i[508];
  assign data_mem_pkt_o[507] = lce_data_cmd_i[507];
  assign data_mem_pkt_o[506] = lce_data_cmd_i[506];
  assign data_mem_pkt_o[505] = lce_data_cmd_i[505];
  assign data_mem_pkt_o[504] = lce_data_cmd_i[504];
  assign data_mem_pkt_o[503] = lce_data_cmd_i[503];
  assign data_mem_pkt_o[502] = lce_data_cmd_i[502];
  assign data_mem_pkt_o[501] = lce_data_cmd_i[501];
  assign data_mem_pkt_o[500] = lce_data_cmd_i[500];
  assign data_mem_pkt_o[499] = lce_data_cmd_i[499];
  assign data_mem_pkt_o[498] = lce_data_cmd_i[498];
  assign data_mem_pkt_o[497] = lce_data_cmd_i[497];
  assign data_mem_pkt_o[496] = lce_data_cmd_i[496];
  assign data_mem_pkt_o[495] = lce_data_cmd_i[495];
  assign data_mem_pkt_o[494] = lce_data_cmd_i[494];
  assign data_mem_pkt_o[493] = lce_data_cmd_i[493];
  assign data_mem_pkt_o[492] = lce_data_cmd_i[492];
  assign data_mem_pkt_o[491] = lce_data_cmd_i[491];
  assign data_mem_pkt_o[490] = lce_data_cmd_i[490];
  assign data_mem_pkt_o[489] = lce_data_cmd_i[489];
  assign data_mem_pkt_o[488] = lce_data_cmd_i[488];
  assign data_mem_pkt_o[487] = lce_data_cmd_i[487];
  assign data_mem_pkt_o[486] = lce_data_cmd_i[486];
  assign data_mem_pkt_o[485] = lce_data_cmd_i[485];
  assign data_mem_pkt_o[484] = lce_data_cmd_i[484];
  assign data_mem_pkt_o[483] = lce_data_cmd_i[483];
  assign data_mem_pkt_o[482] = lce_data_cmd_i[482];
  assign data_mem_pkt_o[481] = lce_data_cmd_i[481];
  assign data_mem_pkt_o[480] = lce_data_cmd_i[480];
  assign data_mem_pkt_o[479] = lce_data_cmd_i[479];
  assign data_mem_pkt_o[478] = lce_data_cmd_i[478];
  assign data_mem_pkt_o[477] = lce_data_cmd_i[477];
  assign data_mem_pkt_o[476] = lce_data_cmd_i[476];
  assign data_mem_pkt_o[475] = lce_data_cmd_i[475];
  assign data_mem_pkt_o[474] = lce_data_cmd_i[474];
  assign data_mem_pkt_o[473] = lce_data_cmd_i[473];
  assign data_mem_pkt_o[472] = lce_data_cmd_i[472];
  assign data_mem_pkt_o[471] = lce_data_cmd_i[471];
  assign data_mem_pkt_o[470] = lce_data_cmd_i[470];
  assign data_mem_pkt_o[469] = lce_data_cmd_i[469];
  assign data_mem_pkt_o[468] = lce_data_cmd_i[468];
  assign data_mem_pkt_o[467] = lce_data_cmd_i[467];
  assign data_mem_pkt_o[466] = lce_data_cmd_i[466];
  assign data_mem_pkt_o[465] = lce_data_cmd_i[465];
  assign data_mem_pkt_o[464] = lce_data_cmd_i[464];
  assign data_mem_pkt_o[463] = lce_data_cmd_i[463];
  assign data_mem_pkt_o[462] = lce_data_cmd_i[462];
  assign data_mem_pkt_o[461] = lce_data_cmd_i[461];
  assign data_mem_pkt_o[460] = lce_data_cmd_i[460];
  assign data_mem_pkt_o[459] = lce_data_cmd_i[459];
  assign data_mem_pkt_o[458] = lce_data_cmd_i[458];
  assign data_mem_pkt_o[457] = lce_data_cmd_i[457];
  assign data_mem_pkt_o[456] = lce_data_cmd_i[456];
  assign data_mem_pkt_o[455] = lce_data_cmd_i[455];
  assign data_mem_pkt_o[454] = lce_data_cmd_i[454];
  assign data_mem_pkt_o[453] = lce_data_cmd_i[453];
  assign data_mem_pkt_o[452] = lce_data_cmd_i[452];
  assign data_mem_pkt_o[451] = lce_data_cmd_i[451];
  assign data_mem_pkt_o[450] = lce_data_cmd_i[450];
  assign data_mem_pkt_o[449] = lce_data_cmd_i[449];
  assign data_mem_pkt_o[448] = lce_data_cmd_i[448];
  assign data_mem_pkt_o[447] = lce_data_cmd_i[447];
  assign data_mem_pkt_o[446] = lce_data_cmd_i[446];
  assign data_mem_pkt_o[445] = lce_data_cmd_i[445];
  assign data_mem_pkt_o[444] = lce_data_cmd_i[444];
  assign data_mem_pkt_o[443] = lce_data_cmd_i[443];
  assign data_mem_pkt_o[442] = lce_data_cmd_i[442];
  assign data_mem_pkt_o[441] = lce_data_cmd_i[441];
  assign data_mem_pkt_o[440] = lce_data_cmd_i[440];
  assign data_mem_pkt_o[439] = lce_data_cmd_i[439];
  assign data_mem_pkt_o[438] = lce_data_cmd_i[438];
  assign data_mem_pkt_o[437] = lce_data_cmd_i[437];
  assign data_mem_pkt_o[436] = lce_data_cmd_i[436];
  assign data_mem_pkt_o[435] = lce_data_cmd_i[435];
  assign data_mem_pkt_o[434] = lce_data_cmd_i[434];
  assign data_mem_pkt_o[433] = lce_data_cmd_i[433];
  assign data_mem_pkt_o[432] = lce_data_cmd_i[432];
  assign data_mem_pkt_o[431] = lce_data_cmd_i[431];
  assign data_mem_pkt_o[430] = lce_data_cmd_i[430];
  assign data_mem_pkt_o[429] = lce_data_cmd_i[429];
  assign data_mem_pkt_o[428] = lce_data_cmd_i[428];
  assign data_mem_pkt_o[427] = lce_data_cmd_i[427];
  assign data_mem_pkt_o[426] = lce_data_cmd_i[426];
  assign data_mem_pkt_o[425] = lce_data_cmd_i[425];
  assign data_mem_pkt_o[424] = lce_data_cmd_i[424];
  assign data_mem_pkt_o[423] = lce_data_cmd_i[423];
  assign data_mem_pkt_o[422] = lce_data_cmd_i[422];
  assign data_mem_pkt_o[421] = lce_data_cmd_i[421];
  assign data_mem_pkt_o[420] = lce_data_cmd_i[420];
  assign data_mem_pkt_o[419] = lce_data_cmd_i[419];
  assign data_mem_pkt_o[418] = lce_data_cmd_i[418];
  assign data_mem_pkt_o[417] = lce_data_cmd_i[417];
  assign data_mem_pkt_o[416] = lce_data_cmd_i[416];
  assign data_mem_pkt_o[415] = lce_data_cmd_i[415];
  assign data_mem_pkt_o[414] = lce_data_cmd_i[414];
  assign data_mem_pkt_o[413] = lce_data_cmd_i[413];
  assign data_mem_pkt_o[412] = lce_data_cmd_i[412];
  assign data_mem_pkt_o[411] = lce_data_cmd_i[411];
  assign data_mem_pkt_o[410] = lce_data_cmd_i[410];
  assign data_mem_pkt_o[409] = lce_data_cmd_i[409];
  assign data_mem_pkt_o[408] = lce_data_cmd_i[408];
  assign data_mem_pkt_o[407] = lce_data_cmd_i[407];
  assign data_mem_pkt_o[406] = lce_data_cmd_i[406];
  assign data_mem_pkt_o[405] = lce_data_cmd_i[405];
  assign data_mem_pkt_o[404] = lce_data_cmd_i[404];
  assign data_mem_pkt_o[403] = lce_data_cmd_i[403];
  assign data_mem_pkt_o[402] = lce_data_cmd_i[402];
  assign data_mem_pkt_o[401] = lce_data_cmd_i[401];
  assign data_mem_pkt_o[400] = lce_data_cmd_i[400];
  assign data_mem_pkt_o[399] = lce_data_cmd_i[399];
  assign data_mem_pkt_o[398] = lce_data_cmd_i[398];
  assign data_mem_pkt_o[397] = lce_data_cmd_i[397];
  assign data_mem_pkt_o[396] = lce_data_cmd_i[396];
  assign data_mem_pkt_o[395] = lce_data_cmd_i[395];
  assign data_mem_pkt_o[394] = lce_data_cmd_i[394];
  assign data_mem_pkt_o[393] = lce_data_cmd_i[393];
  assign data_mem_pkt_o[392] = lce_data_cmd_i[392];
  assign data_mem_pkt_o[391] = lce_data_cmd_i[391];
  assign data_mem_pkt_o[390] = lce_data_cmd_i[390];
  assign data_mem_pkt_o[389] = lce_data_cmd_i[389];
  assign data_mem_pkt_o[388] = lce_data_cmd_i[388];
  assign data_mem_pkt_o[387] = lce_data_cmd_i[387];
  assign data_mem_pkt_o[386] = lce_data_cmd_i[386];
  assign data_mem_pkt_o[385] = lce_data_cmd_i[385];
  assign data_mem_pkt_o[384] = lce_data_cmd_i[384];
  assign data_mem_pkt_o[383] = lce_data_cmd_i[383];
  assign data_mem_pkt_o[382] = lce_data_cmd_i[382];
  assign data_mem_pkt_o[381] = lce_data_cmd_i[381];
  assign data_mem_pkt_o[380] = lce_data_cmd_i[380];
  assign data_mem_pkt_o[379] = lce_data_cmd_i[379];
  assign data_mem_pkt_o[378] = lce_data_cmd_i[378];
  assign data_mem_pkt_o[377] = lce_data_cmd_i[377];
  assign data_mem_pkt_o[376] = lce_data_cmd_i[376];
  assign data_mem_pkt_o[375] = lce_data_cmd_i[375];
  assign data_mem_pkt_o[374] = lce_data_cmd_i[374];
  assign data_mem_pkt_o[373] = lce_data_cmd_i[373];
  assign data_mem_pkt_o[372] = lce_data_cmd_i[372];
  assign data_mem_pkt_o[371] = lce_data_cmd_i[371];
  assign data_mem_pkt_o[370] = lce_data_cmd_i[370];
  assign data_mem_pkt_o[369] = lce_data_cmd_i[369];
  assign data_mem_pkt_o[368] = lce_data_cmd_i[368];
  assign data_mem_pkt_o[367] = lce_data_cmd_i[367];
  assign data_mem_pkt_o[366] = lce_data_cmd_i[366];
  assign data_mem_pkt_o[365] = lce_data_cmd_i[365];
  assign data_mem_pkt_o[364] = lce_data_cmd_i[364];
  assign data_mem_pkt_o[363] = lce_data_cmd_i[363];
  assign data_mem_pkt_o[362] = lce_data_cmd_i[362];
  assign data_mem_pkt_o[361] = lce_data_cmd_i[361];
  assign data_mem_pkt_o[360] = lce_data_cmd_i[360];
  assign data_mem_pkt_o[359] = lce_data_cmd_i[359];
  assign data_mem_pkt_o[358] = lce_data_cmd_i[358];
  assign data_mem_pkt_o[357] = lce_data_cmd_i[357];
  assign data_mem_pkt_o[356] = lce_data_cmd_i[356];
  assign data_mem_pkt_o[355] = lce_data_cmd_i[355];
  assign data_mem_pkt_o[354] = lce_data_cmd_i[354];
  assign data_mem_pkt_o[353] = lce_data_cmd_i[353];
  assign data_mem_pkt_o[352] = lce_data_cmd_i[352];
  assign data_mem_pkt_o[351] = lce_data_cmd_i[351];
  assign data_mem_pkt_o[350] = lce_data_cmd_i[350];
  assign data_mem_pkt_o[349] = lce_data_cmd_i[349];
  assign data_mem_pkt_o[348] = lce_data_cmd_i[348];
  assign data_mem_pkt_o[347] = lce_data_cmd_i[347];
  assign data_mem_pkt_o[346] = lce_data_cmd_i[346];
  assign data_mem_pkt_o[345] = lce_data_cmd_i[345];
  assign data_mem_pkt_o[344] = lce_data_cmd_i[344];
  assign data_mem_pkt_o[343] = lce_data_cmd_i[343];
  assign data_mem_pkt_o[342] = lce_data_cmd_i[342];
  assign data_mem_pkt_o[341] = lce_data_cmd_i[341];
  assign data_mem_pkt_o[340] = lce_data_cmd_i[340];
  assign data_mem_pkt_o[339] = lce_data_cmd_i[339];
  assign data_mem_pkt_o[338] = lce_data_cmd_i[338];
  assign data_mem_pkt_o[337] = lce_data_cmd_i[337];
  assign data_mem_pkt_o[336] = lce_data_cmd_i[336];
  assign data_mem_pkt_o[335] = lce_data_cmd_i[335];
  assign data_mem_pkt_o[334] = lce_data_cmd_i[334];
  assign data_mem_pkt_o[333] = lce_data_cmd_i[333];
  assign data_mem_pkt_o[332] = lce_data_cmd_i[332];
  assign data_mem_pkt_o[331] = lce_data_cmd_i[331];
  assign data_mem_pkt_o[330] = lce_data_cmd_i[330];
  assign data_mem_pkt_o[329] = lce_data_cmd_i[329];
  assign data_mem_pkt_o[328] = lce_data_cmd_i[328];
  assign data_mem_pkt_o[327] = lce_data_cmd_i[327];
  assign data_mem_pkt_o[326] = lce_data_cmd_i[326];
  assign data_mem_pkt_o[325] = lce_data_cmd_i[325];
  assign data_mem_pkt_o[324] = lce_data_cmd_i[324];
  assign data_mem_pkt_o[323] = lce_data_cmd_i[323];
  assign data_mem_pkt_o[322] = lce_data_cmd_i[322];
  assign data_mem_pkt_o[321] = lce_data_cmd_i[321];
  assign data_mem_pkt_o[320] = lce_data_cmd_i[320];
  assign data_mem_pkt_o[319] = lce_data_cmd_i[319];
  assign data_mem_pkt_o[318] = lce_data_cmd_i[318];
  assign data_mem_pkt_o[317] = lce_data_cmd_i[317];
  assign data_mem_pkt_o[316] = lce_data_cmd_i[316];
  assign data_mem_pkt_o[315] = lce_data_cmd_i[315];
  assign data_mem_pkt_o[314] = lce_data_cmd_i[314];
  assign data_mem_pkt_o[313] = lce_data_cmd_i[313];
  assign data_mem_pkt_o[312] = lce_data_cmd_i[312];
  assign data_mem_pkt_o[311] = lce_data_cmd_i[311];
  assign data_mem_pkt_o[310] = lce_data_cmd_i[310];
  assign data_mem_pkt_o[309] = lce_data_cmd_i[309];
  assign data_mem_pkt_o[308] = lce_data_cmd_i[308];
  assign data_mem_pkt_o[307] = lce_data_cmd_i[307];
  assign data_mem_pkt_o[306] = lce_data_cmd_i[306];
  assign data_mem_pkt_o[305] = lce_data_cmd_i[305];
  assign data_mem_pkt_o[304] = lce_data_cmd_i[304];
  assign data_mem_pkt_o[303] = lce_data_cmd_i[303];
  assign data_mem_pkt_o[302] = lce_data_cmd_i[302];
  assign data_mem_pkt_o[301] = lce_data_cmd_i[301];
  assign data_mem_pkt_o[300] = lce_data_cmd_i[300];
  assign data_mem_pkt_o[299] = lce_data_cmd_i[299];
  assign data_mem_pkt_o[298] = lce_data_cmd_i[298];
  assign data_mem_pkt_o[297] = lce_data_cmd_i[297];
  assign data_mem_pkt_o[296] = lce_data_cmd_i[296];
  assign data_mem_pkt_o[295] = lce_data_cmd_i[295];
  assign data_mem_pkt_o[294] = lce_data_cmd_i[294];
  assign data_mem_pkt_o[293] = lce_data_cmd_i[293];
  assign data_mem_pkt_o[292] = lce_data_cmd_i[292];
  assign data_mem_pkt_o[291] = lce_data_cmd_i[291];
  assign data_mem_pkt_o[290] = lce_data_cmd_i[290];
  assign data_mem_pkt_o[289] = lce_data_cmd_i[289];
  assign data_mem_pkt_o[288] = lce_data_cmd_i[288];
  assign data_mem_pkt_o[287] = lce_data_cmd_i[287];
  assign data_mem_pkt_o[286] = lce_data_cmd_i[286];
  assign data_mem_pkt_o[285] = lce_data_cmd_i[285];
  assign data_mem_pkt_o[284] = lce_data_cmd_i[284];
  assign data_mem_pkt_o[283] = lce_data_cmd_i[283];
  assign data_mem_pkt_o[282] = lce_data_cmd_i[282];
  assign data_mem_pkt_o[281] = lce_data_cmd_i[281];
  assign data_mem_pkt_o[280] = lce_data_cmd_i[280];
  assign data_mem_pkt_o[279] = lce_data_cmd_i[279];
  assign data_mem_pkt_o[278] = lce_data_cmd_i[278];
  assign data_mem_pkt_o[277] = lce_data_cmd_i[277];
  assign data_mem_pkt_o[276] = lce_data_cmd_i[276];
  assign data_mem_pkt_o[275] = lce_data_cmd_i[275];
  assign data_mem_pkt_o[274] = lce_data_cmd_i[274];
  assign data_mem_pkt_o[273] = lce_data_cmd_i[273];
  assign data_mem_pkt_o[272] = lce_data_cmd_i[272];
  assign data_mem_pkt_o[271] = lce_data_cmd_i[271];
  assign data_mem_pkt_o[270] = lce_data_cmd_i[270];
  assign data_mem_pkt_o[269] = lce_data_cmd_i[269];
  assign data_mem_pkt_o[268] = lce_data_cmd_i[268];
  assign data_mem_pkt_o[267] = lce_data_cmd_i[267];
  assign data_mem_pkt_o[266] = lce_data_cmd_i[266];
  assign data_mem_pkt_o[265] = lce_data_cmd_i[265];
  assign data_mem_pkt_o[264] = lce_data_cmd_i[264];
  assign data_mem_pkt_o[263] = lce_data_cmd_i[263];
  assign data_mem_pkt_o[262] = lce_data_cmd_i[262];
  assign data_mem_pkt_o[261] = lce_data_cmd_i[261];
  assign data_mem_pkt_o[260] = lce_data_cmd_i[260];
  assign data_mem_pkt_o[259] = lce_data_cmd_i[259];
  assign data_mem_pkt_o[258] = lce_data_cmd_i[258];
  assign data_mem_pkt_o[257] = lce_data_cmd_i[257];
  assign data_mem_pkt_o[256] = lce_data_cmd_i[256];
  assign data_mem_pkt_o[255] = lce_data_cmd_i[255];
  assign data_mem_pkt_o[254] = lce_data_cmd_i[254];
  assign data_mem_pkt_o[253] = lce_data_cmd_i[253];
  assign data_mem_pkt_o[252] = lce_data_cmd_i[252];
  assign data_mem_pkt_o[251] = lce_data_cmd_i[251];
  assign data_mem_pkt_o[250] = lce_data_cmd_i[250];
  assign data_mem_pkt_o[249] = lce_data_cmd_i[249];
  assign data_mem_pkt_o[248] = lce_data_cmd_i[248];
  assign data_mem_pkt_o[247] = lce_data_cmd_i[247];
  assign data_mem_pkt_o[246] = lce_data_cmd_i[246];
  assign data_mem_pkt_o[245] = lce_data_cmd_i[245];
  assign data_mem_pkt_o[244] = lce_data_cmd_i[244];
  assign data_mem_pkt_o[243] = lce_data_cmd_i[243];
  assign data_mem_pkt_o[242] = lce_data_cmd_i[242];
  assign data_mem_pkt_o[241] = lce_data_cmd_i[241];
  assign data_mem_pkt_o[240] = lce_data_cmd_i[240];
  assign data_mem_pkt_o[239] = lce_data_cmd_i[239];
  assign data_mem_pkt_o[238] = lce_data_cmd_i[238];
  assign data_mem_pkt_o[237] = lce_data_cmd_i[237];
  assign data_mem_pkt_o[236] = lce_data_cmd_i[236];
  assign data_mem_pkt_o[235] = lce_data_cmd_i[235];
  assign data_mem_pkt_o[234] = lce_data_cmd_i[234];
  assign data_mem_pkt_o[233] = lce_data_cmd_i[233];
  assign data_mem_pkt_o[232] = lce_data_cmd_i[232];
  assign data_mem_pkt_o[231] = lce_data_cmd_i[231];
  assign data_mem_pkt_o[230] = lce_data_cmd_i[230];
  assign data_mem_pkt_o[229] = lce_data_cmd_i[229];
  assign data_mem_pkt_o[228] = lce_data_cmd_i[228];
  assign data_mem_pkt_o[227] = lce_data_cmd_i[227];
  assign data_mem_pkt_o[226] = lce_data_cmd_i[226];
  assign data_mem_pkt_o[225] = lce_data_cmd_i[225];
  assign data_mem_pkt_o[224] = lce_data_cmd_i[224];
  assign data_mem_pkt_o[223] = lce_data_cmd_i[223];
  assign data_mem_pkt_o[222] = lce_data_cmd_i[222];
  assign data_mem_pkt_o[221] = lce_data_cmd_i[221];
  assign data_mem_pkt_o[220] = lce_data_cmd_i[220];
  assign data_mem_pkt_o[219] = lce_data_cmd_i[219];
  assign data_mem_pkt_o[218] = lce_data_cmd_i[218];
  assign data_mem_pkt_o[217] = lce_data_cmd_i[217];
  assign data_mem_pkt_o[216] = lce_data_cmd_i[216];
  assign data_mem_pkt_o[215] = lce_data_cmd_i[215];
  assign data_mem_pkt_o[214] = lce_data_cmd_i[214];
  assign data_mem_pkt_o[213] = lce_data_cmd_i[213];
  assign data_mem_pkt_o[212] = lce_data_cmd_i[212];
  assign data_mem_pkt_o[211] = lce_data_cmd_i[211];
  assign data_mem_pkt_o[210] = lce_data_cmd_i[210];
  assign data_mem_pkt_o[209] = lce_data_cmd_i[209];
  assign data_mem_pkt_o[208] = lce_data_cmd_i[208];
  assign data_mem_pkt_o[207] = lce_data_cmd_i[207];
  assign data_mem_pkt_o[206] = lce_data_cmd_i[206];
  assign data_mem_pkt_o[205] = lce_data_cmd_i[205];
  assign data_mem_pkt_o[204] = lce_data_cmd_i[204];
  assign data_mem_pkt_o[203] = lce_data_cmd_i[203];
  assign data_mem_pkt_o[202] = lce_data_cmd_i[202];
  assign data_mem_pkt_o[201] = lce_data_cmd_i[201];
  assign data_mem_pkt_o[200] = lce_data_cmd_i[200];
  assign data_mem_pkt_o[199] = lce_data_cmd_i[199];
  assign data_mem_pkt_o[198] = lce_data_cmd_i[198];
  assign data_mem_pkt_o[197] = lce_data_cmd_i[197];
  assign data_mem_pkt_o[196] = lce_data_cmd_i[196];
  assign data_mem_pkt_o[195] = lce_data_cmd_i[195];
  assign data_mem_pkt_o[194] = lce_data_cmd_i[194];
  assign data_mem_pkt_o[193] = lce_data_cmd_i[193];
  assign data_mem_pkt_o[192] = lce_data_cmd_i[192];
  assign data_mem_pkt_o[191] = lce_data_cmd_i[191];
  assign data_mem_pkt_o[190] = lce_data_cmd_i[190];
  assign data_mem_pkt_o[189] = lce_data_cmd_i[189];
  assign data_mem_pkt_o[188] = lce_data_cmd_i[188];
  assign data_mem_pkt_o[187] = lce_data_cmd_i[187];
  assign data_mem_pkt_o[186] = lce_data_cmd_i[186];
  assign data_mem_pkt_o[185] = lce_data_cmd_i[185];
  assign data_mem_pkt_o[184] = lce_data_cmd_i[184];
  assign data_mem_pkt_o[183] = lce_data_cmd_i[183];
  assign data_mem_pkt_o[182] = lce_data_cmd_i[182];
  assign data_mem_pkt_o[181] = lce_data_cmd_i[181];
  assign data_mem_pkt_o[180] = lce_data_cmd_i[180];
  assign data_mem_pkt_o[179] = lce_data_cmd_i[179];
  assign data_mem_pkt_o[178] = lce_data_cmd_i[178];
  assign data_mem_pkt_o[177] = lce_data_cmd_i[177];
  assign data_mem_pkt_o[176] = lce_data_cmd_i[176];
  assign data_mem_pkt_o[175] = lce_data_cmd_i[175];
  assign data_mem_pkt_o[174] = lce_data_cmd_i[174];
  assign data_mem_pkt_o[173] = lce_data_cmd_i[173];
  assign data_mem_pkt_o[172] = lce_data_cmd_i[172];
  assign data_mem_pkt_o[171] = lce_data_cmd_i[171];
  assign data_mem_pkt_o[170] = lce_data_cmd_i[170];
  assign data_mem_pkt_o[169] = lce_data_cmd_i[169];
  assign data_mem_pkt_o[168] = lce_data_cmd_i[168];
  assign data_mem_pkt_o[167] = lce_data_cmd_i[167];
  assign data_mem_pkt_o[166] = lce_data_cmd_i[166];
  assign data_mem_pkt_o[165] = lce_data_cmd_i[165];
  assign data_mem_pkt_o[164] = lce_data_cmd_i[164];
  assign data_mem_pkt_o[163] = lce_data_cmd_i[163];
  assign data_mem_pkt_o[162] = lce_data_cmd_i[162];
  assign data_mem_pkt_o[161] = lce_data_cmd_i[161];
  assign data_mem_pkt_o[160] = lce_data_cmd_i[160];
  assign data_mem_pkt_o[159] = lce_data_cmd_i[159];
  assign data_mem_pkt_o[158] = lce_data_cmd_i[158];
  assign data_mem_pkt_o[157] = lce_data_cmd_i[157];
  assign data_mem_pkt_o[156] = lce_data_cmd_i[156];
  assign data_mem_pkt_o[155] = lce_data_cmd_i[155];
  assign data_mem_pkt_o[154] = lce_data_cmd_i[154];
  assign data_mem_pkt_o[153] = lce_data_cmd_i[153];
  assign data_mem_pkt_o[152] = lce_data_cmd_i[152];
  assign data_mem_pkt_o[151] = lce_data_cmd_i[151];
  assign data_mem_pkt_o[150] = lce_data_cmd_i[150];
  assign data_mem_pkt_o[149] = lce_data_cmd_i[149];
  assign data_mem_pkt_o[148] = lce_data_cmd_i[148];
  assign data_mem_pkt_o[147] = lce_data_cmd_i[147];
  assign data_mem_pkt_o[146] = lce_data_cmd_i[146];
  assign data_mem_pkt_o[145] = lce_data_cmd_i[145];
  assign data_mem_pkt_o[144] = lce_data_cmd_i[144];
  assign data_mem_pkt_o[143] = lce_data_cmd_i[143];
  assign data_mem_pkt_o[142] = lce_data_cmd_i[142];
  assign data_mem_pkt_o[141] = lce_data_cmd_i[141];
  assign data_mem_pkt_o[140] = lce_data_cmd_i[140];
  assign data_mem_pkt_o[139] = lce_data_cmd_i[139];
  assign data_mem_pkt_o[138] = lce_data_cmd_i[138];
  assign data_mem_pkt_o[137] = lce_data_cmd_i[137];
  assign data_mem_pkt_o[136] = lce_data_cmd_i[136];
  assign data_mem_pkt_o[135] = lce_data_cmd_i[135];
  assign data_mem_pkt_o[134] = lce_data_cmd_i[134];
  assign data_mem_pkt_o[133] = lce_data_cmd_i[133];
  assign data_mem_pkt_o[132] = lce_data_cmd_i[132];
  assign data_mem_pkt_o[131] = lce_data_cmd_i[131];
  assign data_mem_pkt_o[130] = lce_data_cmd_i[130];
  assign data_mem_pkt_o[129] = lce_data_cmd_i[129];
  assign data_mem_pkt_o[128] = lce_data_cmd_i[128];
  assign data_mem_pkt_o[127] = lce_data_cmd_i[127];
  assign data_mem_pkt_o[126] = lce_data_cmd_i[126];
  assign data_mem_pkt_o[125] = lce_data_cmd_i[125];
  assign data_mem_pkt_o[124] = lce_data_cmd_i[124];
  assign data_mem_pkt_o[123] = lce_data_cmd_i[123];
  assign data_mem_pkt_o[122] = lce_data_cmd_i[122];
  assign data_mem_pkt_o[121] = lce_data_cmd_i[121];
  assign data_mem_pkt_o[120] = lce_data_cmd_i[120];
  assign data_mem_pkt_o[119] = lce_data_cmd_i[119];
  assign data_mem_pkt_o[118] = lce_data_cmd_i[118];
  assign data_mem_pkt_o[117] = lce_data_cmd_i[117];
  assign data_mem_pkt_o[116] = lce_data_cmd_i[116];
  assign data_mem_pkt_o[115] = lce_data_cmd_i[115];
  assign data_mem_pkt_o[114] = lce_data_cmd_i[114];
  assign data_mem_pkt_o[113] = lce_data_cmd_i[113];
  assign data_mem_pkt_o[112] = lce_data_cmd_i[112];
  assign data_mem_pkt_o[111] = lce_data_cmd_i[111];
  assign data_mem_pkt_o[110] = lce_data_cmd_i[110];
  assign data_mem_pkt_o[109] = lce_data_cmd_i[109];
  assign data_mem_pkt_o[108] = lce_data_cmd_i[108];
  assign data_mem_pkt_o[107] = lce_data_cmd_i[107];
  assign data_mem_pkt_o[106] = lce_data_cmd_i[106];
  assign data_mem_pkt_o[105] = lce_data_cmd_i[105];
  assign data_mem_pkt_o[104] = lce_data_cmd_i[104];
  assign data_mem_pkt_o[103] = lce_data_cmd_i[103];
  assign data_mem_pkt_o[102] = lce_data_cmd_i[102];
  assign data_mem_pkt_o[101] = lce_data_cmd_i[101];
  assign data_mem_pkt_o[100] = lce_data_cmd_i[100];
  assign data_mem_pkt_o[99] = lce_data_cmd_i[99];
  assign data_mem_pkt_o[98] = lce_data_cmd_i[98];
  assign data_mem_pkt_o[97] = lce_data_cmd_i[97];
  assign data_mem_pkt_o[96] = lce_data_cmd_i[96];
  assign data_mem_pkt_o[95] = lce_data_cmd_i[95];
  assign data_mem_pkt_o[94] = lce_data_cmd_i[94];
  assign data_mem_pkt_o[93] = lce_data_cmd_i[93];
  assign data_mem_pkt_o[92] = lce_data_cmd_i[92];
  assign data_mem_pkt_o[91] = lce_data_cmd_i[91];
  assign data_mem_pkt_o[90] = lce_data_cmd_i[90];
  assign data_mem_pkt_o[89] = lce_data_cmd_i[89];
  assign data_mem_pkt_o[88] = lce_data_cmd_i[88];
  assign data_mem_pkt_o[87] = lce_data_cmd_i[87];
  assign data_mem_pkt_o[86] = lce_data_cmd_i[86];
  assign data_mem_pkt_o[85] = lce_data_cmd_i[85];
  assign data_mem_pkt_o[84] = lce_data_cmd_i[84];
  assign data_mem_pkt_o[83] = lce_data_cmd_i[83];
  assign data_mem_pkt_o[82] = lce_data_cmd_i[82];
  assign data_mem_pkt_o[81] = lce_data_cmd_i[81];
  assign data_mem_pkt_o[80] = lce_data_cmd_i[80];
  assign data_mem_pkt_o[79] = lce_data_cmd_i[79];
  assign data_mem_pkt_o[78] = lce_data_cmd_i[78];
  assign data_mem_pkt_o[77] = lce_data_cmd_i[77];
  assign data_mem_pkt_o[76] = lce_data_cmd_i[76];
  assign data_mem_pkt_o[75] = lce_data_cmd_i[75];
  assign data_mem_pkt_o[74] = lce_data_cmd_i[74];
  assign data_mem_pkt_o[73] = lce_data_cmd_i[73];
  assign data_mem_pkt_o[72] = lce_data_cmd_i[72];
  assign data_mem_pkt_o[71] = lce_data_cmd_i[71];
  assign data_mem_pkt_o[70] = lce_data_cmd_i[70];
  assign data_mem_pkt_o[69] = lce_data_cmd_i[69];
  assign data_mem_pkt_o[68] = lce_data_cmd_i[68];
  assign data_mem_pkt_o[67] = lce_data_cmd_i[67];
  assign data_mem_pkt_o[66] = lce_data_cmd_i[66];
  assign data_mem_pkt_o[65] = lce_data_cmd_i[65];
  assign data_mem_pkt_o[64] = lce_data_cmd_i[64];
  assign data_mem_pkt_o[63] = lce_data_cmd_i[63];
  assign data_mem_pkt_o[62] = lce_data_cmd_i[62];
  assign data_mem_pkt_o[61] = lce_data_cmd_i[61];
  assign data_mem_pkt_o[60] = lce_data_cmd_i[60];
  assign data_mem_pkt_o[59] = lce_data_cmd_i[59];
  assign data_mem_pkt_o[58] = lce_data_cmd_i[58];
  assign data_mem_pkt_o[57] = lce_data_cmd_i[57];
  assign data_mem_pkt_o[56] = lce_data_cmd_i[56];
  assign data_mem_pkt_o[55] = lce_data_cmd_i[55];
  assign data_mem_pkt_o[54] = lce_data_cmd_i[54];
  assign data_mem_pkt_o[53] = lce_data_cmd_i[53];
  assign data_mem_pkt_o[52] = lce_data_cmd_i[52];
  assign data_mem_pkt_o[51] = lce_data_cmd_i[51];
  assign data_mem_pkt_o[50] = lce_data_cmd_i[50];
  assign data_mem_pkt_o[49] = lce_data_cmd_i[49];
  assign data_mem_pkt_o[48] = lce_data_cmd_i[48];
  assign data_mem_pkt_o[47] = lce_data_cmd_i[47];
  assign data_mem_pkt_o[46] = lce_data_cmd_i[46];
  assign data_mem_pkt_o[45] = lce_data_cmd_i[45];
  assign data_mem_pkt_o[44] = lce_data_cmd_i[44];
  assign data_mem_pkt_o[43] = lce_data_cmd_i[43];
  assign data_mem_pkt_o[42] = lce_data_cmd_i[42];
  assign data_mem_pkt_o[41] = lce_data_cmd_i[41];
  assign data_mem_pkt_o[40] = lce_data_cmd_i[40];
  assign data_mem_pkt_o[39] = lce_data_cmd_i[39];
  assign data_mem_pkt_o[38] = lce_data_cmd_i[38];
  assign data_mem_pkt_o[37] = lce_data_cmd_i[37];
  assign data_mem_pkt_o[36] = lce_data_cmd_i[36];
  assign data_mem_pkt_o[35] = lce_data_cmd_i[35];
  assign data_mem_pkt_o[34] = lce_data_cmd_i[34];
  assign data_mem_pkt_o[33] = lce_data_cmd_i[33];
  assign data_mem_pkt_o[32] = lce_data_cmd_i[32];
  assign data_mem_pkt_o[31] = lce_data_cmd_i[31];
  assign data_mem_pkt_o[30] = lce_data_cmd_i[30];
  assign data_mem_pkt_o[29] = lce_data_cmd_i[29];
  assign data_mem_pkt_o[28] = lce_data_cmd_i[28];
  assign data_mem_pkt_o[27] = lce_data_cmd_i[27];
  assign data_mem_pkt_o[26] = lce_data_cmd_i[26];
  assign data_mem_pkt_o[25] = lce_data_cmd_i[25];
  assign data_mem_pkt_o[24] = lce_data_cmd_i[24];
  assign data_mem_pkt_o[23] = lce_data_cmd_i[23];
  assign data_mem_pkt_o[22] = lce_data_cmd_i[22];
  assign data_mem_pkt_o[21] = lce_data_cmd_i[21];
  assign data_mem_pkt_o[20] = lce_data_cmd_i[20];
  assign data_mem_pkt_o[19] = lce_data_cmd_i[19];
  assign data_mem_pkt_o[18] = lce_data_cmd_i[18];
  assign data_mem_pkt_o[17] = lce_data_cmd_i[17];
  assign data_mem_pkt_o[16] = lce_data_cmd_i[16];
  assign data_mem_pkt_o[15] = lce_data_cmd_i[15];
  assign data_mem_pkt_o[14] = lce_data_cmd_i[14];
  assign data_mem_pkt_o[13] = lce_data_cmd_i[13];
  assign data_mem_pkt_o[12] = lce_data_cmd_i[12];
  assign data_mem_pkt_o[11] = lce_data_cmd_i[11];
  assign data_mem_pkt_o[10] = lce_data_cmd_i[10];
  assign data_mem_pkt_o[9] = lce_data_cmd_i[9];
  assign data_mem_pkt_o[8] = lce_data_cmd_i[8];
  assign data_mem_pkt_o[7] = lce_data_cmd_i[7];
  assign data_mem_pkt_o[6] = lce_data_cmd_i[6];
  assign data_mem_pkt_o[5] = lce_data_cmd_i[5];
  assign data_mem_pkt_o[4] = lce_data_cmd_i[4];
  assign data_mem_pkt_o[3] = lce_data_cmd_i[3];
  assign data_mem_pkt_o[2] = lce_data_cmd_i[2];
  assign data_mem_pkt_o[1] = lce_data_cmd_i[1];
  assign data_mem_pkt_o[0] = lce_data_cmd_i[0];
  assign cce_data_received_o = lce_data_cmd_v_i & data_mem_pkt_yumi_i;

endmodule



// module bsg_mem_p539
// (
//   w_clk_i,
//   w_reset_i,
//   w_v_i,
//   w_addr_i,
//   w_data_i,
//   r_v_i,
//   r_addr_i,
//   r_data_o
// );

//   input [0:0] w_addr_i;
//   input [538:0] w_data_i;
//   input [0:0] r_addr_i;
//   output [538:0] r_data_o;
//   input w_clk_i;
//   input w_reset_i;
//   input w_v_i;
//   input r_v_i;
//   wire [538:0] r_data_o;
//   wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;
//   reg [1077:0] mem;
//   assign r_data_o[538] = (N3)? mem[538] : 
//                          (N0)? mem[1077] : 1'b0;
//   assign N0 = r_addr_i[0];
//   assign r_data_o[537] = (N3)? mem[537] : 
//                          (N0)? mem[1076] : 1'b0;
//   assign r_data_o[536] = (N3)? mem[536] : 
//                          (N0)? mem[1075] : 1'b0;
//   assign r_data_o[535] = (N3)? mem[535] : 
//                          (N0)? mem[1074] : 1'b0;
//   assign r_data_o[534] = (N3)? mem[534] : 
//                          (N0)? mem[1073] : 1'b0;
//   assign r_data_o[533] = (N3)? mem[533] : 
//                          (N0)? mem[1072] : 1'b0;
//   assign r_data_o[532] = (N3)? mem[532] : 
//                          (N0)? mem[1071] : 1'b0;
//   assign r_data_o[531] = (N3)? mem[531] : 
//                          (N0)? mem[1070] : 1'b0;
//   assign r_data_o[530] = (N3)? mem[530] : 
//                          (N0)? mem[1069] : 1'b0;
//   assign r_data_o[529] = (N3)? mem[529] : 
//                          (N0)? mem[1068] : 1'b0;
//   assign r_data_o[528] = (N3)? mem[528] : 
//                          (N0)? mem[1067] : 1'b0;
//   assign r_data_o[527] = (N3)? mem[527] : 
//                          (N0)? mem[1066] : 1'b0;
//   assign r_data_o[526] = (N3)? mem[526] : 
//                          (N0)? mem[1065] : 1'b0;
//   assign r_data_o[525] = (N3)? mem[525] : 
//                          (N0)? mem[1064] : 1'b0;
//   assign r_data_o[524] = (N3)? mem[524] : 
//                          (N0)? mem[1063] : 1'b0;
//   assign r_data_o[523] = (N3)? mem[523] : 
//                          (N0)? mem[1062] : 1'b0;
//   assign r_data_o[522] = (N3)? mem[522] : 
//                          (N0)? mem[1061] : 1'b0;
//   assign r_data_o[521] = (N3)? mem[521] : 
//                          (N0)? mem[1060] : 1'b0;
//   assign r_data_o[520] = (N3)? mem[520] : 
//                          (N0)? mem[1059] : 1'b0;
//   assign r_data_o[519] = (N3)? mem[519] : 
//                          (N0)? mem[1058] : 1'b0;
//   assign r_data_o[518] = (N3)? mem[518] : 
//                          (N0)? mem[1057] : 1'b0;
//   assign r_data_o[517] = (N3)? mem[517] : 
//                          (N0)? mem[1056] : 1'b0;
//   assign r_data_o[516] = (N3)? mem[516] : 
//                          (N0)? mem[1055] : 1'b0;
//   assign r_data_o[515] = (N3)? mem[515] : 
//                          (N0)? mem[1054] : 1'b0;
//   assign r_data_o[514] = (N3)? mem[514] : 
//                          (N0)? mem[1053] : 1'b0;
//   assign r_data_o[513] = (N3)? mem[513] : 
//                          (N0)? mem[1052] : 1'b0;
//   assign r_data_o[512] = (N3)? mem[512] : 
//                          (N0)? mem[1051] : 1'b0;
//   assign r_data_o[511] = (N3)? mem[511] : 
//                          (N0)? mem[1050] : 1'b0;
//   assign r_data_o[510] = (N3)? mem[510] : 
//                          (N0)? mem[1049] : 1'b0;
//   assign r_data_o[509] = (N3)? mem[509] : 
//                          (N0)? mem[1048] : 1'b0;
//   assign r_data_o[508] = (N3)? mem[508] : 
//                          (N0)? mem[1047] : 1'b0;
//   assign r_data_o[507] = (N3)? mem[507] : 
//                          (N0)? mem[1046] : 1'b0;
//   assign r_data_o[506] = (N3)? mem[506] : 
//                          (N0)? mem[1045] : 1'b0;
//   assign r_data_o[505] = (N3)? mem[505] : 
//                          (N0)? mem[1044] : 1'b0;
//   assign r_data_o[504] = (N3)? mem[504] : 
//                          (N0)? mem[1043] : 1'b0;
//   assign r_data_o[503] = (N3)? mem[503] : 
//                          (N0)? mem[1042] : 1'b0;
//   assign r_data_o[502] = (N3)? mem[502] : 
//                          (N0)? mem[1041] : 1'b0;
//   assign r_data_o[501] = (N3)? mem[501] : 
//                          (N0)? mem[1040] : 1'b0;
//   assign r_data_o[500] = (N3)? mem[500] : 
//                          (N0)? mem[1039] : 1'b0;
//   assign r_data_o[499] = (N3)? mem[499] : 
//                          (N0)? mem[1038] : 1'b0;
//   assign r_data_o[498] = (N3)? mem[498] : 
//                          (N0)? mem[1037] : 1'b0;
//   assign r_data_o[497] = (N3)? mem[497] : 
//                          (N0)? mem[1036] : 1'b0;
//   assign r_data_o[496] = (N3)? mem[496] : 
//                          (N0)? mem[1035] : 1'b0;
//   assign r_data_o[495] = (N3)? mem[495] : 
//                          (N0)? mem[1034] : 1'b0;
//   assign r_data_o[494] = (N3)? mem[494] : 
//                          (N0)? mem[1033] : 1'b0;
//   assign r_data_o[493] = (N3)? mem[493] : 
//                          (N0)? mem[1032] : 1'b0;
//   assign r_data_o[492] = (N3)? mem[492] : 
//                          (N0)? mem[1031] : 1'b0;
//   assign r_data_o[491] = (N3)? mem[491] : 
//                          (N0)? mem[1030] : 1'b0;
//   assign r_data_o[490] = (N3)? mem[490] : 
//                          (N0)? mem[1029] : 1'b0;
//   assign r_data_o[489] = (N3)? mem[489] : 
//                          (N0)? mem[1028] : 1'b0;
//   assign r_data_o[488] = (N3)? mem[488] : 
//                          (N0)? mem[1027] : 1'b0;
//   assign r_data_o[487] = (N3)? mem[487] : 
//                          (N0)? mem[1026] : 1'b0;
//   assign r_data_o[486] = (N3)? mem[486] : 
//                          (N0)? mem[1025] : 1'b0;
//   assign r_data_o[485] = (N3)? mem[485] : 
//                          (N0)? mem[1024] : 1'b0;
//   assign r_data_o[484] = (N3)? mem[484] : 
//                          (N0)? mem[1023] : 1'b0;
//   assign r_data_o[483] = (N3)? mem[483] : 
//                          (N0)? mem[1022] : 1'b0;
//   assign r_data_o[482] = (N3)? mem[482] : 
//                          (N0)? mem[1021] : 1'b0;
//   assign r_data_o[481] = (N3)? mem[481] : 
//                          (N0)? mem[1020] : 1'b0;
//   assign r_data_o[480] = (N3)? mem[480] : 
//                          (N0)? mem[1019] : 1'b0;
//   assign r_data_o[479] = (N3)? mem[479] : 
//                          (N0)? mem[1018] : 1'b0;
//   assign r_data_o[478] = (N3)? mem[478] : 
//                          (N0)? mem[1017] : 1'b0;
//   assign r_data_o[477] = (N3)? mem[477] : 
//                          (N0)? mem[1016] : 1'b0;
//   assign r_data_o[476] = (N3)? mem[476] : 
//                          (N0)? mem[1015] : 1'b0;
//   assign r_data_o[475] = (N3)? mem[475] : 
//                          (N0)? mem[1014] : 1'b0;
//   assign r_data_o[474] = (N3)? mem[474] : 
//                          (N0)? mem[1013] : 1'b0;
//   assign r_data_o[473] = (N3)? mem[473] : 
//                          (N0)? mem[1012] : 1'b0;
//   assign r_data_o[472] = (N3)? mem[472] : 
//                          (N0)? mem[1011] : 1'b0;
//   assign r_data_o[471] = (N3)? mem[471] : 
//                          (N0)? mem[1010] : 1'b0;
//   assign r_data_o[470] = (N3)? mem[470] : 
//                          (N0)? mem[1009] : 1'b0;
//   assign r_data_o[469] = (N3)? mem[469] : 
//                          (N0)? mem[1008] : 1'b0;
//   assign r_data_o[468] = (N3)? mem[468] : 
//                          (N0)? mem[1007] : 1'b0;
//   assign r_data_o[467] = (N3)? mem[467] : 
//                          (N0)? mem[1006] : 1'b0;
//   assign r_data_o[466] = (N3)? mem[466] : 
//                          (N0)? mem[1005] : 1'b0;
//   assign r_data_o[465] = (N3)? mem[465] : 
//                          (N0)? mem[1004] : 1'b0;
//   assign r_data_o[464] = (N3)? mem[464] : 
//                          (N0)? mem[1003] : 1'b0;
//   assign r_data_o[463] = (N3)? mem[463] : 
//                          (N0)? mem[1002] : 1'b0;
//   assign r_data_o[462] = (N3)? mem[462] : 
//                          (N0)? mem[1001] : 1'b0;
//   assign r_data_o[461] = (N3)? mem[461] : 
//                          (N0)? mem[1000] : 1'b0;
//   assign r_data_o[460] = (N3)? mem[460] : 
//                          (N0)? mem[999] : 1'b0;
//   assign r_data_o[459] = (N3)? mem[459] : 
//                          (N0)? mem[998] : 1'b0;
//   assign r_data_o[458] = (N3)? mem[458] : 
//                          (N0)? mem[997] : 1'b0;
//   assign r_data_o[457] = (N3)? mem[457] : 
//                          (N0)? mem[996] : 1'b0;
//   assign r_data_o[456] = (N3)? mem[456] : 
//                          (N0)? mem[995] : 1'b0;
//   assign r_data_o[455] = (N3)? mem[455] : 
//                          (N0)? mem[994] : 1'b0;
//   assign r_data_o[454] = (N3)? mem[454] : 
//                          (N0)? mem[993] : 1'b0;
//   assign r_data_o[453] = (N3)? mem[453] : 
//                          (N0)? mem[992] : 1'b0;
//   assign r_data_o[452] = (N3)? mem[452] : 
//                          (N0)? mem[991] : 1'b0;
//   assign r_data_o[451] = (N3)? mem[451] : 
//                          (N0)? mem[990] : 1'b0;
//   assign r_data_o[450] = (N3)? mem[450] : 
//                          (N0)? mem[989] : 1'b0;
//   assign r_data_o[449] = (N3)? mem[449] : 
//                          (N0)? mem[988] : 1'b0;
//   assign r_data_o[448] = (N3)? mem[448] : 
//                          (N0)? mem[987] : 1'b0;
//   assign r_data_o[447] = (N3)? mem[447] : 
//                          (N0)? mem[986] : 1'b0;
//   assign r_data_o[446] = (N3)? mem[446] : 
//                          (N0)? mem[985] : 1'b0;
//   assign r_data_o[445] = (N3)? mem[445] : 
//                          (N0)? mem[984] : 1'b0;
//   assign r_data_o[444] = (N3)? mem[444] : 
//                          (N0)? mem[983] : 1'b0;
//   assign r_data_o[443] = (N3)? mem[443] : 
//                          (N0)? mem[982] : 1'b0;
//   assign r_data_o[442] = (N3)? mem[442] : 
//                          (N0)? mem[981] : 1'b0;
//   assign r_data_o[441] = (N3)? mem[441] : 
//                          (N0)? mem[980] : 1'b0;
//   assign r_data_o[440] = (N3)? mem[440] : 
//                          (N0)? mem[979] : 1'b0;
//   assign r_data_o[439] = (N3)? mem[439] : 
//                          (N0)? mem[978] : 1'b0;
//   assign r_data_o[438] = (N3)? mem[438] : 
//                          (N0)? mem[977] : 1'b0;
//   assign r_data_o[437] = (N3)? mem[437] : 
//                          (N0)? mem[976] : 1'b0;
//   assign r_data_o[436] = (N3)? mem[436] : 
//                          (N0)? mem[975] : 1'b0;
//   assign r_data_o[435] = (N3)? mem[435] : 
//                          (N0)? mem[974] : 1'b0;
//   assign r_data_o[434] = (N3)? mem[434] : 
//                          (N0)? mem[973] : 1'b0;
//   assign r_data_o[433] = (N3)? mem[433] : 
//                          (N0)? mem[972] : 1'b0;
//   assign r_data_o[432] = (N3)? mem[432] : 
//                          (N0)? mem[971] : 1'b0;
//   assign r_data_o[431] = (N3)? mem[431] : 
//                          (N0)? mem[970] : 1'b0;
//   assign r_data_o[430] = (N3)? mem[430] : 
//                          (N0)? mem[969] : 1'b0;
//   assign r_data_o[429] = (N3)? mem[429] : 
//                          (N0)? mem[968] : 1'b0;
//   assign r_data_o[428] = (N3)? mem[428] : 
//                          (N0)? mem[967] : 1'b0;
//   assign r_data_o[427] = (N3)? mem[427] : 
//                          (N0)? mem[966] : 1'b0;
//   assign r_data_o[426] = (N3)? mem[426] : 
//                          (N0)? mem[965] : 1'b0;
//   assign r_data_o[425] = (N3)? mem[425] : 
//                          (N0)? mem[964] : 1'b0;
//   assign r_data_o[424] = (N3)? mem[424] : 
//                          (N0)? mem[963] : 1'b0;
//   assign r_data_o[423] = (N3)? mem[423] : 
//                          (N0)? mem[962] : 1'b0;
//   assign r_data_o[422] = (N3)? mem[422] : 
//                          (N0)? mem[961] : 1'b0;
//   assign r_data_o[421] = (N3)? mem[421] : 
//                          (N0)? mem[960] : 1'b0;
//   assign r_data_o[420] = (N3)? mem[420] : 
//                          (N0)? mem[959] : 1'b0;
//   assign r_data_o[419] = (N3)? mem[419] : 
//                          (N0)? mem[958] : 1'b0;
//   assign r_data_o[418] = (N3)? mem[418] : 
//                          (N0)? mem[957] : 1'b0;
//   assign r_data_o[417] = (N3)? mem[417] : 
//                          (N0)? mem[956] : 1'b0;
//   assign r_data_o[416] = (N3)? mem[416] : 
//                          (N0)? mem[955] : 1'b0;
//   assign r_data_o[415] = (N3)? mem[415] : 
//                          (N0)? mem[954] : 1'b0;
//   assign r_data_o[414] = (N3)? mem[414] : 
//                          (N0)? mem[953] : 1'b0;
//   assign r_data_o[413] = (N3)? mem[413] : 
//                          (N0)? mem[952] : 1'b0;
//   assign r_data_o[412] = (N3)? mem[412] : 
//                          (N0)? mem[951] : 1'b0;
//   assign r_data_o[411] = (N3)? mem[411] : 
//                          (N0)? mem[950] : 1'b0;
//   assign r_data_o[410] = (N3)? mem[410] : 
//                          (N0)? mem[949] : 1'b0;
//   assign r_data_o[409] = (N3)? mem[409] : 
//                          (N0)? mem[948] : 1'b0;
//   assign r_data_o[408] = (N3)? mem[408] : 
//                          (N0)? mem[947] : 1'b0;
//   assign r_data_o[407] = (N3)? mem[407] : 
//                          (N0)? mem[946] : 1'b0;
//   assign r_data_o[406] = (N3)? mem[406] : 
//                          (N0)? mem[945] : 1'b0;
//   assign r_data_o[405] = (N3)? mem[405] : 
//                          (N0)? mem[944] : 1'b0;
//   assign r_data_o[404] = (N3)? mem[404] : 
//                          (N0)? mem[943] : 1'b0;
//   assign r_data_o[403] = (N3)? mem[403] : 
//                          (N0)? mem[942] : 1'b0;
//   assign r_data_o[402] = (N3)? mem[402] : 
//                          (N0)? mem[941] : 1'b0;
//   assign r_data_o[401] = (N3)? mem[401] : 
//                          (N0)? mem[940] : 1'b0;
//   assign r_data_o[400] = (N3)? mem[400] : 
//                          (N0)? mem[939] : 1'b0;
//   assign r_data_o[399] = (N3)? mem[399] : 
//                          (N0)? mem[938] : 1'b0;
//   assign r_data_o[398] = (N3)? mem[398] : 
//                          (N0)? mem[937] : 1'b0;
//   assign r_data_o[397] = (N3)? mem[397] : 
//                          (N0)? mem[936] : 1'b0;
//   assign r_data_o[396] = (N3)? mem[396] : 
//                          (N0)? mem[935] : 1'b0;
//   assign r_data_o[395] = (N3)? mem[395] : 
//                          (N0)? mem[934] : 1'b0;
//   assign r_data_o[394] = (N3)? mem[394] : 
//                          (N0)? mem[933] : 1'b0;
//   assign r_data_o[393] = (N3)? mem[393] : 
//                          (N0)? mem[932] : 1'b0;
//   assign r_data_o[392] = (N3)? mem[392] : 
//                          (N0)? mem[931] : 1'b0;
//   assign r_data_o[391] = (N3)? mem[391] : 
//                          (N0)? mem[930] : 1'b0;
//   assign r_data_o[390] = (N3)? mem[390] : 
//                          (N0)? mem[929] : 1'b0;
//   assign r_data_o[389] = (N3)? mem[389] : 
//                          (N0)? mem[928] : 1'b0;
//   assign r_data_o[388] = (N3)? mem[388] : 
//                          (N0)? mem[927] : 1'b0;
//   assign r_data_o[387] = (N3)? mem[387] : 
//                          (N0)? mem[926] : 1'b0;
//   assign r_data_o[386] = (N3)? mem[386] : 
//                          (N0)? mem[925] : 1'b0;
//   assign r_data_o[385] = (N3)? mem[385] : 
//                          (N0)? mem[924] : 1'b0;
//   assign r_data_o[384] = (N3)? mem[384] : 
//                          (N0)? mem[923] : 1'b0;
//   assign r_data_o[383] = (N3)? mem[383] : 
//                          (N0)? mem[922] : 1'b0;
//   assign r_data_o[382] = (N3)? mem[382] : 
//                          (N0)? mem[921] : 1'b0;
//   assign r_data_o[381] = (N3)? mem[381] : 
//                          (N0)? mem[920] : 1'b0;
//   assign r_data_o[380] = (N3)? mem[380] : 
//                          (N0)? mem[919] : 1'b0;
//   assign r_data_o[379] = (N3)? mem[379] : 
//                          (N0)? mem[918] : 1'b0;
//   assign r_data_o[378] = (N3)? mem[378] : 
//                          (N0)? mem[917] : 1'b0;
//   assign r_data_o[377] = (N3)? mem[377] : 
//                          (N0)? mem[916] : 1'b0;
//   assign r_data_o[376] = (N3)? mem[376] : 
//                          (N0)? mem[915] : 1'b0;
//   assign r_data_o[375] = (N3)? mem[375] : 
//                          (N0)? mem[914] : 1'b0;
//   assign r_data_o[374] = (N3)? mem[374] : 
//                          (N0)? mem[913] : 1'b0;
//   assign r_data_o[373] = (N3)? mem[373] : 
//                          (N0)? mem[912] : 1'b0;
//   assign r_data_o[372] = (N3)? mem[372] : 
//                          (N0)? mem[911] : 1'b0;
//   assign r_data_o[371] = (N3)? mem[371] : 
//                          (N0)? mem[910] : 1'b0;
//   assign r_data_o[370] = (N3)? mem[370] : 
//                          (N0)? mem[909] : 1'b0;
//   assign r_data_o[369] = (N3)? mem[369] : 
//                          (N0)? mem[908] : 1'b0;
//   assign r_data_o[368] = (N3)? mem[368] : 
//                          (N0)? mem[907] : 1'b0;
//   assign r_data_o[367] = (N3)? mem[367] : 
//                          (N0)? mem[906] : 1'b0;
//   assign r_data_o[366] = (N3)? mem[366] : 
//                          (N0)? mem[905] : 1'b0;
//   assign r_data_o[365] = (N3)? mem[365] : 
//                          (N0)? mem[904] : 1'b0;
//   assign r_data_o[364] = (N3)? mem[364] : 
//                          (N0)? mem[903] : 1'b0;
//   assign r_data_o[363] = (N3)? mem[363] : 
//                          (N0)? mem[902] : 1'b0;
//   assign r_data_o[362] = (N3)? mem[362] : 
//                          (N0)? mem[901] : 1'b0;
//   assign r_data_o[361] = (N3)? mem[361] : 
//                          (N0)? mem[900] : 1'b0;
//   assign r_data_o[360] = (N3)? mem[360] : 
//                          (N0)? mem[899] : 1'b0;
//   assign r_data_o[359] = (N3)? mem[359] : 
//                          (N0)? mem[898] : 1'b0;
//   assign r_data_o[358] = (N3)? mem[358] : 
//                          (N0)? mem[897] : 1'b0;
//   assign r_data_o[357] = (N3)? mem[357] : 
//                          (N0)? mem[896] : 1'b0;
//   assign r_data_o[356] = (N3)? mem[356] : 
//                          (N0)? mem[895] : 1'b0;
//   assign r_data_o[355] = (N3)? mem[355] : 
//                          (N0)? mem[894] : 1'b0;
//   assign r_data_o[354] = (N3)? mem[354] : 
//                          (N0)? mem[893] : 1'b0;
//   assign r_data_o[353] = (N3)? mem[353] : 
//                          (N0)? mem[892] : 1'b0;
//   assign r_data_o[352] = (N3)? mem[352] : 
//                          (N0)? mem[891] : 1'b0;
//   assign r_data_o[351] = (N3)? mem[351] : 
//                          (N0)? mem[890] : 1'b0;
//   assign r_data_o[350] = (N3)? mem[350] : 
//                          (N0)? mem[889] : 1'b0;
//   assign r_data_o[349] = (N3)? mem[349] : 
//                          (N0)? mem[888] : 1'b0;
//   assign r_data_o[348] = (N3)? mem[348] : 
//                          (N0)? mem[887] : 1'b0;
//   assign r_data_o[347] = (N3)? mem[347] : 
//                          (N0)? mem[886] : 1'b0;
//   assign r_data_o[346] = (N3)? mem[346] : 
//                          (N0)? mem[885] : 1'b0;
//   assign r_data_o[345] = (N3)? mem[345] : 
//                          (N0)? mem[884] : 1'b0;
//   assign r_data_o[344] = (N3)? mem[344] : 
//                          (N0)? mem[883] : 1'b0;
//   assign r_data_o[343] = (N3)? mem[343] : 
//                          (N0)? mem[882] : 1'b0;
//   assign r_data_o[342] = (N3)? mem[342] : 
//                          (N0)? mem[881] : 1'b0;
//   assign r_data_o[341] = (N3)? mem[341] : 
//                          (N0)? mem[880] : 1'b0;
//   assign r_data_o[340] = (N3)? mem[340] : 
//                          (N0)? mem[879] : 1'b0;
//   assign r_data_o[339] = (N3)? mem[339] : 
//                          (N0)? mem[878] : 1'b0;
//   assign r_data_o[338] = (N3)? mem[338] : 
//                          (N0)? mem[877] : 1'b0;
//   assign r_data_o[337] = (N3)? mem[337] : 
//                          (N0)? mem[876] : 1'b0;
//   assign r_data_o[336] = (N3)? mem[336] : 
//                          (N0)? mem[875] : 1'b0;
//   assign r_data_o[335] = (N3)? mem[335] : 
//                          (N0)? mem[874] : 1'b0;
//   assign r_data_o[334] = (N3)? mem[334] : 
//                          (N0)? mem[873] : 1'b0;
//   assign r_data_o[333] = (N3)? mem[333] : 
//                          (N0)? mem[872] : 1'b0;
//   assign r_data_o[332] = (N3)? mem[332] : 
//                          (N0)? mem[871] : 1'b0;
//   assign r_data_o[331] = (N3)? mem[331] : 
//                          (N0)? mem[870] : 1'b0;
//   assign r_data_o[330] = (N3)? mem[330] : 
//                          (N0)? mem[869] : 1'b0;
//   assign r_data_o[329] = (N3)? mem[329] : 
//                          (N0)? mem[868] : 1'b0;
//   assign r_data_o[328] = (N3)? mem[328] : 
//                          (N0)? mem[867] : 1'b0;
//   assign r_data_o[327] = (N3)? mem[327] : 
//                          (N0)? mem[866] : 1'b0;
//   assign r_data_o[326] = (N3)? mem[326] : 
//                          (N0)? mem[865] : 1'b0;
//   assign r_data_o[325] = (N3)? mem[325] : 
//                          (N0)? mem[864] : 1'b0;
//   assign r_data_o[324] = (N3)? mem[324] : 
//                          (N0)? mem[863] : 1'b0;
//   assign r_data_o[323] = (N3)? mem[323] : 
//                          (N0)? mem[862] : 1'b0;
//   assign r_data_o[322] = (N3)? mem[322] : 
//                          (N0)? mem[861] : 1'b0;
//   assign r_data_o[321] = (N3)? mem[321] : 
//                          (N0)? mem[860] : 1'b0;
//   assign r_data_o[320] = (N3)? mem[320] : 
//                          (N0)? mem[859] : 1'b0;
//   assign r_data_o[319] = (N3)? mem[319] : 
//                          (N0)? mem[858] : 1'b0;
//   assign r_data_o[318] = (N3)? mem[318] : 
//                          (N0)? mem[857] : 1'b0;
//   assign r_data_o[317] = (N3)? mem[317] : 
//                          (N0)? mem[856] : 1'b0;
//   assign r_data_o[316] = (N3)? mem[316] : 
//                          (N0)? mem[855] : 1'b0;
//   assign r_data_o[315] = (N3)? mem[315] : 
//                          (N0)? mem[854] : 1'b0;
//   assign r_data_o[314] = (N3)? mem[314] : 
//                          (N0)? mem[853] : 1'b0;
//   assign r_data_o[313] = (N3)? mem[313] : 
//                          (N0)? mem[852] : 1'b0;
//   assign r_data_o[312] = (N3)? mem[312] : 
//                          (N0)? mem[851] : 1'b0;
//   assign r_data_o[311] = (N3)? mem[311] : 
//                          (N0)? mem[850] : 1'b0;
//   assign r_data_o[310] = (N3)? mem[310] : 
//                          (N0)? mem[849] : 1'b0;
//   assign r_data_o[309] = (N3)? mem[309] : 
//                          (N0)? mem[848] : 1'b0;
//   assign r_data_o[308] = (N3)? mem[308] : 
//                          (N0)? mem[847] : 1'b0;
//   assign r_data_o[307] = (N3)? mem[307] : 
//                          (N0)? mem[846] : 1'b0;
//   assign r_data_o[306] = (N3)? mem[306] : 
//                          (N0)? mem[845] : 1'b0;
//   assign r_data_o[305] = (N3)? mem[305] : 
//                          (N0)? mem[844] : 1'b0;
//   assign r_data_o[304] = (N3)? mem[304] : 
//                          (N0)? mem[843] : 1'b0;
//   assign r_data_o[303] = (N3)? mem[303] : 
//                          (N0)? mem[842] : 1'b0;
//   assign r_data_o[302] = (N3)? mem[302] : 
//                          (N0)? mem[841] : 1'b0;
//   assign r_data_o[301] = (N3)? mem[301] : 
//                          (N0)? mem[840] : 1'b0;
//   assign r_data_o[300] = (N3)? mem[300] : 
//                          (N0)? mem[839] : 1'b0;
//   assign r_data_o[299] = (N3)? mem[299] : 
//                          (N0)? mem[838] : 1'b0;
//   assign r_data_o[298] = (N3)? mem[298] : 
//                          (N0)? mem[837] : 1'b0;
//   assign r_data_o[297] = (N3)? mem[297] : 
//                          (N0)? mem[836] : 1'b0;
//   assign r_data_o[296] = (N3)? mem[296] : 
//                          (N0)? mem[835] : 1'b0;
//   assign r_data_o[295] = (N3)? mem[295] : 
//                          (N0)? mem[834] : 1'b0;
//   assign r_data_o[294] = (N3)? mem[294] : 
//                          (N0)? mem[833] : 1'b0;
//   assign r_data_o[293] = (N3)? mem[293] : 
//                          (N0)? mem[832] : 1'b0;
//   assign r_data_o[292] = (N3)? mem[292] : 
//                          (N0)? mem[831] : 1'b0;
//   assign r_data_o[291] = (N3)? mem[291] : 
//                          (N0)? mem[830] : 1'b0;
//   assign r_data_o[290] = (N3)? mem[290] : 
//                          (N0)? mem[829] : 1'b0;
//   assign r_data_o[289] = (N3)? mem[289] : 
//                          (N0)? mem[828] : 1'b0;
//   assign r_data_o[288] = (N3)? mem[288] : 
//                          (N0)? mem[827] : 1'b0;
//   assign r_data_o[287] = (N3)? mem[287] : 
//                          (N0)? mem[826] : 1'b0;
//   assign r_data_o[286] = (N3)? mem[286] : 
//                          (N0)? mem[825] : 1'b0;
//   assign r_data_o[285] = (N3)? mem[285] : 
//                          (N0)? mem[824] : 1'b0;
//   assign r_data_o[284] = (N3)? mem[284] : 
//                          (N0)? mem[823] : 1'b0;
//   assign r_data_o[283] = (N3)? mem[283] : 
//                          (N0)? mem[822] : 1'b0;
//   assign r_data_o[282] = (N3)? mem[282] : 
//                          (N0)? mem[821] : 1'b0;
//   assign r_data_o[281] = (N3)? mem[281] : 
//                          (N0)? mem[820] : 1'b0;
//   assign r_data_o[280] = (N3)? mem[280] : 
//                          (N0)? mem[819] : 1'b0;
//   assign r_data_o[279] = (N3)? mem[279] : 
//                          (N0)? mem[818] : 1'b0;
//   assign r_data_o[278] = (N3)? mem[278] : 
//                          (N0)? mem[817] : 1'b0;
//   assign r_data_o[277] = (N3)? mem[277] : 
//                          (N0)? mem[816] : 1'b0;
//   assign r_data_o[276] = (N3)? mem[276] : 
//                          (N0)? mem[815] : 1'b0;
//   assign r_data_o[275] = (N3)? mem[275] : 
//                          (N0)? mem[814] : 1'b0;
//   assign r_data_o[274] = (N3)? mem[274] : 
//                          (N0)? mem[813] : 1'b0;
//   assign r_data_o[273] = (N3)? mem[273] : 
//                          (N0)? mem[812] : 1'b0;
//   assign r_data_o[272] = (N3)? mem[272] : 
//                          (N0)? mem[811] : 1'b0;
//   assign r_data_o[271] = (N3)? mem[271] : 
//                          (N0)? mem[810] : 1'b0;
//   assign r_data_o[270] = (N3)? mem[270] : 
//                          (N0)? mem[809] : 1'b0;
//   assign r_data_o[269] = (N3)? mem[269] : 
//                          (N0)? mem[808] : 1'b0;
//   assign r_data_o[268] = (N3)? mem[268] : 
//                          (N0)? mem[807] : 1'b0;
//   assign r_data_o[267] = (N3)? mem[267] : 
//                          (N0)? mem[806] : 1'b0;
//   assign r_data_o[266] = (N3)? mem[266] : 
//                          (N0)? mem[805] : 1'b0;
//   assign r_data_o[265] = (N3)? mem[265] : 
//                          (N0)? mem[804] : 1'b0;
//   assign r_data_o[264] = (N3)? mem[264] : 
//                          (N0)? mem[803] : 1'b0;
//   assign r_data_o[263] = (N3)? mem[263] : 
//                          (N0)? mem[802] : 1'b0;
//   assign r_data_o[262] = (N3)? mem[262] : 
//                          (N0)? mem[801] : 1'b0;
//   assign r_data_o[261] = (N3)? mem[261] : 
//                          (N0)? mem[800] : 1'b0;
//   assign r_data_o[260] = (N3)? mem[260] : 
//                          (N0)? mem[799] : 1'b0;
//   assign r_data_o[259] = (N3)? mem[259] : 
//                          (N0)? mem[798] : 1'b0;
//   assign r_data_o[258] = (N3)? mem[258] : 
//                          (N0)? mem[797] : 1'b0;
//   assign r_data_o[257] = (N3)? mem[257] : 
//                          (N0)? mem[796] : 1'b0;
//   assign r_data_o[256] = (N3)? mem[256] : 
//                          (N0)? mem[795] : 1'b0;
//   assign r_data_o[255] = (N3)? mem[255] : 
//                          (N0)? mem[794] : 1'b0;
//   assign r_data_o[254] = (N3)? mem[254] : 
//                          (N0)? mem[793] : 1'b0;
//   assign r_data_o[253] = (N3)? mem[253] : 
//                          (N0)? mem[792] : 1'b0;
//   assign r_data_o[252] = (N3)? mem[252] : 
//                          (N0)? mem[791] : 1'b0;
//   assign r_data_o[251] = (N3)? mem[251] : 
//                          (N0)? mem[790] : 1'b0;
//   assign r_data_o[250] = (N3)? mem[250] : 
//                          (N0)? mem[789] : 1'b0;
//   assign r_data_o[249] = (N3)? mem[249] : 
//                          (N0)? mem[788] : 1'b0;
//   assign r_data_o[248] = (N3)? mem[248] : 
//                          (N0)? mem[787] : 1'b0;
//   assign r_data_o[247] = (N3)? mem[247] : 
//                          (N0)? mem[786] : 1'b0;
//   assign r_data_o[246] = (N3)? mem[246] : 
//                          (N0)? mem[785] : 1'b0;
//   assign r_data_o[245] = (N3)? mem[245] : 
//                          (N0)? mem[784] : 1'b0;
//   assign r_data_o[244] = (N3)? mem[244] : 
//                          (N0)? mem[783] : 1'b0;
//   assign r_data_o[243] = (N3)? mem[243] : 
//                          (N0)? mem[782] : 1'b0;
//   assign r_data_o[242] = (N3)? mem[242] : 
//                          (N0)? mem[781] : 1'b0;
//   assign r_data_o[241] = (N3)? mem[241] : 
//                          (N0)? mem[780] : 1'b0;
//   assign r_data_o[240] = (N3)? mem[240] : 
//                          (N0)? mem[779] : 1'b0;
//   assign r_data_o[239] = (N3)? mem[239] : 
//                          (N0)? mem[778] : 1'b0;
//   assign r_data_o[238] = (N3)? mem[238] : 
//                          (N0)? mem[777] : 1'b0;
//   assign r_data_o[237] = (N3)? mem[237] : 
//                          (N0)? mem[776] : 1'b0;
//   assign r_data_o[236] = (N3)? mem[236] : 
//                          (N0)? mem[775] : 1'b0;
//   assign r_data_o[235] = (N3)? mem[235] : 
//                          (N0)? mem[774] : 1'b0;
//   assign r_data_o[234] = (N3)? mem[234] : 
//                          (N0)? mem[773] : 1'b0;
//   assign r_data_o[233] = (N3)? mem[233] : 
//                          (N0)? mem[772] : 1'b0;
//   assign r_data_o[232] = (N3)? mem[232] : 
//                          (N0)? mem[771] : 1'b0;
//   assign r_data_o[231] = (N3)? mem[231] : 
//                          (N0)? mem[770] : 1'b0;
//   assign r_data_o[230] = (N3)? mem[230] : 
//                          (N0)? mem[769] : 1'b0;
//   assign r_data_o[229] = (N3)? mem[229] : 
//                          (N0)? mem[768] : 1'b0;
//   assign r_data_o[228] = (N3)? mem[228] : 
//                          (N0)? mem[767] : 1'b0;
//   assign r_data_o[227] = (N3)? mem[227] : 
//                          (N0)? mem[766] : 1'b0;
//   assign r_data_o[226] = (N3)? mem[226] : 
//                          (N0)? mem[765] : 1'b0;
//   assign r_data_o[225] = (N3)? mem[225] : 
//                          (N0)? mem[764] : 1'b0;
//   assign r_data_o[224] = (N3)? mem[224] : 
//                          (N0)? mem[763] : 1'b0;
//   assign r_data_o[223] = (N3)? mem[223] : 
//                          (N0)? mem[762] : 1'b0;
//   assign r_data_o[222] = (N3)? mem[222] : 
//                          (N0)? mem[761] : 1'b0;
//   assign r_data_o[221] = (N3)? mem[221] : 
//                          (N0)? mem[760] : 1'b0;
//   assign r_data_o[220] = (N3)? mem[220] : 
//                          (N0)? mem[759] : 1'b0;
//   assign r_data_o[219] = (N3)? mem[219] : 
//                          (N0)? mem[758] : 1'b0;
//   assign r_data_o[218] = (N3)? mem[218] : 
//                          (N0)? mem[757] : 1'b0;
//   assign r_data_o[217] = (N3)? mem[217] : 
//                          (N0)? mem[756] : 1'b0;
//   assign r_data_o[216] = (N3)? mem[216] : 
//                          (N0)? mem[755] : 1'b0;
//   assign r_data_o[215] = (N3)? mem[215] : 
//                          (N0)? mem[754] : 1'b0;
//   assign r_data_o[214] = (N3)? mem[214] : 
//                          (N0)? mem[753] : 1'b0;
//   assign r_data_o[213] = (N3)? mem[213] : 
//                          (N0)? mem[752] : 1'b0;
//   assign r_data_o[212] = (N3)? mem[212] : 
//                          (N0)? mem[751] : 1'b0;
//   assign r_data_o[211] = (N3)? mem[211] : 
//                          (N0)? mem[750] : 1'b0;
//   assign r_data_o[210] = (N3)? mem[210] : 
//                          (N0)? mem[749] : 1'b0;
//   assign r_data_o[209] = (N3)? mem[209] : 
//                          (N0)? mem[748] : 1'b0;
//   assign r_data_o[208] = (N3)? mem[208] : 
//                          (N0)? mem[747] : 1'b0;
//   assign r_data_o[207] = (N3)? mem[207] : 
//                          (N0)? mem[746] : 1'b0;
//   assign r_data_o[206] = (N3)? mem[206] : 
//                          (N0)? mem[745] : 1'b0;
//   assign r_data_o[205] = (N3)? mem[205] : 
//                          (N0)? mem[744] : 1'b0;
//   assign r_data_o[204] = (N3)? mem[204] : 
//                          (N0)? mem[743] : 1'b0;
//   assign r_data_o[203] = (N3)? mem[203] : 
//                          (N0)? mem[742] : 1'b0;
//   assign r_data_o[202] = (N3)? mem[202] : 
//                          (N0)? mem[741] : 1'b0;
//   assign r_data_o[201] = (N3)? mem[201] : 
//                          (N0)? mem[740] : 1'b0;
//   assign r_data_o[200] = (N3)? mem[200] : 
//                          (N0)? mem[739] : 1'b0;
//   assign r_data_o[199] = (N3)? mem[199] : 
//                          (N0)? mem[738] : 1'b0;
//   assign r_data_o[198] = (N3)? mem[198] : 
//                          (N0)? mem[737] : 1'b0;
//   assign r_data_o[197] = (N3)? mem[197] : 
//                          (N0)? mem[736] : 1'b0;
//   assign r_data_o[196] = (N3)? mem[196] : 
//                          (N0)? mem[735] : 1'b0;
//   assign r_data_o[195] = (N3)? mem[195] : 
//                          (N0)? mem[734] : 1'b0;
//   assign r_data_o[194] = (N3)? mem[194] : 
//                          (N0)? mem[733] : 1'b0;
//   assign r_data_o[193] = (N3)? mem[193] : 
//                          (N0)? mem[732] : 1'b0;
//   assign r_data_o[192] = (N3)? mem[192] : 
//                          (N0)? mem[731] : 1'b0;
//   assign r_data_o[191] = (N3)? mem[191] : 
//                          (N0)? mem[730] : 1'b0;
//   assign r_data_o[190] = (N3)? mem[190] : 
//                          (N0)? mem[729] : 1'b0;
//   assign r_data_o[189] = (N3)? mem[189] : 
//                          (N0)? mem[728] : 1'b0;
//   assign r_data_o[188] = (N3)? mem[188] : 
//                          (N0)? mem[727] : 1'b0;
//   assign r_data_o[187] = (N3)? mem[187] : 
//                          (N0)? mem[726] : 1'b0;
//   assign r_data_o[186] = (N3)? mem[186] : 
//                          (N0)? mem[725] : 1'b0;
//   assign r_data_o[185] = (N3)? mem[185] : 
//                          (N0)? mem[724] : 1'b0;
//   assign r_data_o[184] = (N3)? mem[184] : 
//                          (N0)? mem[723] : 1'b0;
//   assign r_data_o[183] = (N3)? mem[183] : 
//                          (N0)? mem[722] : 1'b0;
//   assign r_data_o[182] = (N3)? mem[182] : 
//                          (N0)? mem[721] : 1'b0;
//   assign r_data_o[181] = (N3)? mem[181] : 
//                          (N0)? mem[720] : 1'b0;
//   assign r_data_o[180] = (N3)? mem[180] : 
//                          (N0)? mem[719] : 1'b0;
//   assign r_data_o[179] = (N3)? mem[179] : 
//                          (N0)? mem[718] : 1'b0;
//   assign r_data_o[178] = (N3)? mem[178] : 
//                          (N0)? mem[717] : 1'b0;
//   assign r_data_o[177] = (N3)? mem[177] : 
//                          (N0)? mem[716] : 1'b0;
//   assign r_data_o[176] = (N3)? mem[176] : 
//                          (N0)? mem[715] : 1'b0;
//   assign r_data_o[175] = (N3)? mem[175] : 
//                          (N0)? mem[714] : 1'b0;
//   assign r_data_o[174] = (N3)? mem[174] : 
//                          (N0)? mem[713] : 1'b0;
//   assign r_data_o[173] = (N3)? mem[173] : 
//                          (N0)? mem[712] : 1'b0;
//   assign r_data_o[172] = (N3)? mem[172] : 
//                          (N0)? mem[711] : 1'b0;
//   assign r_data_o[171] = (N3)? mem[171] : 
//                          (N0)? mem[710] : 1'b0;
//   assign r_data_o[170] = (N3)? mem[170] : 
//                          (N0)? mem[709] : 1'b0;
//   assign r_data_o[169] = (N3)? mem[169] : 
//                          (N0)? mem[708] : 1'b0;
//   assign r_data_o[168] = (N3)? mem[168] : 
//                          (N0)? mem[707] : 1'b0;
//   assign r_data_o[167] = (N3)? mem[167] : 
//                          (N0)? mem[706] : 1'b0;
//   assign r_data_o[166] = (N3)? mem[166] : 
//                          (N0)? mem[705] : 1'b0;
//   assign r_data_o[165] = (N3)? mem[165] : 
//                          (N0)? mem[704] : 1'b0;
//   assign r_data_o[164] = (N3)? mem[164] : 
//                          (N0)? mem[703] : 1'b0;
//   assign r_data_o[163] = (N3)? mem[163] : 
//                          (N0)? mem[702] : 1'b0;
//   assign r_data_o[162] = (N3)? mem[162] : 
//                          (N0)? mem[701] : 1'b0;
//   assign r_data_o[161] = (N3)? mem[161] : 
//                          (N0)? mem[700] : 1'b0;
//   assign r_data_o[160] = (N3)? mem[160] : 
//                          (N0)? mem[699] : 1'b0;
//   assign r_data_o[159] = (N3)? mem[159] : 
//                          (N0)? mem[698] : 1'b0;
//   assign r_data_o[158] = (N3)? mem[158] : 
//                          (N0)? mem[697] : 1'b0;
//   assign r_data_o[157] = (N3)? mem[157] : 
//                          (N0)? mem[696] : 1'b0;
//   assign r_data_o[156] = (N3)? mem[156] : 
//                          (N0)? mem[695] : 1'b0;
//   assign r_data_o[155] = (N3)? mem[155] : 
//                          (N0)? mem[694] : 1'b0;
//   assign r_data_o[154] = (N3)? mem[154] : 
//                          (N0)? mem[693] : 1'b0;
//   assign r_data_o[153] = (N3)? mem[153] : 
//                          (N0)? mem[692] : 1'b0;
//   assign r_data_o[152] = (N3)? mem[152] : 
//                          (N0)? mem[691] : 1'b0;
//   assign r_data_o[151] = (N3)? mem[151] : 
//                          (N0)? mem[690] : 1'b0;
//   assign r_data_o[150] = (N3)? mem[150] : 
//                          (N0)? mem[689] : 1'b0;
//   assign r_data_o[149] = (N3)? mem[149] : 
//                          (N0)? mem[688] : 1'b0;
//   assign r_data_o[148] = (N3)? mem[148] : 
//                          (N0)? mem[687] : 1'b0;
//   assign r_data_o[147] = (N3)? mem[147] : 
//                          (N0)? mem[686] : 1'b0;
//   assign r_data_o[146] = (N3)? mem[146] : 
//                          (N0)? mem[685] : 1'b0;
//   assign r_data_o[145] = (N3)? mem[145] : 
//                          (N0)? mem[684] : 1'b0;
//   assign r_data_o[144] = (N3)? mem[144] : 
//                          (N0)? mem[683] : 1'b0;
//   assign r_data_o[143] = (N3)? mem[143] : 
//                          (N0)? mem[682] : 1'b0;
//   assign r_data_o[142] = (N3)? mem[142] : 
//                          (N0)? mem[681] : 1'b0;
//   assign r_data_o[141] = (N3)? mem[141] : 
//                          (N0)? mem[680] : 1'b0;
//   assign r_data_o[140] = (N3)? mem[140] : 
//                          (N0)? mem[679] : 1'b0;
//   assign r_data_o[139] = (N3)? mem[139] : 
//                          (N0)? mem[678] : 1'b0;
//   assign r_data_o[138] = (N3)? mem[138] : 
//                          (N0)? mem[677] : 1'b0;
//   assign r_data_o[137] = (N3)? mem[137] : 
//                          (N0)? mem[676] : 1'b0;
//   assign r_data_o[136] = (N3)? mem[136] : 
//                          (N0)? mem[675] : 1'b0;
//   assign r_data_o[135] = (N3)? mem[135] : 
//                          (N0)? mem[674] : 1'b0;
//   assign r_data_o[134] = (N3)? mem[134] : 
//                          (N0)? mem[673] : 1'b0;
//   assign r_data_o[133] = (N3)? mem[133] : 
//                          (N0)? mem[672] : 1'b0;
//   assign r_data_o[132] = (N3)? mem[132] : 
//                          (N0)? mem[671] : 1'b0;
//   assign r_data_o[131] = (N3)? mem[131] : 
//                          (N0)? mem[670] : 1'b0;
//   assign r_data_o[130] = (N3)? mem[130] : 
//                          (N0)? mem[669] : 1'b0;
//   assign r_data_o[129] = (N3)? mem[129] : 
//                          (N0)? mem[668] : 1'b0;
//   assign r_data_o[128] = (N3)? mem[128] : 
//                          (N0)? mem[667] : 1'b0;
//   assign r_data_o[127] = (N3)? mem[127] : 
//                          (N0)? mem[666] : 1'b0;
//   assign r_data_o[126] = (N3)? mem[126] : 
//                          (N0)? mem[665] : 1'b0;
//   assign r_data_o[125] = (N3)? mem[125] : 
//                          (N0)? mem[664] : 1'b0;
//   assign r_data_o[124] = (N3)? mem[124] : 
//                          (N0)? mem[663] : 1'b0;
//   assign r_data_o[123] = (N3)? mem[123] : 
//                          (N0)? mem[662] : 1'b0;
//   assign r_data_o[122] = (N3)? mem[122] : 
//                          (N0)? mem[661] : 1'b0;
//   assign r_data_o[121] = (N3)? mem[121] : 
//                          (N0)? mem[660] : 1'b0;
//   assign r_data_o[120] = (N3)? mem[120] : 
//                          (N0)? mem[659] : 1'b0;
//   assign r_data_o[119] = (N3)? mem[119] : 
//                          (N0)? mem[658] : 1'b0;
//   assign r_data_o[118] = (N3)? mem[118] : 
//                          (N0)? mem[657] : 1'b0;
//   assign r_data_o[117] = (N3)? mem[117] : 
//                          (N0)? mem[656] : 1'b0;
//   assign r_data_o[116] = (N3)? mem[116] : 
//                          (N0)? mem[655] : 1'b0;
//   assign r_data_o[115] = (N3)? mem[115] : 
//                          (N0)? mem[654] : 1'b0;
//   assign r_data_o[114] = (N3)? mem[114] : 
//                          (N0)? mem[653] : 1'b0;
//   assign r_data_o[113] = (N3)? mem[113] : 
//                          (N0)? mem[652] : 1'b0;
//   assign r_data_o[112] = (N3)? mem[112] : 
//                          (N0)? mem[651] : 1'b0;
//   assign r_data_o[111] = (N3)? mem[111] : 
//                          (N0)? mem[650] : 1'b0;
//   assign r_data_o[110] = (N3)? mem[110] : 
//                          (N0)? mem[649] : 1'b0;
//   assign r_data_o[109] = (N3)? mem[109] : 
//                          (N0)? mem[648] : 1'b0;
//   assign r_data_o[108] = (N3)? mem[108] : 
//                          (N0)? mem[647] : 1'b0;
//   assign r_data_o[107] = (N3)? mem[107] : 
//                          (N0)? mem[646] : 1'b0;
//   assign r_data_o[106] = (N3)? mem[106] : 
//                          (N0)? mem[645] : 1'b0;
//   assign r_data_o[105] = (N3)? mem[105] : 
//                          (N0)? mem[644] : 1'b0;
//   assign r_data_o[104] = (N3)? mem[104] : 
//                          (N0)? mem[643] : 1'b0;
//   assign r_data_o[103] = (N3)? mem[103] : 
//                          (N0)? mem[642] : 1'b0;
//   assign r_data_o[102] = (N3)? mem[102] : 
//                          (N0)? mem[641] : 1'b0;
//   assign r_data_o[101] = (N3)? mem[101] : 
//                          (N0)? mem[640] : 1'b0;
//   assign r_data_o[100] = (N3)? mem[100] : 
//                          (N0)? mem[639] : 1'b0;
//   assign r_data_o[99] = (N3)? mem[99] : 
//                         (N0)? mem[638] : 1'b0;
//   assign r_data_o[98] = (N3)? mem[98] : 
//                         (N0)? mem[637] : 1'b0;
//   assign r_data_o[97] = (N3)? mem[97] : 
//                         (N0)? mem[636] : 1'b0;
//   assign r_data_o[96] = (N3)? mem[96] : 
//                         (N0)? mem[635] : 1'b0;
//   assign r_data_o[95] = (N3)? mem[95] : 
//                         (N0)? mem[634] : 1'b0;
//   assign r_data_o[94] = (N3)? mem[94] : 
//                         (N0)? mem[633] : 1'b0;
//   assign r_data_o[93] = (N3)? mem[93] : 
//                         (N0)? mem[632] : 1'b0;
//   assign r_data_o[92] = (N3)? mem[92] : 
//                         (N0)? mem[631] : 1'b0;
//   assign r_data_o[91] = (N3)? mem[91] : 
//                         (N0)? mem[630] : 1'b0;
//   assign r_data_o[90] = (N3)? mem[90] : 
//                         (N0)? mem[629] : 1'b0;
//   assign r_data_o[89] = (N3)? mem[89] : 
//                         (N0)? mem[628] : 1'b0;
//   assign r_data_o[88] = (N3)? mem[88] : 
//                         (N0)? mem[627] : 1'b0;
//   assign r_data_o[87] = (N3)? mem[87] : 
//                         (N0)? mem[626] : 1'b0;
//   assign r_data_o[86] = (N3)? mem[86] : 
//                         (N0)? mem[625] : 1'b0;
//   assign r_data_o[85] = (N3)? mem[85] : 
//                         (N0)? mem[624] : 1'b0;
//   assign r_data_o[84] = (N3)? mem[84] : 
//                         (N0)? mem[623] : 1'b0;
//   assign r_data_o[83] = (N3)? mem[83] : 
//                         (N0)? mem[622] : 1'b0;
//   assign r_data_o[82] = (N3)? mem[82] : 
//                         (N0)? mem[621] : 1'b0;
//   assign r_data_o[81] = (N3)? mem[81] : 
//                         (N0)? mem[620] : 1'b0;
//   assign r_data_o[80] = (N3)? mem[80] : 
//                         (N0)? mem[619] : 1'b0;
//   assign r_data_o[79] = (N3)? mem[79] : 
//                         (N0)? mem[618] : 1'b0;
//   assign r_data_o[78] = (N3)? mem[78] : 
//                         (N0)? mem[617] : 1'b0;
//   assign r_data_o[77] = (N3)? mem[77] : 
//                         (N0)? mem[616] : 1'b0;
//   assign r_data_o[76] = (N3)? mem[76] : 
//                         (N0)? mem[615] : 1'b0;
//   assign r_data_o[75] = (N3)? mem[75] : 
//                         (N0)? mem[614] : 1'b0;
//   assign r_data_o[74] = (N3)? mem[74] : 
//                         (N0)? mem[613] : 1'b0;
//   assign r_data_o[73] = (N3)? mem[73] : 
//                         (N0)? mem[612] : 1'b0;
//   assign r_data_o[72] = (N3)? mem[72] : 
//                         (N0)? mem[611] : 1'b0;
//   assign r_data_o[71] = (N3)? mem[71] : 
//                         (N0)? mem[610] : 1'b0;
//   assign r_data_o[70] = (N3)? mem[70] : 
//                         (N0)? mem[609] : 1'b0;
//   assign r_data_o[69] = (N3)? mem[69] : 
//                         (N0)? mem[608] : 1'b0;
//   assign r_data_o[68] = (N3)? mem[68] : 
//                         (N0)? mem[607] : 1'b0;
//   assign r_data_o[67] = (N3)? mem[67] : 
//                         (N0)? mem[606] : 1'b0;
//   assign r_data_o[66] = (N3)? mem[66] : 
//                         (N0)? mem[605] : 1'b0;
//   assign r_data_o[65] = (N3)? mem[65] : 
//                         (N0)? mem[604] : 1'b0;
//   assign r_data_o[64] = (N3)? mem[64] : 
//                         (N0)? mem[603] : 1'b0;
//   assign r_data_o[63] = (N3)? mem[63] : 
//                         (N0)? mem[602] : 1'b0;
//   assign r_data_o[62] = (N3)? mem[62] : 
//                         (N0)? mem[601] : 1'b0;
//   assign r_data_o[61] = (N3)? mem[61] : 
//                         (N0)? mem[600] : 1'b0;
//   assign r_data_o[60] = (N3)? mem[60] : 
//                         (N0)? mem[599] : 1'b0;
//   assign r_data_o[59] = (N3)? mem[59] : 
//                         (N0)? mem[598] : 1'b0;
//   assign r_data_o[58] = (N3)? mem[58] : 
//                         (N0)? mem[597] : 1'b0;
//   assign r_data_o[57] = (N3)? mem[57] : 
//                         (N0)? mem[596] : 1'b0;
//   assign r_data_o[56] = (N3)? mem[56] : 
//                         (N0)? mem[595] : 1'b0;
//   assign r_data_o[55] = (N3)? mem[55] : 
//                         (N0)? mem[594] : 1'b0;
//   assign r_data_o[54] = (N3)? mem[54] : 
//                         (N0)? mem[593] : 1'b0;
//   assign r_data_o[53] = (N3)? mem[53] : 
//                         (N0)? mem[592] : 1'b0;
//   assign r_data_o[52] = (N3)? mem[52] : 
//                         (N0)? mem[591] : 1'b0;
//   assign r_data_o[51] = (N3)? mem[51] : 
//                         (N0)? mem[590] : 1'b0;
//   assign r_data_o[50] = (N3)? mem[50] : 
//                         (N0)? mem[589] : 1'b0;
//   assign r_data_o[49] = (N3)? mem[49] : 
//                         (N0)? mem[588] : 1'b0;
//   assign r_data_o[48] = (N3)? mem[48] : 
//                         (N0)? mem[587] : 1'b0;
//   assign r_data_o[47] = (N3)? mem[47] : 
//                         (N0)? mem[586] : 1'b0;
//   assign r_data_o[46] = (N3)? mem[46] : 
//                         (N0)? mem[585] : 1'b0;
//   assign r_data_o[45] = (N3)? mem[45] : 
//                         (N0)? mem[584] : 1'b0;
//   assign r_data_o[44] = (N3)? mem[44] : 
//                         (N0)? mem[583] : 1'b0;
//   assign r_data_o[43] = (N3)? mem[43] : 
//                         (N0)? mem[582] : 1'b0;
//   assign r_data_o[42] = (N3)? mem[42] : 
//                         (N0)? mem[581] : 1'b0;
//   assign r_data_o[41] = (N3)? mem[41] : 
//                         (N0)? mem[580] : 1'b0;
//   assign r_data_o[40] = (N3)? mem[40] : 
//                         (N0)? mem[579] : 1'b0;
//   assign r_data_o[39] = (N3)? mem[39] : 
//                         (N0)? mem[578] : 1'b0;
//   assign r_data_o[38] = (N3)? mem[38] : 
//                         (N0)? mem[577] : 1'b0;
//   assign r_data_o[37] = (N3)? mem[37] : 
//                         (N0)? mem[576] : 1'b0;
//   assign r_data_o[36] = (N3)? mem[36] : 
//                         (N0)? mem[575] : 1'b0;
//   assign r_data_o[35] = (N3)? mem[35] : 
//                         (N0)? mem[574] : 1'b0;
//   assign r_data_o[34] = (N3)? mem[34] : 
//                         (N0)? mem[573] : 1'b0;
//   assign r_data_o[33] = (N3)? mem[33] : 
//                         (N0)? mem[572] : 1'b0;
//   assign r_data_o[32] = (N3)? mem[32] : 
//                         (N0)? mem[571] : 1'b0;
//   assign r_data_o[31] = (N3)? mem[31] : 
//                         (N0)? mem[570] : 1'b0;
//   assign r_data_o[30] = (N3)? mem[30] : 
//                         (N0)? mem[569] : 1'b0;
//   assign r_data_o[29] = (N3)? mem[29] : 
//                         (N0)? mem[568] : 1'b0;
//   assign r_data_o[28] = (N3)? mem[28] : 
//                         (N0)? mem[567] : 1'b0;
//   assign r_data_o[27] = (N3)? mem[27] : 
//                         (N0)? mem[566] : 1'b0;
//   assign r_data_o[26] = (N3)? mem[26] : 
//                         (N0)? mem[565] : 1'b0;
//   assign r_data_o[25] = (N3)? mem[25] : 
//                         (N0)? mem[564] : 1'b0;
//   assign r_data_o[24] = (N3)? mem[24] : 
//                         (N0)? mem[563] : 1'b0;
//   assign r_data_o[23] = (N3)? mem[23] : 
//                         (N0)? mem[562] : 1'b0;
//   assign r_data_o[22] = (N3)? mem[22] : 
//                         (N0)? mem[561] : 1'b0;
//   assign r_data_o[21] = (N3)? mem[21] : 
//                         (N0)? mem[560] : 1'b0;
//   assign r_data_o[20] = (N3)? mem[20] : 
//                         (N0)? mem[559] : 1'b0;
//   assign r_data_o[19] = (N3)? mem[19] : 
//                         (N0)? mem[558] : 1'b0;
//   assign r_data_o[18] = (N3)? mem[18] : 
//                         (N0)? mem[557] : 1'b0;
//   assign r_data_o[17] = (N3)? mem[17] : 
//                         (N0)? mem[556] : 1'b0;
//   assign r_data_o[16] = (N3)? mem[16] : 
//                         (N0)? mem[555] : 1'b0;
//   assign r_data_o[15] = (N3)? mem[15] : 
//                         (N0)? mem[554] : 1'b0;
//   assign r_data_o[14] = (N3)? mem[14] : 
//                         (N0)? mem[553] : 1'b0;
//   assign r_data_o[13] = (N3)? mem[13] : 
//                         (N0)? mem[552] : 1'b0;
//   assign r_data_o[12] = (N3)? mem[12] : 
//                         (N0)? mem[551] : 1'b0;
//   assign r_data_o[11] = (N3)? mem[11] : 
//                         (N0)? mem[550] : 1'b0;
//   assign r_data_o[10] = (N3)? mem[10] : 
//                         (N0)? mem[549] : 1'b0;
//   assign r_data_o[9] = (N3)? mem[9] : 
//                        (N0)? mem[548] : 1'b0;
//   assign r_data_o[8] = (N3)? mem[8] : 
//                        (N0)? mem[547] : 1'b0;
//   assign r_data_o[7] = (N3)? mem[7] : 
//                        (N0)? mem[546] : 1'b0;
//   assign r_data_o[6] = (N3)? mem[6] : 
//                        (N0)? mem[545] : 1'b0;
//   assign r_data_o[5] = (N3)? mem[5] : 
//                        (N0)? mem[544] : 1'b0;
//   assign r_data_o[4] = (N3)? mem[4] : 
//                        (N0)? mem[543] : 1'b0;
//   assign r_data_o[3] = (N3)? mem[3] : 
//                        (N0)? mem[542] : 1'b0;
//   assign r_data_o[2] = (N3)? mem[2] : 
//                        (N0)? mem[541] : 1'b0;
//   assign r_data_o[1] = (N3)? mem[1] : 
//                        (N0)? mem[540] : 1'b0;
//   assign r_data_o[0] = (N3)? mem[0] : 
//                        (N0)? mem[539] : 1'b0;
//   assign N5 = ~w_addr_i[0];
//   assign { N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], N5, N5, N5, N5, N5, N5 } : 
//                                                                        (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
//   assign N1 = w_v_i;
//   assign N2 = N4;
//   assign N3 = ~r_addr_i[0];
//   assign N4 = ~w_v_i;

//   always @(posedge w_clk_i) begin
//     if(N13) begin
//       { mem[1077:979], mem[539:539] } <= { w_data_i[538:440], w_data_i[0:0] };
//     end 
//     if(N14) begin
//       { mem[978:880], mem[540:540] } <= { w_data_i[439:341], w_data_i[1:1] };
//     end 
//     if(N15) begin
//       { mem[879:781], mem[541:541] } <= { w_data_i[340:242], w_data_i[2:2] };
//     end 
//     if(N16) begin
//       { mem[780:682], mem[542:542] } <= { w_data_i[241:143], w_data_i[3:3] };
//     end 
//     if(N17) begin
//       { mem[681:583], mem[543:543] } <= { w_data_i[142:44], w_data_i[4:4] };
//     end 
//     if(N18) begin
//       { mem[582:544] } <= { w_data_i[43:5] };
//     end 
//     if(N7) begin
//       { mem[538:440], mem[0:0] } <= { w_data_i[538:440], w_data_i[0:0] };
//     end 
//     if(N8) begin
//       { mem[439:341], mem[1:1] } <= { w_data_i[439:341], w_data_i[1:1] };
//     end 
//     if(N9) begin
//       { mem[340:242], mem[2:2] } <= { w_data_i[340:242], w_data_i[2:2] };
//     end 
//     if(N10) begin
//       { mem[241:143], mem[3:3] } <= { w_data_i[241:143], w_data_i[3:3] };
//     end 
//     if(N11) begin
//       { mem[142:44], mem[4:4] } <= { w_data_i[142:44], w_data_i[4:4] };
//     end 
//     if(N12) begin
//       { mem[43:5] } <= { w_data_i[43:5] };
//     end 
//   end


// endmodule



module bsg_mem_1r1w_width_p539_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [538:0] w_data_i;
  input [0:0] r_addr_i;
  output [538:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [538:0] r_data_o;

  bsg_mem_p539
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p539
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [538:0] data_i;
  output [538:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [538:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p539_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 : 
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 : 
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 : 
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 : 
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 : 
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 : 
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end 
    if(N9) begin
      tail_r <= N10;
    end 
    if(N11) begin
      head_r <= N12;
    end 
  end


endmodule



module bp_fe_lce_tr_resp_in_data_width_p64_lce_data_width_p512_lce_addr_width_p22_lce_sets_p64_ways_p8_num_cce_p1_num_lce_p2_block_size_in_bytes_p8
(
  tr_received_o,
  lce_tr_resp_i,
  lce_tr_resp_v_i,
  lce_tr_resp_yumi_o,
  data_mem_pkt_v_o,
  data_mem_pkt_o,
  data_mem_pkt_yumi_i
);

  input [538:0] lce_tr_resp_i;
  output [521:0] data_mem_pkt_o;
  input lce_tr_resp_v_i;
  input data_mem_pkt_yumi_i;
  output tr_received_o;
  output lce_tr_resp_yumi_o;
  output data_mem_pkt_v_o;
  wire [521:0] data_mem_pkt_o;
  wire tr_received_o,lce_tr_resp_yumi_o,data_mem_pkt_v_o,lce_tr_resp_v_i;
  assign data_mem_pkt_o[512] = 1'b1;
  assign data_mem_pkt_v_o = lce_tr_resp_v_i;
  assign data_mem_pkt_o[521] = lce_tr_resp_i[523];
  assign data_mem_pkt_o[520] = lce_tr_resp_i[522];
  assign data_mem_pkt_o[519] = lce_tr_resp_i[521];
  assign data_mem_pkt_o[518] = lce_tr_resp_i[520];
  assign data_mem_pkt_o[517] = lce_tr_resp_i[519];
  assign data_mem_pkt_o[516] = lce_tr_resp_i[518];
  assign data_mem_pkt_o[515] = lce_tr_resp_i[536];
  assign data_mem_pkt_o[514] = lce_tr_resp_i[535];
  assign data_mem_pkt_o[513] = lce_tr_resp_i[534];
  assign data_mem_pkt_o[511] = lce_tr_resp_i[511];
  assign data_mem_pkt_o[510] = lce_tr_resp_i[510];
  assign data_mem_pkt_o[509] = lce_tr_resp_i[509];
  assign data_mem_pkt_o[508] = lce_tr_resp_i[508];
  assign data_mem_pkt_o[507] = lce_tr_resp_i[507];
  assign data_mem_pkt_o[506] = lce_tr_resp_i[506];
  assign data_mem_pkt_o[505] = lce_tr_resp_i[505];
  assign data_mem_pkt_o[504] = lce_tr_resp_i[504];
  assign data_mem_pkt_o[503] = lce_tr_resp_i[503];
  assign data_mem_pkt_o[502] = lce_tr_resp_i[502];
  assign data_mem_pkt_o[501] = lce_tr_resp_i[501];
  assign data_mem_pkt_o[500] = lce_tr_resp_i[500];
  assign data_mem_pkt_o[499] = lce_tr_resp_i[499];
  assign data_mem_pkt_o[498] = lce_tr_resp_i[498];
  assign data_mem_pkt_o[497] = lce_tr_resp_i[497];
  assign data_mem_pkt_o[496] = lce_tr_resp_i[496];
  assign data_mem_pkt_o[495] = lce_tr_resp_i[495];
  assign data_mem_pkt_o[494] = lce_tr_resp_i[494];
  assign data_mem_pkt_o[493] = lce_tr_resp_i[493];
  assign data_mem_pkt_o[492] = lce_tr_resp_i[492];
  assign data_mem_pkt_o[491] = lce_tr_resp_i[491];
  assign data_mem_pkt_o[490] = lce_tr_resp_i[490];
  assign data_mem_pkt_o[489] = lce_tr_resp_i[489];
  assign data_mem_pkt_o[488] = lce_tr_resp_i[488];
  assign data_mem_pkt_o[487] = lce_tr_resp_i[487];
  assign data_mem_pkt_o[486] = lce_tr_resp_i[486];
  assign data_mem_pkt_o[485] = lce_tr_resp_i[485];
  assign data_mem_pkt_o[484] = lce_tr_resp_i[484];
  assign data_mem_pkt_o[483] = lce_tr_resp_i[483];
  assign data_mem_pkt_o[482] = lce_tr_resp_i[482];
  assign data_mem_pkt_o[481] = lce_tr_resp_i[481];
  assign data_mem_pkt_o[480] = lce_tr_resp_i[480];
  assign data_mem_pkt_o[479] = lce_tr_resp_i[479];
  assign data_mem_pkt_o[478] = lce_tr_resp_i[478];
  assign data_mem_pkt_o[477] = lce_tr_resp_i[477];
  assign data_mem_pkt_o[476] = lce_tr_resp_i[476];
  assign data_mem_pkt_o[475] = lce_tr_resp_i[475];
  assign data_mem_pkt_o[474] = lce_tr_resp_i[474];
  assign data_mem_pkt_o[473] = lce_tr_resp_i[473];
  assign data_mem_pkt_o[472] = lce_tr_resp_i[472];
  assign data_mem_pkt_o[471] = lce_tr_resp_i[471];
  assign data_mem_pkt_o[470] = lce_tr_resp_i[470];
  assign data_mem_pkt_o[469] = lce_tr_resp_i[469];
  assign data_mem_pkt_o[468] = lce_tr_resp_i[468];
  assign data_mem_pkt_o[467] = lce_tr_resp_i[467];
  assign data_mem_pkt_o[466] = lce_tr_resp_i[466];
  assign data_mem_pkt_o[465] = lce_tr_resp_i[465];
  assign data_mem_pkt_o[464] = lce_tr_resp_i[464];
  assign data_mem_pkt_o[463] = lce_tr_resp_i[463];
  assign data_mem_pkt_o[462] = lce_tr_resp_i[462];
  assign data_mem_pkt_o[461] = lce_tr_resp_i[461];
  assign data_mem_pkt_o[460] = lce_tr_resp_i[460];
  assign data_mem_pkt_o[459] = lce_tr_resp_i[459];
  assign data_mem_pkt_o[458] = lce_tr_resp_i[458];
  assign data_mem_pkt_o[457] = lce_tr_resp_i[457];
  assign data_mem_pkt_o[456] = lce_tr_resp_i[456];
  assign data_mem_pkt_o[455] = lce_tr_resp_i[455];
  assign data_mem_pkt_o[454] = lce_tr_resp_i[454];
  assign data_mem_pkt_o[453] = lce_tr_resp_i[453];
  assign data_mem_pkt_o[452] = lce_tr_resp_i[452];
  assign data_mem_pkt_o[451] = lce_tr_resp_i[451];
  assign data_mem_pkt_o[450] = lce_tr_resp_i[450];
  assign data_mem_pkt_o[449] = lce_tr_resp_i[449];
  assign data_mem_pkt_o[448] = lce_tr_resp_i[448];
  assign data_mem_pkt_o[447] = lce_tr_resp_i[447];
  assign data_mem_pkt_o[446] = lce_tr_resp_i[446];
  assign data_mem_pkt_o[445] = lce_tr_resp_i[445];
  assign data_mem_pkt_o[444] = lce_tr_resp_i[444];
  assign data_mem_pkt_o[443] = lce_tr_resp_i[443];
  assign data_mem_pkt_o[442] = lce_tr_resp_i[442];
  assign data_mem_pkt_o[441] = lce_tr_resp_i[441];
  assign data_mem_pkt_o[440] = lce_tr_resp_i[440];
  assign data_mem_pkt_o[439] = lce_tr_resp_i[439];
  assign data_mem_pkt_o[438] = lce_tr_resp_i[438];
  assign data_mem_pkt_o[437] = lce_tr_resp_i[437];
  assign data_mem_pkt_o[436] = lce_tr_resp_i[436];
  assign data_mem_pkt_o[435] = lce_tr_resp_i[435];
  assign data_mem_pkt_o[434] = lce_tr_resp_i[434];
  assign data_mem_pkt_o[433] = lce_tr_resp_i[433];
  assign data_mem_pkt_o[432] = lce_tr_resp_i[432];
  assign data_mem_pkt_o[431] = lce_tr_resp_i[431];
  assign data_mem_pkt_o[430] = lce_tr_resp_i[430];
  assign data_mem_pkt_o[429] = lce_tr_resp_i[429];
  assign data_mem_pkt_o[428] = lce_tr_resp_i[428];
  assign data_mem_pkt_o[427] = lce_tr_resp_i[427];
  assign data_mem_pkt_o[426] = lce_tr_resp_i[426];
  assign data_mem_pkt_o[425] = lce_tr_resp_i[425];
  assign data_mem_pkt_o[424] = lce_tr_resp_i[424];
  assign data_mem_pkt_o[423] = lce_tr_resp_i[423];
  assign data_mem_pkt_o[422] = lce_tr_resp_i[422];
  assign data_mem_pkt_o[421] = lce_tr_resp_i[421];
  assign data_mem_pkt_o[420] = lce_tr_resp_i[420];
  assign data_mem_pkt_o[419] = lce_tr_resp_i[419];
  assign data_mem_pkt_o[418] = lce_tr_resp_i[418];
  assign data_mem_pkt_o[417] = lce_tr_resp_i[417];
  assign data_mem_pkt_o[416] = lce_tr_resp_i[416];
  assign data_mem_pkt_o[415] = lce_tr_resp_i[415];
  assign data_mem_pkt_o[414] = lce_tr_resp_i[414];
  assign data_mem_pkt_o[413] = lce_tr_resp_i[413];
  assign data_mem_pkt_o[412] = lce_tr_resp_i[412];
  assign data_mem_pkt_o[411] = lce_tr_resp_i[411];
  assign data_mem_pkt_o[410] = lce_tr_resp_i[410];
  assign data_mem_pkt_o[409] = lce_tr_resp_i[409];
  assign data_mem_pkt_o[408] = lce_tr_resp_i[408];
  assign data_mem_pkt_o[407] = lce_tr_resp_i[407];
  assign data_mem_pkt_o[406] = lce_tr_resp_i[406];
  assign data_mem_pkt_o[405] = lce_tr_resp_i[405];
  assign data_mem_pkt_o[404] = lce_tr_resp_i[404];
  assign data_mem_pkt_o[403] = lce_tr_resp_i[403];
  assign data_mem_pkt_o[402] = lce_tr_resp_i[402];
  assign data_mem_pkt_o[401] = lce_tr_resp_i[401];
  assign data_mem_pkt_o[400] = lce_tr_resp_i[400];
  assign data_mem_pkt_o[399] = lce_tr_resp_i[399];
  assign data_mem_pkt_o[398] = lce_tr_resp_i[398];
  assign data_mem_pkt_o[397] = lce_tr_resp_i[397];
  assign data_mem_pkt_o[396] = lce_tr_resp_i[396];
  assign data_mem_pkt_o[395] = lce_tr_resp_i[395];
  assign data_mem_pkt_o[394] = lce_tr_resp_i[394];
  assign data_mem_pkt_o[393] = lce_tr_resp_i[393];
  assign data_mem_pkt_o[392] = lce_tr_resp_i[392];
  assign data_mem_pkt_o[391] = lce_tr_resp_i[391];
  assign data_mem_pkt_o[390] = lce_tr_resp_i[390];
  assign data_mem_pkt_o[389] = lce_tr_resp_i[389];
  assign data_mem_pkt_o[388] = lce_tr_resp_i[388];
  assign data_mem_pkt_o[387] = lce_tr_resp_i[387];
  assign data_mem_pkt_o[386] = lce_tr_resp_i[386];
  assign data_mem_pkt_o[385] = lce_tr_resp_i[385];
  assign data_mem_pkt_o[384] = lce_tr_resp_i[384];
  assign data_mem_pkt_o[383] = lce_tr_resp_i[383];
  assign data_mem_pkt_o[382] = lce_tr_resp_i[382];
  assign data_mem_pkt_o[381] = lce_tr_resp_i[381];
  assign data_mem_pkt_o[380] = lce_tr_resp_i[380];
  assign data_mem_pkt_o[379] = lce_tr_resp_i[379];
  assign data_mem_pkt_o[378] = lce_tr_resp_i[378];
  assign data_mem_pkt_o[377] = lce_tr_resp_i[377];
  assign data_mem_pkt_o[376] = lce_tr_resp_i[376];
  assign data_mem_pkt_o[375] = lce_tr_resp_i[375];
  assign data_mem_pkt_o[374] = lce_tr_resp_i[374];
  assign data_mem_pkt_o[373] = lce_tr_resp_i[373];
  assign data_mem_pkt_o[372] = lce_tr_resp_i[372];
  assign data_mem_pkt_o[371] = lce_tr_resp_i[371];
  assign data_mem_pkt_o[370] = lce_tr_resp_i[370];
  assign data_mem_pkt_o[369] = lce_tr_resp_i[369];
  assign data_mem_pkt_o[368] = lce_tr_resp_i[368];
  assign data_mem_pkt_o[367] = lce_tr_resp_i[367];
  assign data_mem_pkt_o[366] = lce_tr_resp_i[366];
  assign data_mem_pkt_o[365] = lce_tr_resp_i[365];
  assign data_mem_pkt_o[364] = lce_tr_resp_i[364];
  assign data_mem_pkt_o[363] = lce_tr_resp_i[363];
  assign data_mem_pkt_o[362] = lce_tr_resp_i[362];
  assign data_mem_pkt_o[361] = lce_tr_resp_i[361];
  assign data_mem_pkt_o[360] = lce_tr_resp_i[360];
  assign data_mem_pkt_o[359] = lce_tr_resp_i[359];
  assign data_mem_pkt_o[358] = lce_tr_resp_i[358];
  assign data_mem_pkt_o[357] = lce_tr_resp_i[357];
  assign data_mem_pkt_o[356] = lce_tr_resp_i[356];
  assign data_mem_pkt_o[355] = lce_tr_resp_i[355];
  assign data_mem_pkt_o[354] = lce_tr_resp_i[354];
  assign data_mem_pkt_o[353] = lce_tr_resp_i[353];
  assign data_mem_pkt_o[352] = lce_tr_resp_i[352];
  assign data_mem_pkt_o[351] = lce_tr_resp_i[351];
  assign data_mem_pkt_o[350] = lce_tr_resp_i[350];
  assign data_mem_pkt_o[349] = lce_tr_resp_i[349];
  assign data_mem_pkt_o[348] = lce_tr_resp_i[348];
  assign data_mem_pkt_o[347] = lce_tr_resp_i[347];
  assign data_mem_pkt_o[346] = lce_tr_resp_i[346];
  assign data_mem_pkt_o[345] = lce_tr_resp_i[345];
  assign data_mem_pkt_o[344] = lce_tr_resp_i[344];
  assign data_mem_pkt_o[343] = lce_tr_resp_i[343];
  assign data_mem_pkt_o[342] = lce_tr_resp_i[342];
  assign data_mem_pkt_o[341] = lce_tr_resp_i[341];
  assign data_mem_pkt_o[340] = lce_tr_resp_i[340];
  assign data_mem_pkt_o[339] = lce_tr_resp_i[339];
  assign data_mem_pkt_o[338] = lce_tr_resp_i[338];
  assign data_mem_pkt_o[337] = lce_tr_resp_i[337];
  assign data_mem_pkt_o[336] = lce_tr_resp_i[336];
  assign data_mem_pkt_o[335] = lce_tr_resp_i[335];
  assign data_mem_pkt_o[334] = lce_tr_resp_i[334];
  assign data_mem_pkt_o[333] = lce_tr_resp_i[333];
  assign data_mem_pkt_o[332] = lce_tr_resp_i[332];
  assign data_mem_pkt_o[331] = lce_tr_resp_i[331];
  assign data_mem_pkt_o[330] = lce_tr_resp_i[330];
  assign data_mem_pkt_o[329] = lce_tr_resp_i[329];
  assign data_mem_pkt_o[328] = lce_tr_resp_i[328];
  assign data_mem_pkt_o[327] = lce_tr_resp_i[327];
  assign data_mem_pkt_o[326] = lce_tr_resp_i[326];
  assign data_mem_pkt_o[325] = lce_tr_resp_i[325];
  assign data_mem_pkt_o[324] = lce_tr_resp_i[324];
  assign data_mem_pkt_o[323] = lce_tr_resp_i[323];
  assign data_mem_pkt_o[322] = lce_tr_resp_i[322];
  assign data_mem_pkt_o[321] = lce_tr_resp_i[321];
  assign data_mem_pkt_o[320] = lce_tr_resp_i[320];
  assign data_mem_pkt_o[319] = lce_tr_resp_i[319];
  assign data_mem_pkt_o[318] = lce_tr_resp_i[318];
  assign data_mem_pkt_o[317] = lce_tr_resp_i[317];
  assign data_mem_pkt_o[316] = lce_tr_resp_i[316];
  assign data_mem_pkt_o[315] = lce_tr_resp_i[315];
  assign data_mem_pkt_o[314] = lce_tr_resp_i[314];
  assign data_mem_pkt_o[313] = lce_tr_resp_i[313];
  assign data_mem_pkt_o[312] = lce_tr_resp_i[312];
  assign data_mem_pkt_o[311] = lce_tr_resp_i[311];
  assign data_mem_pkt_o[310] = lce_tr_resp_i[310];
  assign data_mem_pkt_o[309] = lce_tr_resp_i[309];
  assign data_mem_pkt_o[308] = lce_tr_resp_i[308];
  assign data_mem_pkt_o[307] = lce_tr_resp_i[307];
  assign data_mem_pkt_o[306] = lce_tr_resp_i[306];
  assign data_mem_pkt_o[305] = lce_tr_resp_i[305];
  assign data_mem_pkt_o[304] = lce_tr_resp_i[304];
  assign data_mem_pkt_o[303] = lce_tr_resp_i[303];
  assign data_mem_pkt_o[302] = lce_tr_resp_i[302];
  assign data_mem_pkt_o[301] = lce_tr_resp_i[301];
  assign data_mem_pkt_o[300] = lce_tr_resp_i[300];
  assign data_mem_pkt_o[299] = lce_tr_resp_i[299];
  assign data_mem_pkt_o[298] = lce_tr_resp_i[298];
  assign data_mem_pkt_o[297] = lce_tr_resp_i[297];
  assign data_mem_pkt_o[296] = lce_tr_resp_i[296];
  assign data_mem_pkt_o[295] = lce_tr_resp_i[295];
  assign data_mem_pkt_o[294] = lce_tr_resp_i[294];
  assign data_mem_pkt_o[293] = lce_tr_resp_i[293];
  assign data_mem_pkt_o[292] = lce_tr_resp_i[292];
  assign data_mem_pkt_o[291] = lce_tr_resp_i[291];
  assign data_mem_pkt_o[290] = lce_tr_resp_i[290];
  assign data_mem_pkt_o[289] = lce_tr_resp_i[289];
  assign data_mem_pkt_o[288] = lce_tr_resp_i[288];
  assign data_mem_pkt_o[287] = lce_tr_resp_i[287];
  assign data_mem_pkt_o[286] = lce_tr_resp_i[286];
  assign data_mem_pkt_o[285] = lce_tr_resp_i[285];
  assign data_mem_pkt_o[284] = lce_tr_resp_i[284];
  assign data_mem_pkt_o[283] = lce_tr_resp_i[283];
  assign data_mem_pkt_o[282] = lce_tr_resp_i[282];
  assign data_mem_pkt_o[281] = lce_tr_resp_i[281];
  assign data_mem_pkt_o[280] = lce_tr_resp_i[280];
  assign data_mem_pkt_o[279] = lce_tr_resp_i[279];
  assign data_mem_pkt_o[278] = lce_tr_resp_i[278];
  assign data_mem_pkt_o[277] = lce_tr_resp_i[277];
  assign data_mem_pkt_o[276] = lce_tr_resp_i[276];
  assign data_mem_pkt_o[275] = lce_tr_resp_i[275];
  assign data_mem_pkt_o[274] = lce_tr_resp_i[274];
  assign data_mem_pkt_o[273] = lce_tr_resp_i[273];
  assign data_mem_pkt_o[272] = lce_tr_resp_i[272];
  assign data_mem_pkt_o[271] = lce_tr_resp_i[271];
  assign data_mem_pkt_o[270] = lce_tr_resp_i[270];
  assign data_mem_pkt_o[269] = lce_tr_resp_i[269];
  assign data_mem_pkt_o[268] = lce_tr_resp_i[268];
  assign data_mem_pkt_o[267] = lce_tr_resp_i[267];
  assign data_mem_pkt_o[266] = lce_tr_resp_i[266];
  assign data_mem_pkt_o[265] = lce_tr_resp_i[265];
  assign data_mem_pkt_o[264] = lce_tr_resp_i[264];
  assign data_mem_pkt_o[263] = lce_tr_resp_i[263];
  assign data_mem_pkt_o[262] = lce_tr_resp_i[262];
  assign data_mem_pkt_o[261] = lce_tr_resp_i[261];
  assign data_mem_pkt_o[260] = lce_tr_resp_i[260];
  assign data_mem_pkt_o[259] = lce_tr_resp_i[259];
  assign data_mem_pkt_o[258] = lce_tr_resp_i[258];
  assign data_mem_pkt_o[257] = lce_tr_resp_i[257];
  assign data_mem_pkt_o[256] = lce_tr_resp_i[256];
  assign data_mem_pkt_o[255] = lce_tr_resp_i[255];
  assign data_mem_pkt_o[254] = lce_tr_resp_i[254];
  assign data_mem_pkt_o[253] = lce_tr_resp_i[253];
  assign data_mem_pkt_o[252] = lce_tr_resp_i[252];
  assign data_mem_pkt_o[251] = lce_tr_resp_i[251];
  assign data_mem_pkt_o[250] = lce_tr_resp_i[250];
  assign data_mem_pkt_o[249] = lce_tr_resp_i[249];
  assign data_mem_pkt_o[248] = lce_tr_resp_i[248];
  assign data_mem_pkt_o[247] = lce_tr_resp_i[247];
  assign data_mem_pkt_o[246] = lce_tr_resp_i[246];
  assign data_mem_pkt_o[245] = lce_tr_resp_i[245];
  assign data_mem_pkt_o[244] = lce_tr_resp_i[244];
  assign data_mem_pkt_o[243] = lce_tr_resp_i[243];
  assign data_mem_pkt_o[242] = lce_tr_resp_i[242];
  assign data_mem_pkt_o[241] = lce_tr_resp_i[241];
  assign data_mem_pkt_o[240] = lce_tr_resp_i[240];
  assign data_mem_pkt_o[239] = lce_tr_resp_i[239];
  assign data_mem_pkt_o[238] = lce_tr_resp_i[238];
  assign data_mem_pkt_o[237] = lce_tr_resp_i[237];
  assign data_mem_pkt_o[236] = lce_tr_resp_i[236];
  assign data_mem_pkt_o[235] = lce_tr_resp_i[235];
  assign data_mem_pkt_o[234] = lce_tr_resp_i[234];
  assign data_mem_pkt_o[233] = lce_tr_resp_i[233];
  assign data_mem_pkt_o[232] = lce_tr_resp_i[232];
  assign data_mem_pkt_o[231] = lce_tr_resp_i[231];
  assign data_mem_pkt_o[230] = lce_tr_resp_i[230];
  assign data_mem_pkt_o[229] = lce_tr_resp_i[229];
  assign data_mem_pkt_o[228] = lce_tr_resp_i[228];
  assign data_mem_pkt_o[227] = lce_tr_resp_i[227];
  assign data_mem_pkt_o[226] = lce_tr_resp_i[226];
  assign data_mem_pkt_o[225] = lce_tr_resp_i[225];
  assign data_mem_pkt_o[224] = lce_tr_resp_i[224];
  assign data_mem_pkt_o[223] = lce_tr_resp_i[223];
  assign data_mem_pkt_o[222] = lce_tr_resp_i[222];
  assign data_mem_pkt_o[221] = lce_tr_resp_i[221];
  assign data_mem_pkt_o[220] = lce_tr_resp_i[220];
  assign data_mem_pkt_o[219] = lce_tr_resp_i[219];
  assign data_mem_pkt_o[218] = lce_tr_resp_i[218];
  assign data_mem_pkt_o[217] = lce_tr_resp_i[217];
  assign data_mem_pkt_o[216] = lce_tr_resp_i[216];
  assign data_mem_pkt_o[215] = lce_tr_resp_i[215];
  assign data_mem_pkt_o[214] = lce_tr_resp_i[214];
  assign data_mem_pkt_o[213] = lce_tr_resp_i[213];
  assign data_mem_pkt_o[212] = lce_tr_resp_i[212];
  assign data_mem_pkt_o[211] = lce_tr_resp_i[211];
  assign data_mem_pkt_o[210] = lce_tr_resp_i[210];
  assign data_mem_pkt_o[209] = lce_tr_resp_i[209];
  assign data_mem_pkt_o[208] = lce_tr_resp_i[208];
  assign data_mem_pkt_o[207] = lce_tr_resp_i[207];
  assign data_mem_pkt_o[206] = lce_tr_resp_i[206];
  assign data_mem_pkt_o[205] = lce_tr_resp_i[205];
  assign data_mem_pkt_o[204] = lce_tr_resp_i[204];
  assign data_mem_pkt_o[203] = lce_tr_resp_i[203];
  assign data_mem_pkt_o[202] = lce_tr_resp_i[202];
  assign data_mem_pkt_o[201] = lce_tr_resp_i[201];
  assign data_mem_pkt_o[200] = lce_tr_resp_i[200];
  assign data_mem_pkt_o[199] = lce_tr_resp_i[199];
  assign data_mem_pkt_o[198] = lce_tr_resp_i[198];
  assign data_mem_pkt_o[197] = lce_tr_resp_i[197];
  assign data_mem_pkt_o[196] = lce_tr_resp_i[196];
  assign data_mem_pkt_o[195] = lce_tr_resp_i[195];
  assign data_mem_pkt_o[194] = lce_tr_resp_i[194];
  assign data_mem_pkt_o[193] = lce_tr_resp_i[193];
  assign data_mem_pkt_o[192] = lce_tr_resp_i[192];
  assign data_mem_pkt_o[191] = lce_tr_resp_i[191];
  assign data_mem_pkt_o[190] = lce_tr_resp_i[190];
  assign data_mem_pkt_o[189] = lce_tr_resp_i[189];
  assign data_mem_pkt_o[188] = lce_tr_resp_i[188];
  assign data_mem_pkt_o[187] = lce_tr_resp_i[187];
  assign data_mem_pkt_o[186] = lce_tr_resp_i[186];
  assign data_mem_pkt_o[185] = lce_tr_resp_i[185];
  assign data_mem_pkt_o[184] = lce_tr_resp_i[184];
  assign data_mem_pkt_o[183] = lce_tr_resp_i[183];
  assign data_mem_pkt_o[182] = lce_tr_resp_i[182];
  assign data_mem_pkt_o[181] = lce_tr_resp_i[181];
  assign data_mem_pkt_o[180] = lce_tr_resp_i[180];
  assign data_mem_pkt_o[179] = lce_tr_resp_i[179];
  assign data_mem_pkt_o[178] = lce_tr_resp_i[178];
  assign data_mem_pkt_o[177] = lce_tr_resp_i[177];
  assign data_mem_pkt_o[176] = lce_tr_resp_i[176];
  assign data_mem_pkt_o[175] = lce_tr_resp_i[175];
  assign data_mem_pkt_o[174] = lce_tr_resp_i[174];
  assign data_mem_pkt_o[173] = lce_tr_resp_i[173];
  assign data_mem_pkt_o[172] = lce_tr_resp_i[172];
  assign data_mem_pkt_o[171] = lce_tr_resp_i[171];
  assign data_mem_pkt_o[170] = lce_tr_resp_i[170];
  assign data_mem_pkt_o[169] = lce_tr_resp_i[169];
  assign data_mem_pkt_o[168] = lce_tr_resp_i[168];
  assign data_mem_pkt_o[167] = lce_tr_resp_i[167];
  assign data_mem_pkt_o[166] = lce_tr_resp_i[166];
  assign data_mem_pkt_o[165] = lce_tr_resp_i[165];
  assign data_mem_pkt_o[164] = lce_tr_resp_i[164];
  assign data_mem_pkt_o[163] = lce_tr_resp_i[163];
  assign data_mem_pkt_o[162] = lce_tr_resp_i[162];
  assign data_mem_pkt_o[161] = lce_tr_resp_i[161];
  assign data_mem_pkt_o[160] = lce_tr_resp_i[160];
  assign data_mem_pkt_o[159] = lce_tr_resp_i[159];
  assign data_mem_pkt_o[158] = lce_tr_resp_i[158];
  assign data_mem_pkt_o[157] = lce_tr_resp_i[157];
  assign data_mem_pkt_o[156] = lce_tr_resp_i[156];
  assign data_mem_pkt_o[155] = lce_tr_resp_i[155];
  assign data_mem_pkt_o[154] = lce_tr_resp_i[154];
  assign data_mem_pkt_o[153] = lce_tr_resp_i[153];
  assign data_mem_pkt_o[152] = lce_tr_resp_i[152];
  assign data_mem_pkt_o[151] = lce_tr_resp_i[151];
  assign data_mem_pkt_o[150] = lce_tr_resp_i[150];
  assign data_mem_pkt_o[149] = lce_tr_resp_i[149];
  assign data_mem_pkt_o[148] = lce_tr_resp_i[148];
  assign data_mem_pkt_o[147] = lce_tr_resp_i[147];
  assign data_mem_pkt_o[146] = lce_tr_resp_i[146];
  assign data_mem_pkt_o[145] = lce_tr_resp_i[145];
  assign data_mem_pkt_o[144] = lce_tr_resp_i[144];
  assign data_mem_pkt_o[143] = lce_tr_resp_i[143];
  assign data_mem_pkt_o[142] = lce_tr_resp_i[142];
  assign data_mem_pkt_o[141] = lce_tr_resp_i[141];
  assign data_mem_pkt_o[140] = lce_tr_resp_i[140];
  assign data_mem_pkt_o[139] = lce_tr_resp_i[139];
  assign data_mem_pkt_o[138] = lce_tr_resp_i[138];
  assign data_mem_pkt_o[137] = lce_tr_resp_i[137];
  assign data_mem_pkt_o[136] = lce_tr_resp_i[136];
  assign data_mem_pkt_o[135] = lce_tr_resp_i[135];
  assign data_mem_pkt_o[134] = lce_tr_resp_i[134];
  assign data_mem_pkt_o[133] = lce_tr_resp_i[133];
  assign data_mem_pkt_o[132] = lce_tr_resp_i[132];
  assign data_mem_pkt_o[131] = lce_tr_resp_i[131];
  assign data_mem_pkt_o[130] = lce_tr_resp_i[130];
  assign data_mem_pkt_o[129] = lce_tr_resp_i[129];
  assign data_mem_pkt_o[128] = lce_tr_resp_i[128];
  assign data_mem_pkt_o[127] = lce_tr_resp_i[127];
  assign data_mem_pkt_o[126] = lce_tr_resp_i[126];
  assign data_mem_pkt_o[125] = lce_tr_resp_i[125];
  assign data_mem_pkt_o[124] = lce_tr_resp_i[124];
  assign data_mem_pkt_o[123] = lce_tr_resp_i[123];
  assign data_mem_pkt_o[122] = lce_tr_resp_i[122];
  assign data_mem_pkt_o[121] = lce_tr_resp_i[121];
  assign data_mem_pkt_o[120] = lce_tr_resp_i[120];
  assign data_mem_pkt_o[119] = lce_tr_resp_i[119];
  assign data_mem_pkt_o[118] = lce_tr_resp_i[118];
  assign data_mem_pkt_o[117] = lce_tr_resp_i[117];
  assign data_mem_pkt_o[116] = lce_tr_resp_i[116];
  assign data_mem_pkt_o[115] = lce_tr_resp_i[115];
  assign data_mem_pkt_o[114] = lce_tr_resp_i[114];
  assign data_mem_pkt_o[113] = lce_tr_resp_i[113];
  assign data_mem_pkt_o[112] = lce_tr_resp_i[112];
  assign data_mem_pkt_o[111] = lce_tr_resp_i[111];
  assign data_mem_pkt_o[110] = lce_tr_resp_i[110];
  assign data_mem_pkt_o[109] = lce_tr_resp_i[109];
  assign data_mem_pkt_o[108] = lce_tr_resp_i[108];
  assign data_mem_pkt_o[107] = lce_tr_resp_i[107];
  assign data_mem_pkt_o[106] = lce_tr_resp_i[106];
  assign data_mem_pkt_o[105] = lce_tr_resp_i[105];
  assign data_mem_pkt_o[104] = lce_tr_resp_i[104];
  assign data_mem_pkt_o[103] = lce_tr_resp_i[103];
  assign data_mem_pkt_o[102] = lce_tr_resp_i[102];
  assign data_mem_pkt_o[101] = lce_tr_resp_i[101];
  assign data_mem_pkt_o[100] = lce_tr_resp_i[100];
  assign data_mem_pkt_o[99] = lce_tr_resp_i[99];
  assign data_mem_pkt_o[98] = lce_tr_resp_i[98];
  assign data_mem_pkt_o[97] = lce_tr_resp_i[97];
  assign data_mem_pkt_o[96] = lce_tr_resp_i[96];
  assign data_mem_pkt_o[95] = lce_tr_resp_i[95];
  assign data_mem_pkt_o[94] = lce_tr_resp_i[94];
  assign data_mem_pkt_o[93] = lce_tr_resp_i[93];
  assign data_mem_pkt_o[92] = lce_tr_resp_i[92];
  assign data_mem_pkt_o[91] = lce_tr_resp_i[91];
  assign data_mem_pkt_o[90] = lce_tr_resp_i[90];
  assign data_mem_pkt_o[89] = lce_tr_resp_i[89];
  assign data_mem_pkt_o[88] = lce_tr_resp_i[88];
  assign data_mem_pkt_o[87] = lce_tr_resp_i[87];
  assign data_mem_pkt_o[86] = lce_tr_resp_i[86];
  assign data_mem_pkt_o[85] = lce_tr_resp_i[85];
  assign data_mem_pkt_o[84] = lce_tr_resp_i[84];
  assign data_mem_pkt_o[83] = lce_tr_resp_i[83];
  assign data_mem_pkt_o[82] = lce_tr_resp_i[82];
  assign data_mem_pkt_o[81] = lce_tr_resp_i[81];
  assign data_mem_pkt_o[80] = lce_tr_resp_i[80];
  assign data_mem_pkt_o[79] = lce_tr_resp_i[79];
  assign data_mem_pkt_o[78] = lce_tr_resp_i[78];
  assign data_mem_pkt_o[77] = lce_tr_resp_i[77];
  assign data_mem_pkt_o[76] = lce_tr_resp_i[76];
  assign data_mem_pkt_o[75] = lce_tr_resp_i[75];
  assign data_mem_pkt_o[74] = lce_tr_resp_i[74];
  assign data_mem_pkt_o[73] = lce_tr_resp_i[73];
  assign data_mem_pkt_o[72] = lce_tr_resp_i[72];
  assign data_mem_pkt_o[71] = lce_tr_resp_i[71];
  assign data_mem_pkt_o[70] = lce_tr_resp_i[70];
  assign data_mem_pkt_o[69] = lce_tr_resp_i[69];
  assign data_mem_pkt_o[68] = lce_tr_resp_i[68];
  assign data_mem_pkt_o[67] = lce_tr_resp_i[67];
  assign data_mem_pkt_o[66] = lce_tr_resp_i[66];
  assign data_mem_pkt_o[65] = lce_tr_resp_i[65];
  assign data_mem_pkt_o[64] = lce_tr_resp_i[64];
  assign data_mem_pkt_o[63] = lce_tr_resp_i[63];
  assign data_mem_pkt_o[62] = lce_tr_resp_i[62];
  assign data_mem_pkt_o[61] = lce_tr_resp_i[61];
  assign data_mem_pkt_o[60] = lce_tr_resp_i[60];
  assign data_mem_pkt_o[59] = lce_tr_resp_i[59];
  assign data_mem_pkt_o[58] = lce_tr_resp_i[58];
  assign data_mem_pkt_o[57] = lce_tr_resp_i[57];
  assign data_mem_pkt_o[56] = lce_tr_resp_i[56];
  assign data_mem_pkt_o[55] = lce_tr_resp_i[55];
  assign data_mem_pkt_o[54] = lce_tr_resp_i[54];
  assign data_mem_pkt_o[53] = lce_tr_resp_i[53];
  assign data_mem_pkt_o[52] = lce_tr_resp_i[52];
  assign data_mem_pkt_o[51] = lce_tr_resp_i[51];
  assign data_mem_pkt_o[50] = lce_tr_resp_i[50];
  assign data_mem_pkt_o[49] = lce_tr_resp_i[49];
  assign data_mem_pkt_o[48] = lce_tr_resp_i[48];
  assign data_mem_pkt_o[47] = lce_tr_resp_i[47];
  assign data_mem_pkt_o[46] = lce_tr_resp_i[46];
  assign data_mem_pkt_o[45] = lce_tr_resp_i[45];
  assign data_mem_pkt_o[44] = lce_tr_resp_i[44];
  assign data_mem_pkt_o[43] = lce_tr_resp_i[43];
  assign data_mem_pkt_o[42] = lce_tr_resp_i[42];
  assign data_mem_pkt_o[41] = lce_tr_resp_i[41];
  assign data_mem_pkt_o[40] = lce_tr_resp_i[40];
  assign data_mem_pkt_o[39] = lce_tr_resp_i[39];
  assign data_mem_pkt_o[38] = lce_tr_resp_i[38];
  assign data_mem_pkt_o[37] = lce_tr_resp_i[37];
  assign data_mem_pkt_o[36] = lce_tr_resp_i[36];
  assign data_mem_pkt_o[35] = lce_tr_resp_i[35];
  assign data_mem_pkt_o[34] = lce_tr_resp_i[34];
  assign data_mem_pkt_o[33] = lce_tr_resp_i[33];
  assign data_mem_pkt_o[32] = lce_tr_resp_i[32];
  assign data_mem_pkt_o[31] = lce_tr_resp_i[31];
  assign data_mem_pkt_o[30] = lce_tr_resp_i[30];
  assign data_mem_pkt_o[29] = lce_tr_resp_i[29];
  assign data_mem_pkt_o[28] = lce_tr_resp_i[28];
  assign data_mem_pkt_o[27] = lce_tr_resp_i[27];
  assign data_mem_pkt_o[26] = lce_tr_resp_i[26];
  assign data_mem_pkt_o[25] = lce_tr_resp_i[25];
  assign data_mem_pkt_o[24] = lce_tr_resp_i[24];
  assign data_mem_pkt_o[23] = lce_tr_resp_i[23];
  assign data_mem_pkt_o[22] = lce_tr_resp_i[22];
  assign data_mem_pkt_o[21] = lce_tr_resp_i[21];
  assign data_mem_pkt_o[20] = lce_tr_resp_i[20];
  assign data_mem_pkt_o[19] = lce_tr_resp_i[19];
  assign data_mem_pkt_o[18] = lce_tr_resp_i[18];
  assign data_mem_pkt_o[17] = lce_tr_resp_i[17];
  assign data_mem_pkt_o[16] = lce_tr_resp_i[16];
  assign data_mem_pkt_o[15] = lce_tr_resp_i[15];
  assign data_mem_pkt_o[14] = lce_tr_resp_i[14];
  assign data_mem_pkt_o[13] = lce_tr_resp_i[13];
  assign data_mem_pkt_o[12] = lce_tr_resp_i[12];
  assign data_mem_pkt_o[11] = lce_tr_resp_i[11];
  assign data_mem_pkt_o[10] = lce_tr_resp_i[10];
  assign data_mem_pkt_o[9] = lce_tr_resp_i[9];
  assign data_mem_pkt_o[8] = lce_tr_resp_i[8];
  assign data_mem_pkt_o[7] = lce_tr_resp_i[7];
  assign data_mem_pkt_o[6] = lce_tr_resp_i[6];
  assign data_mem_pkt_o[5] = lce_tr_resp_i[5];
  assign data_mem_pkt_o[4] = lce_tr_resp_i[4];
  assign data_mem_pkt_o[3] = lce_tr_resp_i[3];
  assign data_mem_pkt_o[2] = lce_tr_resp_i[2];
  assign data_mem_pkt_o[1] = lce_tr_resp_i[1];
  assign data_mem_pkt_o[0] = lce_tr_resp_i[0];
  assign lce_tr_resp_yumi_o = data_mem_pkt_yumi_i & lce_tr_resp_v_i;
  assign tr_received_o = data_mem_pkt_yumi_i & lce_tr_resp_v_i;

endmodule



module bp_fe_sub_module1
(
  clk_i,
  reset_i,
  id_i,
  ready_o,
  cache_miss_o,
  miss_i,
  miss_addr_i,
  data_mem_data_i,
  data_mem_pkt_o,
  data_mem_pkt_v_o,
  data_mem_pkt_yumi_i,
  tag_mem_pkt_o,
  tag_mem_pkt_v_o,
  tag_mem_pkt_yumi_i,
  metadata_mem_pkt_v_o,
  metadata_mem_pkt_o,
  lru_way_i,
  metadata_mem_pkt_yumi_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  lce_tr_resp_i,
  lce_tr_resp_v_i,
  lce_tr_resp_ready_o,
  lce_tr_resp_o,
  lce_tr_resp_v_o,
  lce_tr_resp_ready_i
);

  input [0:0] id_i;
  input [21:0] miss_addr_i;
  input [511:0] data_mem_data_i;
  output [521:0] data_mem_pkt_o;
  output [22:0] tag_mem_pkt_o;
  output [9:0] metadata_mem_pkt_o;
  input [2:0] lru_way_i;
  output [29:0] lce_req_o;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  input [35:0] lce_cmd_i;
  input [539:0] lce_data_cmd_i;
  input [538:0] lce_tr_resp_i;
  output [538:0] lce_tr_resp_o;
  input clk_i;
  input reset_i;
  input miss_i;
  input data_mem_pkt_yumi_i;
  input tag_mem_pkt_yumi_i;
  input metadata_mem_pkt_yumi_i;
  input lce_req_ready_i;
  input lce_resp_ready_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_v_i;
  input lce_tr_resp_v_i;
  input lce_tr_resp_ready_i;
  output ready_o;
  output cache_miss_o;
  output data_mem_pkt_v_o;
  output tag_mem_pkt_v_o;
  output metadata_mem_pkt_v_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_ready_o;
  output lce_data_cmd_ready_o;
  output lce_tr_resp_ready_o;
  output lce_tr_resp_v_o;
  wire [521:0] data_mem_pkt_o,lce_cmd_data_mem_pkt_lo,lce_data_cmd_data_mem_pkt_lo,
  lce_tr_resp_in_data_mem_pkt_lo;
  wire [22:0] tag_mem_pkt_o;
  wire [9:0] metadata_mem_pkt_o;
  wire [29:0] lce_req_o;
  wire [25:0] lce_resp_o,lce_req_lce_resp_lo,lce_cmd_lce_resp_lo;
  wire [536:0] lce_data_resp_o;
  wire [538:0] lce_tr_resp_o,lce_tr_resp_in_fifo_data_lo;
  wire ready_o,cache_miss_o,data_mem_pkt_v_o,tag_mem_pkt_v_o,metadata_mem_pkt_v_o,
  lce_req_v_o,lce_resp_v_o,lce_data_resp_v_o,lce_cmd_ready_o,lce_data_cmd_ready_o,
  lce_tr_resp_ready_o,lce_tr_resp_v_o,N0,N1,N2,N3,N4,N5,tr_received_li,
  cce_data_received_li,tag_set_li,tag_set_wakeup_li,lce_req_lce_resp_v_lo,
  lce_req_lce_resp_yumi_li,lce_cmd_fifo_v_lo,lce_cmd_fifo_yumi_li,lce_ready_lo,lce_cmd_data_mem_pkt_v_lo,
  lce_cmd_data_mem_pkt_yumi_li,lce_cmd_lce_resp_v_lo,lce_cmd_lce_resp_yumi_li,
  lce_data_cmd_fifo_v_lo,lce_data_cmd_fifo_yumi_li,lce_data_cmd_data_mem_pkt_v_lo,
  lce_data_cmd_data_mem_pkt_yumi_li,lce_tr_resp_in_fifo_v_lo,
  lce_tr_resp_in_fifo_yumi_li,lce_tr_resp_in_data_mem_pkt_v_lo,lce_tr_resp_in_data_mem_pkt_yumi_li,N6,N7,N8,
  N9,N10,N11,N12,N13,N14;
  wire [35:0] lce_cmd_fifo_data_lo;
  wire [539:0] lce_data_cmd_fifo_data_lo;

  bp_fe_lce_req_data_width_p64_lce_addr_width_p22_num_cce_p1_num_lce_p2_lce_sets_p64_ways_p8_block_size_in_bytes_p8
  lce_req
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .id_i(id_i[0]),
    .miss_i(miss_i),
    .miss_addr_i(miss_addr_i),
    .lru_way_i(lru_way_i),
    .cache_miss_o(cache_miss_o),
    .tr_received_i(tr_received_li),
    .cce_data_received_i(cce_data_received_li),
    .tag_set_i(tag_set_li),
    .tag_set_wakeup_i(tag_set_wakeup_li),
    .lce_req_o(lce_req_o),
    .lce_req_v_o(lce_req_v_o),
    .lce_req_ready_i(lce_req_ready_i),
    .lce_resp_o(lce_req_lce_resp_lo),
    .lce_resp_v_o(lce_req_lce_resp_v_lo),
    .lce_resp_yumi_i(lce_req_lce_resp_yumi_li)
  );


  bsg_two_fifo_width_p36
  lce_cmd_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(lce_cmd_ready_o),
    .data_i(lce_cmd_i),
    .v_i(lce_cmd_v_i),
    .v_o(lce_cmd_fifo_v_lo),
    .data_o(lce_cmd_fifo_data_lo),
    .yumi_i(lce_cmd_fifo_yumi_li)
  );


  bp_fe_lce_cmd_data_width_p64_lce_data_width_p512_lce_addr_width_p22_lce_sets_p64_ways_p8_tag_width_p10_num_cce_p1_num_lce_p2_block_size_in_bytes_p8
  lce_cmd
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .id_i(id_i[0]),
    .lce_ready_o(lce_ready_lo),
    .tag_set_o(tag_set_li),
    .tag_set_wakeup_o(tag_set_wakeup_li),
    .data_mem_data_i(data_mem_data_i),
    .data_mem_pkt_o(lce_cmd_data_mem_pkt_lo),
    .data_mem_pkt_v_o(lce_cmd_data_mem_pkt_v_lo),
    .data_mem_pkt_yumi_i(lce_cmd_data_mem_pkt_yumi_li),
    .tag_mem_pkt_o(tag_mem_pkt_o),
    .tag_mem_pkt_v_o(tag_mem_pkt_v_o),
    .tag_mem_pkt_yumi_i(tag_mem_pkt_yumi_i),
    .metadata_mem_pkt_v_o(metadata_mem_pkt_v_o),
    .metadata_mem_pkt_o(metadata_mem_pkt_o),
    .metadata_mem_pkt_yumi_i(metadata_mem_pkt_yumi_i),
    .lce_resp_o(lce_cmd_lce_resp_lo),
    .lce_resp_v_o(lce_cmd_lce_resp_v_lo),
    .lce_resp_yumi_i(lce_cmd_lce_resp_yumi_li),
    .lce_data_resp_o(lce_data_resp_o),
    .lce_data_resp_v_o(lce_data_resp_v_o),
    .lce_data_resp_ready_i(lce_data_resp_ready_i),
    .lce_cmd_i(lce_cmd_fifo_data_lo),
    .lce_cmd_v_i(lce_cmd_fifo_v_lo),
    .lce_cmd_yumi_o(lce_cmd_fifo_yumi_li),
    .lce_tr_resp_o(lce_tr_resp_o),
    .lce_tr_resp_v_o(lce_tr_resp_v_o),
    .lce_tr_resp_ready_i(lce_tr_resp_ready_i)
  );


  bsg_two_fifo_width_p540
  lce_data_cmd_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(lce_data_cmd_ready_o),
    .data_i(lce_data_cmd_i),
    .v_i(lce_data_cmd_v_i),
    .v_o(lce_data_cmd_fifo_v_lo),
    .data_o(lce_data_cmd_fifo_data_lo),
    .yumi_i(lce_data_cmd_fifo_yumi_li)
  );


  bp_fe_lce_data_cmd_data_width_p64_lce_addr_width_p22_lce_data_width_p512_num_cce_p1_num_lce_p2_lce_sets_p64_ways_p8_block_size_in_bytes_p8
  lce_data_cmd
  (
    .cce_data_received_o(cce_data_received_li),
    .lce_data_cmd_i(lce_data_cmd_fifo_data_lo),
    .lce_data_cmd_v_i(lce_data_cmd_fifo_v_lo),
    .lce_data_cmd_yumi_o(lce_data_cmd_fifo_yumi_li),
    .data_mem_pkt_v_o(lce_data_cmd_data_mem_pkt_v_lo),
    .data_mem_pkt_o(lce_data_cmd_data_mem_pkt_lo),
    .data_mem_pkt_yumi_i(lce_data_cmd_data_mem_pkt_yumi_li)
  );


  bsg_two_fifo_width_p539
  lce_tr_resp_in_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(lce_tr_resp_ready_o),
    .data_i(lce_tr_resp_i),
    .v_i(lce_tr_resp_v_i),
    .v_o(lce_tr_resp_in_fifo_v_lo),
    .data_o(lce_tr_resp_in_fifo_data_lo),
    .yumi_i(lce_tr_resp_in_fifo_yumi_li)
  );


  bp_fe_lce_tr_resp_in_data_width_p64_lce_data_width_p512_lce_addr_width_p22_lce_sets_p64_ways_p8_num_cce_p1_num_lce_p2_block_size_in_bytes_p8
  lce_tr_resp_in
  (
    .tr_received_o(tr_received_li),
    .lce_tr_resp_i(lce_tr_resp_in_fifo_data_lo),
    .lce_tr_resp_v_i(lce_tr_resp_in_fifo_v_lo),
    .lce_tr_resp_yumi_o(lce_tr_resp_in_fifo_yumi_li),
    .data_mem_pkt_v_o(lce_tr_resp_in_data_mem_pkt_v_lo),
    .data_mem_pkt_o(lce_tr_resp_in_data_mem_pkt_lo),
    .data_mem_pkt_yumi_i(lce_tr_resp_in_data_mem_pkt_yumi_li)
  );

  assign data_mem_pkt_v_o = (N0)? 1'b1 : 
                            (N9)? 1'b1 : 
                            (N7)? lce_cmd_data_mem_pkt_v_lo : 1'b0;
  assign N0 = lce_tr_resp_in_data_mem_pkt_v_lo;
  assign data_mem_pkt_o = (N0)? lce_tr_resp_in_data_mem_pkt_lo : 
                          (N9)? lce_data_cmd_data_mem_pkt_lo : 
                          (N7)? lce_cmd_data_mem_pkt_lo : 1'b0;
  assign lce_tr_resp_in_data_mem_pkt_yumi_li = (N0)? data_mem_pkt_yumi_i : 
                                               (N8)? 1'b0 : 
                                               (N1)? 1'b0 : 1'b0;
  assign N1 = 1'b0;
  assign lce_data_cmd_data_mem_pkt_yumi_li = (N0)? 1'b0 : 
                                             (N9)? data_mem_pkt_yumi_i : 
                                             (N7)? 1'b0 : 1'b0;
  assign lce_cmd_data_mem_pkt_yumi_li = (N0)? 1'b0 : 
                                        (N9)? 1'b0 : 
                                        (N7)? data_mem_pkt_yumi_i : 1'b0;
  assign lce_resp_v_o = (N2)? 1'b1 : 
                        (N3)? lce_cmd_lce_resp_v_lo : 1'b0;
  assign N2 = lce_req_lce_resp_v_lo;
  assign N3 = N10;
  assign lce_resp_o = (N2)? lce_req_lce_resp_lo : 
                      (N3)? lce_cmd_lce_resp_lo : 1'b0;
  assign lce_req_lce_resp_yumi_li = (N2)? lce_resp_ready_i : 
                                    (N3)? 1'b0 : 1'b0;
  assign lce_cmd_lce_resp_yumi_li = (N4)? lce_resp_ready_i : 
                                    (N5)? 1'b0 : 1'b0;
  assign N4 = lce_cmd_lce_resp_v_lo;
  assign N5 = N11;
  assign N6 = lce_data_cmd_data_mem_pkt_v_lo | lce_tr_resp_in_data_mem_pkt_v_lo;
  assign N7 = ~N6;
  assign N8 = ~lce_tr_resp_in_data_mem_pkt_v_lo;
  assign N9 = lce_data_cmd_data_mem_pkt_v_lo & N8;
  assign N10 = ~lce_req_lce_resp_v_lo;
  assign N11 = ~lce_cmd_lce_resp_v_lo;
  assign ready_o = N13 & N14;
  assign N13 = lce_ready_lo & N12;
  assign N12 = ~1'b0;
  assign N14 = ~cache_miss_o;

endmodule



module bsg_mux_width_p64_els_p8
(
  data_i,
  sel_i,
  data_o
);

  input [511:0] data_i;
  input [2:0] sel_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;
  assign data_o[63] = (N7)? data_i[63] : 
                      (N9)? data_i[127] : 
                      (N11)? data_i[191] : 
                      (N13)? data_i[255] : 
                      (N8)? data_i[319] : 
                      (N10)? data_i[383] : 
                      (N12)? data_i[447] : 
                      (N14)? data_i[511] : 1'b0;
  assign data_o[62] = (N7)? data_i[62] : 
                      (N9)? data_i[126] : 
                      (N11)? data_i[190] : 
                      (N13)? data_i[254] : 
                      (N8)? data_i[318] : 
                      (N10)? data_i[382] : 
                      (N12)? data_i[446] : 
                      (N14)? data_i[510] : 1'b0;
  assign data_o[61] = (N7)? data_i[61] : 
                      (N9)? data_i[125] : 
                      (N11)? data_i[189] : 
                      (N13)? data_i[253] : 
                      (N8)? data_i[317] : 
                      (N10)? data_i[381] : 
                      (N12)? data_i[445] : 
                      (N14)? data_i[509] : 1'b0;
  assign data_o[60] = (N7)? data_i[60] : 
                      (N9)? data_i[124] : 
                      (N11)? data_i[188] : 
                      (N13)? data_i[252] : 
                      (N8)? data_i[316] : 
                      (N10)? data_i[380] : 
                      (N12)? data_i[444] : 
                      (N14)? data_i[508] : 1'b0;
  assign data_o[59] = (N7)? data_i[59] : 
                      (N9)? data_i[123] : 
                      (N11)? data_i[187] : 
                      (N13)? data_i[251] : 
                      (N8)? data_i[315] : 
                      (N10)? data_i[379] : 
                      (N12)? data_i[443] : 
                      (N14)? data_i[507] : 1'b0;
  assign data_o[58] = (N7)? data_i[58] : 
                      (N9)? data_i[122] : 
                      (N11)? data_i[186] : 
                      (N13)? data_i[250] : 
                      (N8)? data_i[314] : 
                      (N10)? data_i[378] : 
                      (N12)? data_i[442] : 
                      (N14)? data_i[506] : 1'b0;
  assign data_o[57] = (N7)? data_i[57] : 
                      (N9)? data_i[121] : 
                      (N11)? data_i[185] : 
                      (N13)? data_i[249] : 
                      (N8)? data_i[313] : 
                      (N10)? data_i[377] : 
                      (N12)? data_i[441] : 
                      (N14)? data_i[505] : 1'b0;
  assign data_o[56] = (N7)? data_i[56] : 
                      (N9)? data_i[120] : 
                      (N11)? data_i[184] : 
                      (N13)? data_i[248] : 
                      (N8)? data_i[312] : 
                      (N10)? data_i[376] : 
                      (N12)? data_i[440] : 
                      (N14)? data_i[504] : 1'b0;
  assign data_o[55] = (N7)? data_i[55] : 
                      (N9)? data_i[119] : 
                      (N11)? data_i[183] : 
                      (N13)? data_i[247] : 
                      (N8)? data_i[311] : 
                      (N10)? data_i[375] : 
                      (N12)? data_i[439] : 
                      (N14)? data_i[503] : 1'b0;
  assign data_o[54] = (N7)? data_i[54] : 
                      (N9)? data_i[118] : 
                      (N11)? data_i[182] : 
                      (N13)? data_i[246] : 
                      (N8)? data_i[310] : 
                      (N10)? data_i[374] : 
                      (N12)? data_i[438] : 
                      (N14)? data_i[502] : 1'b0;
  assign data_o[53] = (N7)? data_i[53] : 
                      (N9)? data_i[117] : 
                      (N11)? data_i[181] : 
                      (N13)? data_i[245] : 
                      (N8)? data_i[309] : 
                      (N10)? data_i[373] : 
                      (N12)? data_i[437] : 
                      (N14)? data_i[501] : 1'b0;
  assign data_o[52] = (N7)? data_i[52] : 
                      (N9)? data_i[116] : 
                      (N11)? data_i[180] : 
                      (N13)? data_i[244] : 
                      (N8)? data_i[308] : 
                      (N10)? data_i[372] : 
                      (N12)? data_i[436] : 
                      (N14)? data_i[500] : 1'b0;
  assign data_o[51] = (N7)? data_i[51] : 
                      (N9)? data_i[115] : 
                      (N11)? data_i[179] : 
                      (N13)? data_i[243] : 
                      (N8)? data_i[307] : 
                      (N10)? data_i[371] : 
                      (N12)? data_i[435] : 
                      (N14)? data_i[499] : 1'b0;
  assign data_o[50] = (N7)? data_i[50] : 
                      (N9)? data_i[114] : 
                      (N11)? data_i[178] : 
                      (N13)? data_i[242] : 
                      (N8)? data_i[306] : 
                      (N10)? data_i[370] : 
                      (N12)? data_i[434] : 
                      (N14)? data_i[498] : 1'b0;
  assign data_o[49] = (N7)? data_i[49] : 
                      (N9)? data_i[113] : 
                      (N11)? data_i[177] : 
                      (N13)? data_i[241] : 
                      (N8)? data_i[305] : 
                      (N10)? data_i[369] : 
                      (N12)? data_i[433] : 
                      (N14)? data_i[497] : 1'b0;
  assign data_o[48] = (N7)? data_i[48] : 
                      (N9)? data_i[112] : 
                      (N11)? data_i[176] : 
                      (N13)? data_i[240] : 
                      (N8)? data_i[304] : 
                      (N10)? data_i[368] : 
                      (N12)? data_i[432] : 
                      (N14)? data_i[496] : 1'b0;
  assign data_o[47] = (N7)? data_i[47] : 
                      (N9)? data_i[111] : 
                      (N11)? data_i[175] : 
                      (N13)? data_i[239] : 
                      (N8)? data_i[303] : 
                      (N10)? data_i[367] : 
                      (N12)? data_i[431] : 
                      (N14)? data_i[495] : 1'b0;
  assign data_o[46] = (N7)? data_i[46] : 
                      (N9)? data_i[110] : 
                      (N11)? data_i[174] : 
                      (N13)? data_i[238] : 
                      (N8)? data_i[302] : 
                      (N10)? data_i[366] : 
                      (N12)? data_i[430] : 
                      (N14)? data_i[494] : 1'b0;
  assign data_o[45] = (N7)? data_i[45] : 
                      (N9)? data_i[109] : 
                      (N11)? data_i[173] : 
                      (N13)? data_i[237] : 
                      (N8)? data_i[301] : 
                      (N10)? data_i[365] : 
                      (N12)? data_i[429] : 
                      (N14)? data_i[493] : 1'b0;
  assign data_o[44] = (N7)? data_i[44] : 
                      (N9)? data_i[108] : 
                      (N11)? data_i[172] : 
                      (N13)? data_i[236] : 
                      (N8)? data_i[300] : 
                      (N10)? data_i[364] : 
                      (N12)? data_i[428] : 
                      (N14)? data_i[492] : 1'b0;
  assign data_o[43] = (N7)? data_i[43] : 
                      (N9)? data_i[107] : 
                      (N11)? data_i[171] : 
                      (N13)? data_i[235] : 
                      (N8)? data_i[299] : 
                      (N10)? data_i[363] : 
                      (N12)? data_i[427] : 
                      (N14)? data_i[491] : 1'b0;
  assign data_o[42] = (N7)? data_i[42] : 
                      (N9)? data_i[106] : 
                      (N11)? data_i[170] : 
                      (N13)? data_i[234] : 
                      (N8)? data_i[298] : 
                      (N10)? data_i[362] : 
                      (N12)? data_i[426] : 
                      (N14)? data_i[490] : 1'b0;
  assign data_o[41] = (N7)? data_i[41] : 
                      (N9)? data_i[105] : 
                      (N11)? data_i[169] : 
                      (N13)? data_i[233] : 
                      (N8)? data_i[297] : 
                      (N10)? data_i[361] : 
                      (N12)? data_i[425] : 
                      (N14)? data_i[489] : 1'b0;
  assign data_o[40] = (N7)? data_i[40] : 
                      (N9)? data_i[104] : 
                      (N11)? data_i[168] : 
                      (N13)? data_i[232] : 
                      (N8)? data_i[296] : 
                      (N10)? data_i[360] : 
                      (N12)? data_i[424] : 
                      (N14)? data_i[488] : 1'b0;
  assign data_o[39] = (N7)? data_i[39] : 
                      (N9)? data_i[103] : 
                      (N11)? data_i[167] : 
                      (N13)? data_i[231] : 
                      (N8)? data_i[295] : 
                      (N10)? data_i[359] : 
                      (N12)? data_i[423] : 
                      (N14)? data_i[487] : 1'b0;
  assign data_o[38] = (N7)? data_i[38] : 
                      (N9)? data_i[102] : 
                      (N11)? data_i[166] : 
                      (N13)? data_i[230] : 
                      (N8)? data_i[294] : 
                      (N10)? data_i[358] : 
                      (N12)? data_i[422] : 
                      (N14)? data_i[486] : 1'b0;
  assign data_o[37] = (N7)? data_i[37] : 
                      (N9)? data_i[101] : 
                      (N11)? data_i[165] : 
                      (N13)? data_i[229] : 
                      (N8)? data_i[293] : 
                      (N10)? data_i[357] : 
                      (N12)? data_i[421] : 
                      (N14)? data_i[485] : 1'b0;
  assign data_o[36] = (N7)? data_i[36] : 
                      (N9)? data_i[100] : 
                      (N11)? data_i[164] : 
                      (N13)? data_i[228] : 
                      (N8)? data_i[292] : 
                      (N10)? data_i[356] : 
                      (N12)? data_i[420] : 
                      (N14)? data_i[484] : 1'b0;
  assign data_o[35] = (N7)? data_i[35] : 
                      (N9)? data_i[99] : 
                      (N11)? data_i[163] : 
                      (N13)? data_i[227] : 
                      (N8)? data_i[291] : 
                      (N10)? data_i[355] : 
                      (N12)? data_i[419] : 
                      (N14)? data_i[483] : 1'b0;
  assign data_o[34] = (N7)? data_i[34] : 
                      (N9)? data_i[98] : 
                      (N11)? data_i[162] : 
                      (N13)? data_i[226] : 
                      (N8)? data_i[290] : 
                      (N10)? data_i[354] : 
                      (N12)? data_i[418] : 
                      (N14)? data_i[482] : 1'b0;
  assign data_o[33] = (N7)? data_i[33] : 
                      (N9)? data_i[97] : 
                      (N11)? data_i[161] : 
                      (N13)? data_i[225] : 
                      (N8)? data_i[289] : 
                      (N10)? data_i[353] : 
                      (N12)? data_i[417] : 
                      (N14)? data_i[481] : 1'b0;
  assign data_o[32] = (N7)? data_i[32] : 
                      (N9)? data_i[96] : 
                      (N11)? data_i[160] : 
                      (N13)? data_i[224] : 
                      (N8)? data_i[288] : 
                      (N10)? data_i[352] : 
                      (N12)? data_i[416] : 
                      (N14)? data_i[480] : 1'b0;
  assign data_o[31] = (N7)? data_i[31] : 
                      (N9)? data_i[95] : 
                      (N11)? data_i[159] : 
                      (N13)? data_i[223] : 
                      (N8)? data_i[287] : 
                      (N10)? data_i[351] : 
                      (N12)? data_i[415] : 
                      (N14)? data_i[479] : 1'b0;
  assign data_o[30] = (N7)? data_i[30] : 
                      (N9)? data_i[94] : 
                      (N11)? data_i[158] : 
                      (N13)? data_i[222] : 
                      (N8)? data_i[286] : 
                      (N10)? data_i[350] : 
                      (N12)? data_i[414] : 
                      (N14)? data_i[478] : 1'b0;
  assign data_o[29] = (N7)? data_i[29] : 
                      (N9)? data_i[93] : 
                      (N11)? data_i[157] : 
                      (N13)? data_i[221] : 
                      (N8)? data_i[285] : 
                      (N10)? data_i[349] : 
                      (N12)? data_i[413] : 
                      (N14)? data_i[477] : 1'b0;
  assign data_o[28] = (N7)? data_i[28] : 
                      (N9)? data_i[92] : 
                      (N11)? data_i[156] : 
                      (N13)? data_i[220] : 
                      (N8)? data_i[284] : 
                      (N10)? data_i[348] : 
                      (N12)? data_i[412] : 
                      (N14)? data_i[476] : 1'b0;
  assign data_o[27] = (N7)? data_i[27] : 
                      (N9)? data_i[91] : 
                      (N11)? data_i[155] : 
                      (N13)? data_i[219] : 
                      (N8)? data_i[283] : 
                      (N10)? data_i[347] : 
                      (N12)? data_i[411] : 
                      (N14)? data_i[475] : 1'b0;
  assign data_o[26] = (N7)? data_i[26] : 
                      (N9)? data_i[90] : 
                      (N11)? data_i[154] : 
                      (N13)? data_i[218] : 
                      (N8)? data_i[282] : 
                      (N10)? data_i[346] : 
                      (N12)? data_i[410] : 
                      (N14)? data_i[474] : 1'b0;
  assign data_o[25] = (N7)? data_i[25] : 
                      (N9)? data_i[89] : 
                      (N11)? data_i[153] : 
                      (N13)? data_i[217] : 
                      (N8)? data_i[281] : 
                      (N10)? data_i[345] : 
                      (N12)? data_i[409] : 
                      (N14)? data_i[473] : 1'b0;
  assign data_o[24] = (N7)? data_i[24] : 
                      (N9)? data_i[88] : 
                      (N11)? data_i[152] : 
                      (N13)? data_i[216] : 
                      (N8)? data_i[280] : 
                      (N10)? data_i[344] : 
                      (N12)? data_i[408] : 
                      (N14)? data_i[472] : 1'b0;
  assign data_o[23] = (N7)? data_i[23] : 
                      (N9)? data_i[87] : 
                      (N11)? data_i[151] : 
                      (N13)? data_i[215] : 
                      (N8)? data_i[279] : 
                      (N10)? data_i[343] : 
                      (N12)? data_i[407] : 
                      (N14)? data_i[471] : 1'b0;
  assign data_o[22] = (N7)? data_i[22] : 
                      (N9)? data_i[86] : 
                      (N11)? data_i[150] : 
                      (N13)? data_i[214] : 
                      (N8)? data_i[278] : 
                      (N10)? data_i[342] : 
                      (N12)? data_i[406] : 
                      (N14)? data_i[470] : 1'b0;
  assign data_o[21] = (N7)? data_i[21] : 
                      (N9)? data_i[85] : 
                      (N11)? data_i[149] : 
                      (N13)? data_i[213] : 
                      (N8)? data_i[277] : 
                      (N10)? data_i[341] : 
                      (N12)? data_i[405] : 
                      (N14)? data_i[469] : 1'b0;
  assign data_o[20] = (N7)? data_i[20] : 
                      (N9)? data_i[84] : 
                      (N11)? data_i[148] : 
                      (N13)? data_i[212] : 
                      (N8)? data_i[276] : 
                      (N10)? data_i[340] : 
                      (N12)? data_i[404] : 
                      (N14)? data_i[468] : 1'b0;
  assign data_o[19] = (N7)? data_i[19] : 
                      (N9)? data_i[83] : 
                      (N11)? data_i[147] : 
                      (N13)? data_i[211] : 
                      (N8)? data_i[275] : 
                      (N10)? data_i[339] : 
                      (N12)? data_i[403] : 
                      (N14)? data_i[467] : 1'b0;
  assign data_o[18] = (N7)? data_i[18] : 
                      (N9)? data_i[82] : 
                      (N11)? data_i[146] : 
                      (N13)? data_i[210] : 
                      (N8)? data_i[274] : 
                      (N10)? data_i[338] : 
                      (N12)? data_i[402] : 
                      (N14)? data_i[466] : 1'b0;
  assign data_o[17] = (N7)? data_i[17] : 
                      (N9)? data_i[81] : 
                      (N11)? data_i[145] : 
                      (N13)? data_i[209] : 
                      (N8)? data_i[273] : 
                      (N10)? data_i[337] : 
                      (N12)? data_i[401] : 
                      (N14)? data_i[465] : 1'b0;
  assign data_o[16] = (N7)? data_i[16] : 
                      (N9)? data_i[80] : 
                      (N11)? data_i[144] : 
                      (N13)? data_i[208] : 
                      (N8)? data_i[272] : 
                      (N10)? data_i[336] : 
                      (N12)? data_i[400] : 
                      (N14)? data_i[464] : 1'b0;
  assign data_o[15] = (N7)? data_i[15] : 
                      (N9)? data_i[79] : 
                      (N11)? data_i[143] : 
                      (N13)? data_i[207] : 
                      (N8)? data_i[271] : 
                      (N10)? data_i[335] : 
                      (N12)? data_i[399] : 
                      (N14)? data_i[463] : 1'b0;
  assign data_o[14] = (N7)? data_i[14] : 
                      (N9)? data_i[78] : 
                      (N11)? data_i[142] : 
                      (N13)? data_i[206] : 
                      (N8)? data_i[270] : 
                      (N10)? data_i[334] : 
                      (N12)? data_i[398] : 
                      (N14)? data_i[462] : 1'b0;
  assign data_o[13] = (N7)? data_i[13] : 
                      (N9)? data_i[77] : 
                      (N11)? data_i[141] : 
                      (N13)? data_i[205] : 
                      (N8)? data_i[269] : 
                      (N10)? data_i[333] : 
                      (N12)? data_i[397] : 
                      (N14)? data_i[461] : 1'b0;
  assign data_o[12] = (N7)? data_i[12] : 
                      (N9)? data_i[76] : 
                      (N11)? data_i[140] : 
                      (N13)? data_i[204] : 
                      (N8)? data_i[268] : 
                      (N10)? data_i[332] : 
                      (N12)? data_i[396] : 
                      (N14)? data_i[460] : 1'b0;
  assign data_o[11] = (N7)? data_i[11] : 
                      (N9)? data_i[75] : 
                      (N11)? data_i[139] : 
                      (N13)? data_i[203] : 
                      (N8)? data_i[267] : 
                      (N10)? data_i[331] : 
                      (N12)? data_i[395] : 
                      (N14)? data_i[459] : 1'b0;
  assign data_o[10] = (N7)? data_i[10] : 
                      (N9)? data_i[74] : 
                      (N11)? data_i[138] : 
                      (N13)? data_i[202] : 
                      (N8)? data_i[266] : 
                      (N10)? data_i[330] : 
                      (N12)? data_i[394] : 
                      (N14)? data_i[458] : 1'b0;
  assign data_o[9] = (N7)? data_i[9] : 
                     (N9)? data_i[73] : 
                     (N11)? data_i[137] : 
                     (N13)? data_i[201] : 
                     (N8)? data_i[265] : 
                     (N10)? data_i[329] : 
                     (N12)? data_i[393] : 
                     (N14)? data_i[457] : 1'b0;
  assign data_o[8] = (N7)? data_i[8] : 
                     (N9)? data_i[72] : 
                     (N11)? data_i[136] : 
                     (N13)? data_i[200] : 
                     (N8)? data_i[264] : 
                     (N10)? data_i[328] : 
                     (N12)? data_i[392] : 
                     (N14)? data_i[456] : 1'b0;
  assign data_o[7] = (N7)? data_i[7] : 
                     (N9)? data_i[71] : 
                     (N11)? data_i[135] : 
                     (N13)? data_i[199] : 
                     (N8)? data_i[263] : 
                     (N10)? data_i[327] : 
                     (N12)? data_i[391] : 
                     (N14)? data_i[455] : 1'b0;
  assign data_o[6] = (N7)? data_i[6] : 
                     (N9)? data_i[70] : 
                     (N11)? data_i[134] : 
                     (N13)? data_i[198] : 
                     (N8)? data_i[262] : 
                     (N10)? data_i[326] : 
                     (N12)? data_i[390] : 
                     (N14)? data_i[454] : 1'b0;
  assign data_o[5] = (N7)? data_i[5] : 
                     (N9)? data_i[69] : 
                     (N11)? data_i[133] : 
                     (N13)? data_i[197] : 
                     (N8)? data_i[261] : 
                     (N10)? data_i[325] : 
                     (N12)? data_i[389] : 
                     (N14)? data_i[453] : 1'b0;
  assign data_o[4] = (N7)? data_i[4] : 
                     (N9)? data_i[68] : 
                     (N11)? data_i[132] : 
                     (N13)? data_i[196] : 
                     (N8)? data_i[260] : 
                     (N10)? data_i[324] : 
                     (N12)? data_i[388] : 
                     (N14)? data_i[452] : 1'b0;
  assign data_o[3] = (N7)? data_i[3] : 
                     (N9)? data_i[67] : 
                     (N11)? data_i[131] : 
                     (N13)? data_i[195] : 
                     (N8)? data_i[259] : 
                     (N10)? data_i[323] : 
                     (N12)? data_i[387] : 
                     (N14)? data_i[451] : 1'b0;
  assign data_o[2] = (N7)? data_i[2] : 
                     (N9)? data_i[66] : 
                     (N11)? data_i[130] : 
                     (N13)? data_i[194] : 
                     (N8)? data_i[258] : 
                     (N10)? data_i[322] : 
                     (N12)? data_i[386] : 
                     (N14)? data_i[450] : 1'b0;
  assign data_o[1] = (N7)? data_i[1] : 
                     (N9)? data_i[65] : 
                     (N11)? data_i[129] : 
                     (N13)? data_i[193] : 
                     (N8)? data_i[257] : 
                     (N10)? data_i[321] : 
                     (N12)? data_i[385] : 
                     (N14)? data_i[449] : 1'b0;
  assign data_o[0] = (N7)? data_i[0] : 
                     (N9)? data_i[64] : 
                     (N11)? data_i[128] : 
                     (N13)? data_i[192] : 
                     (N8)? data_i[256] : 
                     (N10)? data_i[320] : 
                     (N12)? data_i[384] : 
                     (N14)? data_i[448] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];
  assign N6 = ~sel_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & sel_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & sel_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & sel_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & sel_i[2];

endmodule



module bp_be_dcache_lru_decode_ways_p8
(
  way_id_i,
  data_o,
  mask_o
);

  input [2:0] way_id_i;
  output [6:0] data_o;
  output [6:0] mask_o;
  wire [6:0] data_o,mask_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30;
  assign mask_o[0] = 1'b1;
  assign N11 = N8 & N9;
  assign N12 = N11 & N10;
  assign N13 = way_id_i[2] | way_id_i[1];
  assign N14 = N13 | N10;
  assign N16 = way_id_i[2] | N9;
  assign N17 = N16 | way_id_i[0];
  assign N19 = N16 | N10;
  assign N21 = N8 | way_id_i[1];
  assign N22 = N21 | way_id_i[0];
  assign N24 = N21 | N10;
  assign N26 = N8 | N9;
  assign N27 = N26 | way_id_i[0];
  assign N29 = way_id_i[2] & way_id_i[1];
  assign N30 = N29 & way_id_i[0];
  assign data_o = (N0)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                  (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                  (N2)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                  (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                  (N4)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                  (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                  (N6)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                  (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N12;
  assign N1 = N15;
  assign N2 = N18;
  assign N3 = N20;
  assign N4 = N23;
  assign N5 = N25;
  assign N6 = N28;
  assign N7 = N30;
  assign mask_o[6:1] = (N0)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                       (N1)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                       (N2)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                       (N3)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                       (N4)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                       (N5)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                       (N6)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                       (N7)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 1'b0;
  assign N8 = ~way_id_i[2];
  assign N9 = ~way_id_i[1];
  assign N10 = ~way_id_i[0];
  assign N15 = ~N14;
  assign N18 = ~N17;
  assign N20 = ~N19;
  assign N23 = ~N22;
  assign N25 = ~N24;
  assign N28 = ~N27;

endmodule



module icache_eaddr_width_p64_data_width_p64_inst_width_p32_tag_width_p10_num_cce_p1_num_lce_p2_ways_p8_lce_sets_p64_block_size_in_bytes_p8
(
  clk_i,
  reset_i,
  id_i,
  pc_gen_icache_vaddr_i,
  pc_gen_icache_vaddr_v_i,
  pc_gen_icache_vaddr_ready_o,
  icache_pc_gen_data_o,
  icache_pc_gen_data_v_o,
  icache_pc_gen_data_ready_i,
  itlb_icache_data_resp_i,
  itlb_icache_data_resp_v_i,
  itlb_icache_data_resp_ready_o,
  cache_miss_o,
  poison_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  lce_tr_resp_i,
  lce_tr_resp_v_i,
  lce_tr_resp_ready_o,
  lce_tr_resp_o,
  lce_tr_resp_v_o,
  lce_tr_resp_ready_i
);

  input [0:0] id_i;
  input [63:0] pc_gen_icache_vaddr_i;
  output [95:0] icache_pc_gen_data_o;
  input [9:0] itlb_icache_data_resp_i;
  output [29:0] lce_req_o;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  input [35:0] lce_cmd_i;
  input [539:0] lce_data_cmd_i;
  input [538:0] lce_tr_resp_i;
  output [538:0] lce_tr_resp_o;
  input clk_i;
  input reset_i;
  input pc_gen_icache_vaddr_v_i;
  input icache_pc_gen_data_ready_i;
  input itlb_icache_data_resp_v_i;
  input poison_i;
  input lce_req_ready_i;
  input lce_resp_ready_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_v_i;
  input lce_tr_resp_v_i;
  input lce_tr_resp_ready_i;
  output pc_gen_icache_vaddr_ready_o;
  output icache_pc_gen_data_v_o;
  output itlb_icache_data_resp_ready_o;
  output cache_miss_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_ready_o;
  output lce_data_cmd_ready_o;
  output lce_tr_resp_ready_o;
  output lce_tr_resp_v_o;
  wire [29:0] lce_req_o;
  wire [25:0] lce_resp_o;
  wire [536:0] lce_data_resp_o;
  wire [538:0] lce_tr_resp_o;
  wire pc_gen_icache_vaddr_ready_o,icache_pc_gen_data_v_o,cache_miss_o,lce_req_v_o,
  lce_resp_v_o,lce_data_resp_v_o,lce_cmd_ready_o,lce_data_cmd_ready_o,
  lce_tr_resp_ready_o,lce_tr_resp_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  N17,N18,tl_we,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,
  N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,
  N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,
  N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,n_0_net_,tag_mem_w_li,tag_mem_v_li,
  n_1_net_,n_2_net_,n_3_net_,n_4_net_,n_5_net_,n_6_net_,n_7_net_,n_8_net_,tv_we,
  N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,
  N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,
  N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,
  N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,
  N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,
  N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,
  N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,
  N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,
  N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,
  N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,
  N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,
  N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,
  N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,
  N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,
  N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,
  N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,
  N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,
  N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,
  N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,
  N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,
  N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,
  N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,
  N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,
  N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,
  N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,
  N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,
  N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,
  N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,
  N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,
  N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,
  N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,
  N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,
  N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,
  N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,
  N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,
  N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,
  N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,
  N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,
  N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
  N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,
  N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,
  N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,
  N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,
  N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,
  N794,N795,N796,N797,N798,hit,miss_v,n_9_net_,metadata_mem_w_li,metadata_mem_v_li,
  n_10_net__7_,n_10_net__6_,n_10_net__5_,n_10_net__4_,n_10_net__3_,n_10_net__2_,
  n_10_net__1_,n_10_net__0_,invalid_exist,N799,data_mem_pkt_v_lo,
  data_mem_pkt_yumi_li,tag_mem_pkt_v_lo,tag_mem_pkt_yumi_li,metadata_mem_pkt_v_lo,
  metadata_mem_pkt_yumi_li,n_11_net__2_,n_11_net__1_,n_11_net__0_,N800,N801,N802,N803,n_15_net__0_,
  N804,n_17_net__1_,N805,N806,n_19_net__1_,n_19_net__0_,N807,n_21_net__2_,N808,N809,
  n_23_net__2_,n_23_net__0_,N810,N811,n_25_net__2_,n_25_net__1_,N812,N813,N814,
  n_27_net__2_,n_27_net__1_,n_27_net__0_,N815,N816,N817,N818,N819,N820,N821,N822,
  N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,N838,
  N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,N854,
  N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,N870,
  N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,N886,
  N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,N902,
  N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,N918,
  N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,N934,
  N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,N950,
  N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,N966,
  N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,N982,
  N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,N998,
  N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012,
  N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,N1025,
  N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038,
  N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,
  N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  n_29_net__0_,n_30_net__1_,n_31_net__1_,n_31_net__0_,n_32_net__2_,n_33_net__2_,
  n_33_net__0_,n_34_net__2_,n_34_net__1_,n_35_net__2_,n_35_net__1_,n_35_net__0_,N1065,N1066,
  N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079,
  N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091,N1092,
  N1093,N1094,N1095,N1096,N1097,N1098,N1099;
  wire [95:0] tag_mem_data_li,tag_mem_w_mask_li,tag_mem_data_lo;
  wire [5:0] tag_mem_addr_li,metadata_mem_addr_li;
  wire [71:0] data_mem_bank_addr_li;
  wire [7:0] data_mem_bank_w_li,data_mem_bank_v_li,hit_v;
  wire [511:0] data_mem_bank_data_lo,data_mem_data_li,data_mem_write_data;
  wire [2:0] hit_index,lru_encode,way_invalid_index,lru_way_li,lru_decode_way_li;
  wire [6:0] metadata_mem_data_li,metadata_mem_mask_li,metadata_mem_data_lo,
  lru_decode_data_lo,lru_decode_mask_lo;
  wire [521:0] data_mem_pkt;
  wire [22:0] tag_mem_pkt;
  wire [9:0] metadata_mem_pkt;
  wire [63:0] ld_data_way_picked;
  reg [63:0] eaddr_tl_r;
  reg itlb_icache_data_resp_ready_o,v_tv_r;
  reg [11:0] vaddr_tl_r;
  reg [511:0] ld_data_tv_r;
  reg [21:0] addr_tv_r;
  reg [95:0] icache_pc_gen_data_o;
  reg [79:0] tag_tv_r;
  reg [15:0] state_tv_r;
  reg [2:0] data_mem_pkt_way_r;

  bsg_mem_1rw_sync_mask_write_bit_width_p96_els_p64
  tag_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(tag_mem_data_li),
    .addr_i(tag_mem_addr_li),
    .v_i(n_0_net_),
    .w_mask_i(tag_mem_w_mask_li),
    .w_i(tag_mem_w_li),
    .data_o(tag_mem_data_lo)
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_banks_0__data_mem_bank
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_1_net_),
    .w_i(data_mem_bank_w_li[0]),
    .addr_i(data_mem_bank_addr_li[8:0]),
    .data_i(data_mem_write_data[63:0]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_bank_data_lo[63:0])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_banks_1__data_mem_bank
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_2_net_),
    .w_i(data_mem_bank_w_li[1]),
    .addr_i(data_mem_bank_addr_li[17:9]),
    .data_i(data_mem_write_data[127:64]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_bank_data_lo[127:64])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_banks_2__data_mem_bank
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_3_net_),
    .w_i(data_mem_bank_w_li[2]),
    .addr_i(data_mem_bank_addr_li[26:18]),
    .data_i(data_mem_write_data[191:128]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_bank_data_lo[191:128])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_banks_3__data_mem_bank
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_4_net_),
    .w_i(data_mem_bank_w_li[3]),
    .addr_i(data_mem_bank_addr_li[35:27]),
    .data_i(data_mem_write_data[255:192]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_bank_data_lo[255:192])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_banks_4__data_mem_bank
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_5_net_),
    .w_i(data_mem_bank_w_li[4]),
    .addr_i(data_mem_bank_addr_li[44:36]),
    .data_i(data_mem_write_data[319:256]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_bank_data_lo[319:256])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_banks_5__data_mem_bank
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_6_net_),
    .w_i(data_mem_bank_w_li[5]),
    .addr_i(data_mem_bank_addr_li[53:45]),
    .data_i(data_mem_write_data[383:320]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_bank_data_lo[383:320])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_banks_6__data_mem_bank
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_7_net_),
    .w_i(data_mem_bank_w_li[6]),
    .addr_i(data_mem_bank_addr_li[62:54]),
    .data_i(data_mem_write_data[447:384]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_bank_data_lo[447:384])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_banks_7__data_mem_bank
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_8_net_),
    .w_i(data_mem_bank_w_li[7]),
    .addr_i(data_mem_bank_addr_li[71:63]),
    .data_i(data_mem_write_data[511:448]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_bank_data_lo[511:448])
  );

  assign N791 = tag_tv_r[9:0] == addr_tv_r[21:12];
  assign N792 = tag_tv_r[19:10] == addr_tv_r[21:12];
  assign N793 = tag_tv_r[29:20] == addr_tv_r[21:12];
  assign N794 = tag_tv_r[39:30] == addr_tv_r[21:12];
  assign N795 = tag_tv_r[49:40] == addr_tv_r[21:12];
  assign N796 = tag_tv_r[59:50] == addr_tv_r[21:12];
  assign N797 = tag_tv_r[69:60] == addr_tv_r[21:12];
  assign N798 = tag_tv_r[79:70] == addr_tv_r[21:12];

  bsg_priority_encode_width_p8_lo_to_hi_p1
  pe_load_hit
  (
    .i(hit_v),
    .addr_o(hit_index),
    .v_o(hit)
  );


  bsg_mem_1rw_sync_mask_write_bit_width_p7_els_p64
  metadata_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(metadata_mem_data_li),
    .addr_i(metadata_mem_addr_li),
    .v_i(n_9_net_),
    .w_mask_i(metadata_mem_mask_li),
    .w_i(metadata_mem_w_li),
    .data_o(metadata_mem_data_lo)
  );


  bp_be_dcache_lru_encode_ways_p8
  lru_encoder
  (
    .lru_i(metadata_mem_data_lo),
    .way_id_o(lru_encode)
  );


  bsg_priority_encode_width_p8_lo_to_hi_p1
  pe_invalid
  (
    .i({ n_10_net__7_, n_10_net__6_, n_10_net__5_, n_10_net__4_, n_10_net__3_, n_10_net__2_, n_10_net__1_, n_10_net__0_ }),
    .addr_o(way_invalid_index),
    .v_o(invalid_exist)
  );


  bp_fe_sub_module1
  lce
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .id_i(id_i[0]),
    .ready_o(pc_gen_icache_vaddr_ready_o),
    .cache_miss_o(cache_miss_o),
    .miss_i(miss_v),
    .miss_addr_i(addr_tv_r),
    .data_mem_data_i(data_mem_data_li),
    .data_mem_pkt_o(data_mem_pkt),
    .data_mem_pkt_v_o(data_mem_pkt_v_lo),
    .data_mem_pkt_yumi_i(data_mem_pkt_yumi_li),
    .tag_mem_pkt_o(tag_mem_pkt),
    .tag_mem_pkt_v_o(tag_mem_pkt_v_lo),
    .tag_mem_pkt_yumi_i(tag_mem_pkt_yumi_li),
    .metadata_mem_pkt_v_o(metadata_mem_pkt_v_lo),
    .metadata_mem_pkt_o(metadata_mem_pkt),
    .lru_way_i(lru_way_li),
    .metadata_mem_pkt_yumi_i(metadata_mem_pkt_yumi_li),
    .lce_req_o(lce_req_o),
    .lce_req_v_o(lce_req_v_o),
    .lce_req_ready_i(lce_req_ready_i),
    .lce_resp_o(lce_resp_o),
    .lce_resp_v_o(lce_resp_v_o),
    .lce_resp_ready_i(lce_resp_ready_i),
    .lce_data_resp_o(lce_data_resp_o),
    .lce_data_resp_v_o(lce_data_resp_v_o),
    .lce_data_resp_ready_i(lce_data_resp_ready_i),
    .lce_cmd_i(lce_cmd_i),
    .lce_cmd_v_i(lce_cmd_v_i),
    .lce_cmd_ready_o(lce_cmd_ready_o),
    .lce_data_cmd_i(lce_data_cmd_i),
    .lce_data_cmd_v_i(lce_data_cmd_v_i),
    .lce_data_cmd_ready_o(lce_data_cmd_ready_o),
    .lce_tr_resp_i(lce_tr_resp_i),
    .lce_tr_resp_v_i(lce_tr_resp_v_i),
    .lce_tr_resp_ready_o(lce_tr_resp_ready_o),
    .lce_tr_resp_o(lce_tr_resp_o),
    .lce_tr_resp_v_o(lce_tr_resp_v_o),
    .lce_tr_resp_ready_i(lce_tr_resp_ready_i)
  );


  bsg_mux_width_p64_els_p8
  data_set_select_mux
  (
    .data_i(ld_data_tv_r),
    .sel_i({ n_11_net__2_, n_11_net__1_, n_11_net__0_ }),
    .data_o(ld_data_way_picked)
  );


  bsg_mux_width_p64_els_p8
  genblk4_0__data_mem_write_mux
  (
    .data_i(data_mem_pkt[511:0]),
    .sel_i(data_mem_pkt[515:513]),
    .data_o(data_mem_write_data[63:0])
  );


  bsg_mux_width_p64_els_p8
  genblk4_1__data_mem_write_mux
  (
    .data_i(data_mem_pkt[511:0]),
    .sel_i({ data_mem_pkt[515:514], n_15_net__0_ }),
    .data_o(data_mem_write_data[127:64])
  );


  bsg_mux_width_p64_els_p8
  genblk4_2__data_mem_write_mux
  (
    .data_i(data_mem_pkt[511:0]),
    .sel_i({ data_mem_pkt[515:515], n_17_net__1_, data_mem_pkt[513:513] }),
    .data_o(data_mem_write_data[191:128])
  );


  bsg_mux_width_p64_els_p8
  genblk4_3__data_mem_write_mux
  (
    .data_i(data_mem_pkt[511:0]),
    .sel_i({ data_mem_pkt[515:515], n_19_net__1_, n_19_net__0_ }),
    .data_o(data_mem_write_data[255:192])
  );


  bsg_mux_width_p64_els_p8
  genblk4_4__data_mem_write_mux
  (
    .data_i(data_mem_pkt[511:0]),
    .sel_i({ n_21_net__2_, data_mem_pkt[514:513] }),
    .data_o(data_mem_write_data[319:256])
  );


  bsg_mux_width_p64_els_p8
  genblk4_5__data_mem_write_mux
  (
    .data_i(data_mem_pkt[511:0]),
    .sel_i({ n_23_net__2_, data_mem_pkt[514:514], n_23_net__0_ }),
    .data_o(data_mem_write_data[383:320])
  );


  bsg_mux_width_p64_els_p8
  genblk4_6__data_mem_write_mux
  (
    .data_i(data_mem_pkt[511:0]),
    .sel_i({ n_25_net__2_, n_25_net__1_, data_mem_pkt[513:513] }),
    .data_o(data_mem_write_data[447:384])
  );


  bsg_mux_width_p64_els_p8
  genblk4_7__data_mem_write_mux
  (
    .data_i(data_mem_pkt[511:0]),
    .sel_i({ n_27_net__2_, n_27_net__1_, n_27_net__0_ }),
    .data_o(data_mem_write_data[511:448])
  );

  assign N817 = N815 & N816;
  assign N818 = tag_mem_pkt[1] | N816;
  assign N820 = N815 | tag_mem_pkt[0];
  assign N822 = tag_mem_pkt[1] & tag_mem_pkt[0];
  assign { N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } << { N837, N836, N835, N834, N833, N832, N831, N830 };
  assign { N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } << { N940, N939, N938, N937, N936, N935, N934 };

  bp_be_dcache_lru_decode_ways_p8
  lru_decode
  (
    .way_id_i(lru_decode_way_li),
    .data_o(lru_decode_data_lo),
    .mask_o(lru_decode_mask_lo)
  );


  bsg_mux_width_p64_els_p8
  genblk5_0__lce_data_mem_read_mux
  (
    .data_i(data_mem_bank_data_lo),
    .sel_i(data_mem_pkt_way_r),
    .data_o(data_mem_data_li[63:0])
  );


  bsg_mux_width_p64_els_p8
  genblk5_1__lce_data_mem_read_mux
  (
    .data_i(data_mem_bank_data_lo),
    .sel_i({ data_mem_pkt_way_r[2:1], n_29_net__0_ }),
    .data_o(data_mem_data_li[127:64])
  );


  bsg_mux_width_p64_els_p8
  genblk5_2__lce_data_mem_read_mux
  (
    .data_i(data_mem_bank_data_lo),
    .sel_i({ data_mem_pkt_way_r[2:2], n_30_net__1_, data_mem_pkt_way_r[0:0] }),
    .data_o(data_mem_data_li[191:128])
  );


  bsg_mux_width_p64_els_p8
  genblk5_3__lce_data_mem_read_mux
  (
    .data_i(data_mem_bank_data_lo),
    .sel_i({ data_mem_pkt_way_r[2:2], n_31_net__1_, n_31_net__0_ }),
    .data_o(data_mem_data_li[255:192])
  );


  bsg_mux_width_p64_els_p8
  genblk5_4__lce_data_mem_read_mux
  (
    .data_i(data_mem_bank_data_lo),
    .sel_i({ n_32_net__2_, data_mem_pkt_way_r[1:0] }),
    .data_o(data_mem_data_li[319:256])
  );


  bsg_mux_width_p64_els_p8
  genblk5_5__lce_data_mem_read_mux
  (
    .data_i(data_mem_bank_data_lo),
    .sel_i({ n_33_net__2_, data_mem_pkt_way_r[1:1], n_33_net__0_ }),
    .data_o(data_mem_data_li[383:320])
  );


  bsg_mux_width_p64_els_p8
  genblk5_6__lce_data_mem_read_mux
  (
    .data_i(data_mem_bank_data_lo),
    .sel_i({ n_34_net__2_, n_34_net__1_, data_mem_pkt_way_r[0:0] }),
    .data_o(data_mem_data_li[447:384])
  );


  bsg_mux_width_p64_els_p8
  genblk5_7__lce_data_mem_read_mux
  (
    .data_i(data_mem_bank_data_lo),
    .sel_i({ n_35_net__2_, n_35_net__1_, n_35_net__0_ }),
    .data_o(data_mem_data_li[511:448])
  );

  assign N1065 = state_tv_r[14] | state_tv_r[15];
  assign N1066 = state_tv_r[12] | state_tv_r[13];
  assign N1067 = state_tv_r[10] | state_tv_r[11];
  assign N1068 = state_tv_r[8] | state_tv_r[9];
  assign N1069 = state_tv_r[6] | state_tv_r[7];
  assign N1070 = state_tv_r[4] | state_tv_r[5];
  assign N1071 = state_tv_r[2] | state_tv_r[3];
  assign N1072 = state_tv_r[0] | state_tv_r[1];
  assign N1073 = state_tv_r[14] | state_tv_r[15];
  assign N1074 = state_tv_r[12] | state_tv_r[13];
  assign N1075 = state_tv_r[10] | state_tv_r[11];
  assign N1076 = state_tv_r[8] | state_tv_r[9];
  assign N1077 = state_tv_r[6] | state_tv_r[7];
  assign N1078 = state_tv_r[4] | state_tv_r[5];
  assign N1079 = state_tv_r[2] | state_tv_r[3];
  assign N1080 = state_tv_r[0] | state_tv_r[1];
  assign { N940, N939, N938, N937, N936, N935, N934 } = tag_mem_pkt[16:14] * { 1'b1, 1'b1, 1'b0, 1'b0 };
  assign { N829, N828, N827, N826, N825, N824, N823 } = tag_mem_pkt[16:14] * { 1'b1, 1'b1, 1'b0, 1'b0 };
  assign { N837, N836, N835, N834, N833, N832, N831, N830 } = { N829, N828, N827, N826, N825, N824, N823 } + { 1'b1, 1'b0, 1'b1, 1'b0 };
  assign N21 = (N0)? 1'b0 : 
               (N1)? tl_we : 1'b0;
  assign N0 = N20;
  assign N1 = N19;
  assign N22 = (N0)? 1'b1 : 
               (N1)? tl_we : 1'b0;
  assign { N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                          (N1)? pc_gen_icache_vaddr_i[11:0] : 1'b0;
  assign { N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                  (N1)? pc_gen_icache_vaddr_i[63:12] : 1'b0;
  assign N89 = (N2)? 1'b0 : 
               (N3)? tv_we : 1'b0;
  assign N2 = N88;
  assign N3 = N87;
  assign { N102, N100, N98, N96, N94, N92, N90 } = (N2)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                   (N3)? { tv_we, tv_we, tv_we, tv_we, tv_we, tv_we, tv_we } : 1'b0;
  assign { N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N101, N99, N97, N95, N93, N91 } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                             (N3)? { itlb_icache_data_resp_i, vaddr_tl_r } : 1'b0;
  assign { N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119 } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N3)? eaddr_tl_r : 1'b0;
  assign { N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183 } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3)? { tag_mem_data_lo[93:84], tag_mem_data_lo[81:72], tag_mem_data_lo[69:60], tag_mem_data_lo[57:48], tag_mem_data_lo[45:36], tag_mem_data_lo[33:24], tag_mem_data_lo[21:12], tag_mem_data_lo[9:0] } : 1'b0;
  assign { N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263 } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                              (N3)? { tag_mem_data_lo[95:94], tag_mem_data_lo[83:82], tag_mem_data_lo[71:70], tag_mem_data_lo[59:58], tag_mem_data_lo[47:46], tag_mem_data_lo[35:34], tag_mem_data_lo[23:22], tag_mem_data_lo[11:10] } : 1'b0;
  assign { N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279 } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3)? data_mem_bank_data_lo : 1'b0;
  assign lru_way_li = (N4)? way_invalid_index : 
                      (N5)? lru_encode : 1'b0;
  assign N4 = invalid_exist;
  assign N5 = N799;
  assign icache_pc_gen_data_o[95:64] = (N6)? ld_data_way_picked[63:32] : 
                                       (N7)? ld_data_way_picked[31:0] : 1'b0;
  assign N6 = N801;
  assign N7 = N800;
  assign data_mem_bank_v_li = (N8)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                              (N9)? { data_mem_pkt_yumi_li, data_mem_pkt_yumi_li, data_mem_pkt_yumi_li, data_mem_pkt_yumi_li, data_mem_pkt_yumi_li, data_mem_pkt_yumi_li, data_mem_pkt_yumi_li, data_mem_pkt_yumi_li } : 1'b0;
  assign N8 = tl_we;
  assign N9 = N802;
  assign data_mem_bank_addr_li[8:0] = (N8)? pc_gen_icache_vaddr_i[11:3] : 
                                      (N9)? data_mem_pkt[521:513] : 1'b0;
  assign data_mem_bank_addr_li[17:9] = (N8)? pc_gen_icache_vaddr_i[11:3] : 
                                       (N9)? { data_mem_pkt[521:514], N803 } : 1'b0;
  assign data_mem_bank_addr_li[26:18] = (N8)? pc_gen_icache_vaddr_i[11:3] : 
                                        (N9)? { data_mem_pkt[521:515], N804, data_mem_pkt[513:513] } : 1'b0;
  assign data_mem_bank_addr_li[35:27] = (N8)? pc_gen_icache_vaddr_i[11:3] : 
                                        (N9)? { data_mem_pkt[521:515], N805, N806 } : 1'b0;
  assign data_mem_bank_addr_li[44:36] = (N8)? pc_gen_icache_vaddr_i[11:3] : 
                                        (N9)? { data_mem_pkt[521:516], N807, data_mem_pkt[514:513] } : 1'b0;
  assign data_mem_bank_addr_li[53:45] = (N8)? pc_gen_icache_vaddr_i[11:3] : 
                                        (N9)? { data_mem_pkt[521:516], N808, data_mem_pkt[514:514], N809 } : 1'b0;
  assign data_mem_bank_addr_li[62:54] = (N8)? pc_gen_icache_vaddr_i[11:3] : 
                                        (N9)? { data_mem_pkt[521:516], N810, N811, data_mem_pkt[513:513] } : 1'b0;
  assign data_mem_bank_addr_li[71:63] = (N8)? pc_gen_icache_vaddr_i[11:3] : 
                                        (N9)? { data_mem_pkt[521:516], N812, N813, N814 } : 1'b0;
  assign tag_mem_addr_li = (N8)? pc_gen_icache_vaddr_i[11:6] : 
                           (N9)? tag_mem_pkt[22:17] : 1'b0;
  assign tag_mem_data_li = (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N12)? { tag_mem_pkt[13:2], tag_mem_pkt[13:2], tag_mem_pkt[13:2], tag_mem_pkt[13:2], tag_mem_pkt[13:2], tag_mem_pkt[13:2], tag_mem_pkt[13:2], tag_mem_pkt[13:2] } : 
                           (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = N817;
  assign N11 = N819;
  assign N12 = N821;
  assign N13 = N822;
  assign tag_mem_w_mask_li = (N10)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                             (N11)? { N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838 } : 
                             (N12)? { N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941 } : 
                             (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign metadata_mem_addr_li = (N14)? addr_tv_r[11:6] : 
                                (N15)? metadata_mem_pkt[9:4] : 1'b0;
  assign N14 = v_tv_r;
  assign N15 = N1037;
  assign { N1052, N1051, N1050, N1049, N1048, N1047, N1046 } = (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N17)? { N1039, N1040, N1041, N1042, N1043, N1044, N1045 } : 1'b0;
  assign N16 = N1038;
  assign N17 = metadata_mem_pkt[0];
  assign { N1059, N1058, N1057, N1056, N1055, N1054, N1053 } = (N16)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                               (N17)? lru_decode_mask_lo : 1'b0;
  assign lru_decode_way_li = (N14)? hit_index : 
                             (N15)? metadata_mem_pkt[3:1] : 1'b0;
  assign metadata_mem_data_li = (N14)? lru_decode_data_lo : 
                                (N15)? { N1052, N1051, N1050, N1049, N1048, N1047, N1046 } : 1'b0;
  assign metadata_mem_mask_li = (N14)? lru_decode_mask_lo : 
                                (N15)? { N1059, N1058, N1057, N1056, N1055, N1054, N1053 } : 1'b0;
  assign { N1064, N1063, N1062 } = (N18)? data_mem_pkt[515:513] : 
                                   (N1061)? data_mem_pkt_way_r : 1'b0;
  assign N18 = N1060;
  assign tl_we = N1081 & N1082;
  assign N1081 = pc_gen_icache_vaddr_v_i & pc_gen_icache_vaddr_ready_o;
  assign N1082 = ~poison_i;
  assign N19 = ~reset_i;
  assign N20 = reset_i;
  assign n_0_net_ = N1083 & tag_mem_v_li;
  assign N1083 = ~reset_i;
  assign n_1_net_ = N1084 & data_mem_bank_v_li[0];
  assign N1084 = ~reset_i;
  assign n_2_net_ = N1085 & data_mem_bank_v_li[1];
  assign N1085 = ~reset_i;
  assign n_3_net_ = N1086 & data_mem_bank_v_li[2];
  assign N1086 = ~reset_i;
  assign n_4_net_ = N1087 & data_mem_bank_v_li[3];
  assign N1087 = ~reset_i;
  assign n_5_net_ = N1088 & data_mem_bank_v_li[4];
  assign N1088 = ~reset_i;
  assign n_6_net_ = N1089 & data_mem_bank_v_li[5];
  assign N1089 = ~reset_i;
  assign n_7_net_ = N1090 & data_mem_bank_v_li[6];
  assign N1090 = ~reset_i;
  assign n_8_net_ = N1091 & data_mem_bank_v_li[7];
  assign N1091 = ~reset_i;
  assign tv_we = N1092 & itlb_icache_data_resp_v_i;
  assign N1092 = itlb_icache_data_resp_ready_o & N1082;
  assign N87 = ~reset_i;
  assign N88 = reset_i;
  assign hit_v[0] = N791 & N1072;
  assign hit_v[1] = N792 & N1071;
  assign hit_v[2] = N793 & N1070;
  assign hit_v[3] = N794 & N1069;
  assign hit_v[4] = N795 & N1068;
  assign hit_v[5] = N796 & N1067;
  assign hit_v[6] = N797 & N1066;
  assign hit_v[7] = N798 & N1065;
  assign miss_v = N1093 & v_tv_r;
  assign N1093 = ~hit;
  assign n_9_net_ = N1094 & metadata_mem_v_li;
  assign N1094 = ~reset_i;
  assign n_10_net__7_ = ~N1073;
  assign n_10_net__6_ = ~N1074;
  assign n_10_net__5_ = ~N1075;
  assign n_10_net__4_ = ~N1076;
  assign n_10_net__3_ = ~N1077;
  assign n_10_net__2_ = ~N1078;
  assign n_10_net__1_ = ~N1079;
  assign n_10_net__0_ = ~N1080;
  assign N799 = ~invalid_exist;
  assign icache_pc_gen_data_v_o = N1096 & N1097;
  assign N1096 = v_tv_r & N1095;
  assign N1095 = ~miss_v;
  assign N1097 = ~reset_i;
  assign n_11_net__2_ = hit_index[2] ^ addr_tv_r[5];
  assign n_11_net__1_ = hit_index[1] ^ addr_tv_r[4];
  assign n_11_net__0_ = hit_index[0] ^ addr_tv_r[3];
  assign N800 = ~addr_tv_r[2];
  assign N801 = addr_tv_r[2];
  assign N802 = ~tl_we;
  assign data_mem_bank_w_li[7] = data_mem_pkt_yumi_li & data_mem_pkt[512];
  assign data_mem_bank_w_li[6] = data_mem_pkt_yumi_li & data_mem_pkt[512];
  assign data_mem_bank_w_li[5] = data_mem_pkt_yumi_li & data_mem_pkt[512];
  assign data_mem_bank_w_li[4] = data_mem_pkt_yumi_li & data_mem_pkt[512];
  assign data_mem_bank_w_li[3] = data_mem_pkt_yumi_li & data_mem_pkt[512];
  assign data_mem_bank_w_li[2] = data_mem_pkt_yumi_li & data_mem_pkt[512];
  assign data_mem_bank_w_li[1] = data_mem_pkt_yumi_li & data_mem_pkt[512];
  assign data_mem_bank_w_li[0] = data_mem_pkt_yumi_li & data_mem_pkt[512];
  assign N803 = ~data_mem_pkt[513];
  assign n_15_net__0_ = ~data_mem_pkt[513];
  assign N804 = ~data_mem_pkt[514];
  assign n_17_net__1_ = ~data_mem_pkt[514];
  assign N805 = ~data_mem_pkt[514];
  assign N806 = ~data_mem_pkt[513];
  assign n_19_net__1_ = ~data_mem_pkt[514];
  assign n_19_net__0_ = ~data_mem_pkt[513];
  assign N807 = ~data_mem_pkt[515];
  assign n_21_net__2_ = ~data_mem_pkt[515];
  assign N808 = ~data_mem_pkt[515];
  assign N809 = ~data_mem_pkt[513];
  assign n_23_net__2_ = ~data_mem_pkt[515];
  assign n_23_net__0_ = ~data_mem_pkt[513];
  assign N810 = ~data_mem_pkt[515];
  assign N811 = ~data_mem_pkt[514];
  assign n_25_net__2_ = ~data_mem_pkt[515];
  assign n_25_net__1_ = ~data_mem_pkt[514];
  assign N812 = ~data_mem_pkt[515];
  assign N813 = ~data_mem_pkt[514];
  assign N814 = ~data_mem_pkt[513];
  assign n_27_net__2_ = ~data_mem_pkt[515];
  assign n_27_net__1_ = ~data_mem_pkt[514];
  assign n_27_net__0_ = ~data_mem_pkt[513];
  assign tag_mem_v_li = tl_we | tag_mem_pkt_yumi_li;
  assign tag_mem_w_li = N802 & tag_mem_pkt_v_lo;
  assign N815 = ~tag_mem_pkt[1];
  assign N816 = ~tag_mem_pkt[0];
  assign N819 = ~N818;
  assign N821 = ~N820;
  assign metadata_mem_v_li = v_tv_r | metadata_mem_pkt_yumi_li;
  assign metadata_mem_w_li = N1099 | metadata_mem_pkt_yumi_li;
  assign N1099 = v_tv_r & N1098;
  assign N1098 = ~miss_v;
  assign N1037 = ~v_tv_r;
  assign N1038 = ~metadata_mem_pkt[0];
  assign N1039 = ~lru_decode_data_lo[6];
  assign N1040 = ~lru_decode_data_lo[5];
  assign N1041 = ~lru_decode_data_lo[4];
  assign N1042 = ~lru_decode_data_lo[3];
  assign N1043 = ~lru_decode_data_lo[2];
  assign N1044 = ~lru_decode_data_lo[1];
  assign N1045 = ~lru_decode_data_lo[0];
  assign N1060 = data_mem_pkt_v_lo & data_mem_pkt_yumi_li;
  assign N1061 = ~N1060;
  assign n_29_net__0_ = ~data_mem_pkt_way_r[0];
  assign n_30_net__1_ = ~data_mem_pkt_way_r[1];
  assign n_31_net__1_ = ~data_mem_pkt_way_r[1];
  assign n_31_net__0_ = ~data_mem_pkt_way_r[0];
  assign n_32_net__2_ = ~data_mem_pkt_way_r[2];
  assign n_33_net__2_ = ~data_mem_pkt_way_r[2];
  assign n_33_net__0_ = ~data_mem_pkt_way_r[0];
  assign n_34_net__2_ = ~data_mem_pkt_way_r[2];
  assign n_34_net__1_ = ~data_mem_pkt_way_r[1];
  assign n_35_net__2_ = ~data_mem_pkt_way_r[2];
  assign n_35_net__1_ = ~data_mem_pkt_way_r[1];
  assign n_35_net__0_ = ~data_mem_pkt_way_r[0];
  assign data_mem_pkt_yumi_li = data_mem_pkt_v_lo & N802;
  assign tag_mem_pkt_yumi_li = tag_mem_pkt_v_lo & N802;
  assign metadata_mem_pkt_yumi_li = N1037 & metadata_mem_pkt_v_lo;

  always @(posedge clk_i) begin
    if(N22) begin
      { eaddr_tl_r[63:0] } <= { N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23 };
      { vaddr_tl_r[11:0] } <= { N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23 };
    end 
    if(1'b1) begin
      itlb_icache_data_resp_ready_o <= N21;
      v_tv_r <= N89;
      { data_mem_pkt_way_r[2:0] } <= { N1064, N1063, N1062 };
    end 
    if(N90) begin
      { ld_data_tv_r[511:413] } <= { N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692 };
      { addr_tv_r[0:0] } <= { N91 };
    end 
    if(N92) begin
      { ld_data_tv_r[412:314] } <= { N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593 };
      { addr_tv_r[1:1] } <= { N93 };
    end 
    if(N94) begin
      { ld_data_tv_r[313:215] } <= { N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494 };
      { addr_tv_r[2:2] } <= { N95 };
    end 
    if(N96) begin
      { ld_data_tv_r[214:116] } <= { N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395 };
      { addr_tv_r[3:3] } <= { N97 };
    end 
    if(N98) begin
      { ld_data_tv_r[115:17] } <= { N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296 };
      { addr_tv_r[4:4] } <= { N99 };
    end 
    if(N100) begin
      { ld_data_tv_r[16:0] } <= { N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279 };
      { addr_tv_r[5:5] } <= { N101 };
      { tag_tv_r[79:14] } <= { N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197 };
      { state_tv_r[15:0] } <= { N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263 };
    end 
    if(N102) begin
      { addr_tv_r[21:6] } <= { N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103 };
      { icache_pc_gen_data_o[63:0] } <= { N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119 };
      { tag_tv_r[13:0] } <= { N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183 };
    end 
  end


endmodule



module itlb_vaddr_width_p56_paddr_width_p22_eaddr_width_p64_btb_indx_width_p9_bht_indx_width_p5_ras_addr_width_p22_asid_width_p10_ppn_start_bit_p12_tag_width_p10
(
  clk_i,
  reset_i,
  fe_itlb_i,
  fe_itlb_v_i,
  fe_itlb_ready_o,
  pc_gen_itlb_i,
  pc_gen_itlb_v_i,
  pc_gen_itlb_ready_o,
  itlb_icache_o,
  itlb_icache_data_resp_v_o,
  itlb_icache_data_resp_ready_i,
  itlb_fe_o,
  itlb_fe_v_o,
  itlb_fe_ready_i
);

  input [108:0] fe_itlb_i;
  input [63:0] pc_gen_itlb_i;
  output [9:0] itlb_icache_o;
  output [133:0] itlb_fe_o;
  input clk_i;
  input reset_i;
  input fe_itlb_v_i;
  input pc_gen_itlb_v_i;
  input itlb_icache_data_resp_ready_i;
  input itlb_fe_ready_i;
  output fe_itlb_ready_o;
  output pc_gen_itlb_ready_o;
  output itlb_icache_data_resp_v_o;
  output itlb_fe_v_o;
  wire [133:0] itlb_fe_o;
  wire fe_itlb_ready_o,pc_gen_itlb_ready_o,itlb_icache_data_resp_v_o,itlb_fe_v_o;
  reg [9:0] itlb_icache_o;
  assign pc_gen_itlb_ready_o = 1'b1;
  assign itlb_icache_data_resp_v_o = 1'b1;
  assign fe_itlb_ready_o = 1'b0;
  assign itlb_fe_v_o = 1'b0;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { itlb_icache_o[9:0] } <= { pc_gen_itlb_i[21:12] };
    end 
  end


endmodule



module bp_fe_top
(
  clk_i,
  reset_i,
  icache_id_i,
  bp_fe_cmd_i,
  bp_fe_cmd_v_i,
  bp_fe_cmd_ready_o,
  bp_fe_queue_o,
  bp_fe_queue_v_o,
  bp_fe_queue_ready_i,
  lce_cce_req_o,
  lce_cce_req_v_o,
  lce_cce_req_ready_i,
  lce_cce_resp_o,
  lce_cce_resp_v_o,
  lce_cce_resp_ready_i,
  lce_cce_data_resp_o,
  lce_cce_data_resp_v_o,
  lce_cce_data_resp_ready_i,
  cce_lce_cmd_i,
  cce_lce_cmd_v_i,
  cce_lce_cmd_ready_o,
  cce_lce_data_cmd_i,
  cce_lce_data_cmd_v_i,
  cce_lce_data_cmd_ready_o,
  lce_lce_tr_resp_i,
  lce_lce_tr_resp_v_i,
  lce_lce_tr_resp_ready_o,
  lce_lce_tr_resp_o,
  lce_lce_tr_resp_v_o,
  lce_lce_tr_resp_ready_i
);

  input [0:0] icache_id_i;
  input [108:0] bp_fe_cmd_i;
  output [133:0] bp_fe_queue_o;
  output [29:0] lce_cce_req_o;
  output [25:0] lce_cce_resp_o;
  output [536:0] lce_cce_data_resp_o;
  input [35:0] cce_lce_cmd_i;
  input [539:0] cce_lce_data_cmd_i;
  input [538:0] lce_lce_tr_resp_i;
  output [538:0] lce_lce_tr_resp_o;
  input clk_i;
  input reset_i;
  input bp_fe_cmd_v_i;
  input bp_fe_queue_ready_i;
  input lce_cce_req_ready_i;
  input lce_cce_resp_ready_i;
  input lce_cce_data_resp_ready_i;
  input cce_lce_cmd_v_i;
  input cce_lce_data_cmd_v_i;
  input lce_lce_tr_resp_v_i;
  input lce_lce_tr_resp_ready_i;
  output bp_fe_cmd_ready_o;
  output bp_fe_queue_v_o;
  output lce_cce_req_v_o;
  output lce_cce_resp_v_o;
  output lce_cce_data_resp_v_o;
  output cce_lce_cmd_ready_o;
  output cce_lce_data_cmd_ready_o;
  output lce_lce_tr_resp_ready_o;
  output lce_lce_tr_resp_v_o;
  wire [133:0] bp_fe_queue_o,itlb_fe_queue;
  wire [29:0] lce_cce_req_o;
  wire [25:0] lce_cce_resp_o;
  wire [536:0] lce_cce_data_resp_o;
  wire [538:0] lce_lce_tr_resp_o;
  wire bp_fe_cmd_ready_o,bp_fe_queue_v_o,lce_cce_req_v_o,lce_cce_resp_v_o,
  lce_cce_data_resp_v_o,cce_lce_cmd_ready_o,cce_lce_data_cmd_ready_o,lce_lce_tr_resp_ready_o,
  lce_lce_tr_resp_v_o,N0,N1,pc_gen_queue_scan_instr__68_,
  pc_gen_queue_scan_instr__67_,pc_gen_queue_scan_instr__66_,pc_gen_queue_scan_instr__65_,
  pc_gen_queue_scan_instr__64_,pc_gen_queue_scan_instr__63_,pc_gen_queue_scan_instr__62_,
  pc_gen_queue_scan_instr__61_,pc_gen_queue_scan_instr__60_,pc_gen_queue_scan_instr__59_,
  pc_gen_queue_scan_instr__58_,pc_gen_queue_scan_instr__57_,
  pc_gen_queue_scan_instr__56_,pc_gen_queue_scan_instr__55_,pc_gen_queue_scan_instr__54_,
  pc_gen_queue_scan_instr__53_,pc_gen_queue_scan_instr__52_,pc_gen_queue_scan_instr__51_,
  pc_gen_queue_scan_instr__50_,pc_gen_queue_scan_instr__49_,pc_gen_queue_scan_instr__48_,
  pc_gen_queue_scan_instr__47_,pc_gen_queue_scan_instr__46_,pc_gen_queue_scan_instr__45_,
  pc_gen_queue_scan_instr__44_,pc_gen_queue_scan_instr__43_,
  pc_gen_queue_scan_instr__42_,pc_gen_queue_scan_instr__41_,pc_gen_queue_scan_instr__40_,
  pc_gen_queue_scan_instr__39_,pc_gen_queue_scan_instr__38_,pc_gen_queue_scan_instr__37_,
  pc_gen_queue_scan_instr__36_,pc_gen_queue_scan_instr__35_,pc_gen_queue_scan_instr__34_,
  pc_gen_queue_scan_instr__33_,pc_gen_queue_scan_instr__32_,
  pc_gen_queue_scan_instr__31_,pc_gen_queue_scan_instr__30_,pc_gen_queue_scan_instr__29_,
  pc_gen_queue_scan_instr__28_,pc_gen_queue_scan_instr__27_,pc_gen_queue_scan_instr__26_,
  pc_gen_queue_scan_instr__25_,pc_gen_queue_scan_instr__24_,pc_gen_queue_scan_instr__23_,
  pc_gen_queue_scan_instr__22_,pc_gen_queue_scan_instr__21_,
  pc_gen_queue_scan_instr__20_,pc_gen_queue_scan_instr__19_,pc_gen_queue_scan_instr__18_,
  pc_gen_queue_scan_instr__17_,pc_gen_queue_scan_instr__16_,pc_gen_queue_scan_instr__15_,
  pc_gen_queue_scan_instr__14_,pc_gen_queue_scan_instr__13_,pc_gen_queue_scan_instr__12_,
  pc_gen_queue_scan_instr__11_,pc_gen_queue_scan_instr__10_,
  pc_gen_queue_scan_instr__9_,pc_gen_queue_scan_instr__8_,pc_gen_queue_scan_instr__7_,
  pc_gen_queue_scan_instr__6_,pc_gen_queue_scan_instr__5_,pc_gen_queue_scan_instr__4_,
  pc_gen_queue_scan_instr__3_,pc_gen_queue_scan_instr__2_,pc_gen_queue_scan_instr__1_,
  pc_gen_queue_scan_instr__0_,fe_pc_gen_branch_metadata_fwd__35_,
  fe_pc_gen_branch_metadata_fwd__34_,fe_pc_gen_branch_metadata_fwd__33_,fe_pc_gen_branch_metadata_fwd__32_,
  fe_pc_gen_branch_metadata_fwd__31_,fe_pc_gen_branch_metadata_fwd__30_,
  fe_pc_gen_branch_metadata_fwd__29_,fe_pc_gen_branch_metadata_fwd__28_,
  fe_pc_gen_branch_metadata_fwd__27_,fe_pc_gen_branch_metadata_fwd__26_,fe_pc_gen_branch_metadata_fwd__25_,
  fe_pc_gen_branch_metadata_fwd__24_,fe_pc_gen_branch_metadata_fwd__23_,
  fe_pc_gen_branch_metadata_fwd__22_,fe_pc_gen_branch_metadata_fwd__21_,
  fe_pc_gen_branch_metadata_fwd__20_,fe_pc_gen_branch_metadata_fwd__19_,
  fe_pc_gen_branch_metadata_fwd__18_,fe_pc_gen_branch_metadata_fwd__17_,fe_pc_gen_branch_metadata_fwd__16_,
  fe_pc_gen_branch_metadata_fwd__15_,fe_pc_gen_branch_metadata_fwd__14_,
  fe_pc_gen_branch_metadata_fwd__13_,fe_pc_gen_branch_metadata_fwd__12_,
  fe_pc_gen_branch_metadata_fwd__11_,fe_pc_gen_branch_metadata_fwd__10_,fe_pc_gen_branch_metadata_fwd__9_,
  fe_pc_gen_branch_metadata_fwd__8_,fe_pc_gen_branch_metadata_fwd__7_,
  fe_pc_gen_branch_metadata_fwd__6_,fe_pc_gen_branch_metadata_fwd__5_,
  fe_pc_gen_branch_metadata_fwd__4_,fe_pc_gen_branch_metadata_fwd__3_,fe_pc_gen_branch_metadata_fwd__2_,
  fe_pc_gen_branch_metadata_fwd__1_,fe_pc_gen_branch_metadata_fwd__0_,
  fe_pc_gen_pc_redirect_valid_,N2,N3,cache_miss,poison,pc_gen_icache_v,pc_gen_icache_ready,
  icache_pc_gen_v,icache_pc_gen_ready,pc_gen_itlb_v,pc_gen_itlb_ready,
  itlb_icache_data_resp_v,itlb_icache_data_resp_ready,fe_itlb_ready,itlb_fe_v,N4,N5,N6,N7,N8,N9,N10,
  N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28;
  wire [63:0] pc_gen_icache,pc_gen_itlb;
  wire [95:0] icache_pc_gen;
  wire [9:0] itlb_icache;

  bp_fe_pc_gen_56_22_64_9_5_22_32_10_80000124_1
  bp_fe_pc_gen_1
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(1'b1),
    .pc_gen_icache_o(pc_gen_icache),
    .pc_gen_icache_v_o(pc_gen_icache_v),
    .pc_gen_icache_ready_i(pc_gen_icache_ready),
    .icache_pc_gen_i(icache_pc_gen),
    .icache_pc_gen_v_i(icache_pc_gen_v),
    .icache_pc_gen_ready_o(icache_pc_gen_ready),
    .icache_miss_i(cache_miss),
    .pc_gen_itlb_o(pc_gen_itlb),
    .pc_gen_itlb_v_o(pc_gen_itlb_v),
    .pc_gen_itlb_ready_i(pc_gen_itlb_ready),
    .pc_gen_fe_o({ bp_fe_queue_o[133:133], pc_gen_queue_scan_instr__68_, pc_gen_queue_scan_instr__67_, pc_gen_queue_scan_instr__66_, pc_gen_queue_scan_instr__65_, pc_gen_queue_scan_instr__64_, pc_gen_queue_scan_instr__63_, pc_gen_queue_scan_instr__62_, pc_gen_queue_scan_instr__61_, pc_gen_queue_scan_instr__60_, pc_gen_queue_scan_instr__59_, pc_gen_queue_scan_instr__58_, pc_gen_queue_scan_instr__57_, pc_gen_queue_scan_instr__56_, pc_gen_queue_scan_instr__55_, pc_gen_queue_scan_instr__54_, pc_gen_queue_scan_instr__53_, pc_gen_queue_scan_instr__52_, pc_gen_queue_scan_instr__51_, pc_gen_queue_scan_instr__50_, pc_gen_queue_scan_instr__49_, pc_gen_queue_scan_instr__48_, pc_gen_queue_scan_instr__47_, pc_gen_queue_scan_instr__46_, pc_gen_queue_scan_instr__45_, pc_gen_queue_scan_instr__44_, pc_gen_queue_scan_instr__43_, pc_gen_queue_scan_instr__42_, pc_gen_queue_scan_instr__41_, pc_gen_queue_scan_instr__40_, pc_gen_queue_scan_instr__39_, pc_gen_queue_scan_instr__38_, pc_gen_queue_scan_instr__37_, pc_gen_queue_scan_instr__36_, pc_gen_queue_scan_instr__35_, pc_gen_queue_scan_instr__34_, pc_gen_queue_scan_instr__33_, pc_gen_queue_scan_instr__32_, pc_gen_queue_scan_instr__31_, pc_gen_queue_scan_instr__30_, pc_gen_queue_scan_instr__29_, pc_gen_queue_scan_instr__28_, pc_gen_queue_scan_instr__27_, pc_gen_queue_scan_instr__26_, pc_gen_queue_scan_instr__25_, pc_gen_queue_scan_instr__24_, pc_gen_queue_scan_instr__23_, pc_gen_queue_scan_instr__22_, pc_gen_queue_scan_instr__21_, pc_gen_queue_scan_instr__20_, pc_gen_queue_scan_instr__19_, pc_gen_queue_scan_instr__18_, pc_gen_queue_scan_instr__17_, pc_gen_queue_scan_instr__16_, pc_gen_queue_scan_instr__15_, pc_gen_queue_scan_instr__14_, pc_gen_queue_scan_instr__13_, pc_gen_queue_scan_instr__12_, pc_gen_queue_scan_instr__11_, pc_gen_queue_scan_instr__10_, pc_gen_queue_scan_instr__9_, pc_gen_queue_scan_instr__8_, pc_gen_queue_scan_instr__7_, pc_gen_queue_scan_instr__6_, pc_gen_queue_scan_instr__5_, pc_gen_queue_scan_instr__4_, pc_gen_queue_scan_instr__3_, pc_gen_queue_scan_instr__2_, pc_gen_queue_scan_instr__1_, pc_gen_queue_scan_instr__0_, bp_fe_queue_o[132:0] }),
    .pc_gen_fe_v_o(bp_fe_queue_v_o),
    .pc_gen_fe_ready_i(bp_fe_queue_ready_i),
    .fe_pc_gen_i({ bp_fe_cmd_i[105:42], fe_pc_gen_branch_metadata_fwd__35_, fe_pc_gen_branch_metadata_fwd__34_, fe_pc_gen_branch_metadata_fwd__33_, fe_pc_gen_branch_metadata_fwd__32_, fe_pc_gen_branch_metadata_fwd__31_, fe_pc_gen_branch_metadata_fwd__30_, fe_pc_gen_branch_metadata_fwd__29_, fe_pc_gen_branch_metadata_fwd__28_, fe_pc_gen_branch_metadata_fwd__27_, fe_pc_gen_branch_metadata_fwd__26_, fe_pc_gen_branch_metadata_fwd__25_, fe_pc_gen_branch_metadata_fwd__24_, fe_pc_gen_branch_metadata_fwd__23_, fe_pc_gen_branch_metadata_fwd__22_, fe_pc_gen_branch_metadata_fwd__21_, fe_pc_gen_branch_metadata_fwd__20_, fe_pc_gen_branch_metadata_fwd__19_, fe_pc_gen_branch_metadata_fwd__18_, fe_pc_gen_branch_metadata_fwd__17_, fe_pc_gen_branch_metadata_fwd__16_, fe_pc_gen_branch_metadata_fwd__15_, fe_pc_gen_branch_metadata_fwd__14_, fe_pc_gen_branch_metadata_fwd__13_, fe_pc_gen_branch_metadata_fwd__12_, fe_pc_gen_branch_metadata_fwd__11_, fe_pc_gen_branch_metadata_fwd__10_, fe_pc_gen_branch_metadata_fwd__9_, fe_pc_gen_branch_metadata_fwd__8_, fe_pc_gen_branch_metadata_fwd__7_, fe_pc_gen_branch_metadata_fwd__6_, fe_pc_gen_branch_metadata_fwd__5_, fe_pc_gen_branch_metadata_fwd__4_, fe_pc_gen_branch_metadata_fwd__3_, fe_pc_gen_branch_metadata_fwd__2_, fe_pc_gen_branch_metadata_fwd__1_, fe_pc_gen_branch_metadata_fwd__0_, fe_pc_gen_pc_redirect_valid_, N7 }),
    .fe_pc_gen_v_i(bp_fe_cmd_v_i),
    .fe_pc_gen_ready_o(bp_fe_cmd_ready_o)
  );


  icache_eaddr_width_p64_data_width_p64_inst_width_p32_tag_width_p10_num_cce_p1_num_lce_p2_ways_p8_lce_sets_p64_block_size_in_bytes_p8
  icache_1
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .id_i(icache_id_i[0]),
    .pc_gen_icache_vaddr_i(pc_gen_icache),
    .pc_gen_icache_vaddr_v_i(pc_gen_icache_v),
    .pc_gen_icache_vaddr_ready_o(pc_gen_icache_ready),
    .icache_pc_gen_data_o(icache_pc_gen),
    .icache_pc_gen_data_v_o(icache_pc_gen_v),
    .icache_pc_gen_data_ready_i(icache_pc_gen_ready),
    .itlb_icache_data_resp_i(itlb_icache),
    .itlb_icache_data_resp_v_i(itlb_icache_data_resp_v),
    .itlb_icache_data_resp_ready_o(itlb_icache_data_resp_ready),
    .cache_miss_o(cache_miss),
    .poison_i(poison),
    .lce_req_o(lce_cce_req_o),
    .lce_req_v_o(lce_cce_req_v_o),
    .lce_req_ready_i(lce_cce_req_ready_i),
    .lce_resp_o(lce_cce_resp_o),
    .lce_resp_v_o(lce_cce_resp_v_o),
    .lce_resp_ready_i(lce_cce_resp_ready_i),
    .lce_data_resp_o(lce_cce_data_resp_o),
    .lce_data_resp_v_o(lce_cce_data_resp_v_o),
    .lce_data_resp_ready_i(lce_cce_data_resp_ready_i),
    .lce_cmd_i(cce_lce_cmd_i),
    .lce_cmd_v_i(cce_lce_cmd_v_i),
    .lce_cmd_ready_o(cce_lce_cmd_ready_o),
    .lce_data_cmd_i(cce_lce_data_cmd_i),
    .lce_data_cmd_v_i(cce_lce_data_cmd_v_i),
    .lce_data_cmd_ready_o(cce_lce_data_cmd_ready_o),
    .lce_tr_resp_i(lce_lce_tr_resp_i),
    .lce_tr_resp_v_i(lce_lce_tr_resp_v_i),
    .lce_tr_resp_ready_o(lce_lce_tr_resp_ready_o),
    .lce_tr_resp_o(lce_lce_tr_resp_o),
    .lce_tr_resp_v_o(lce_lce_tr_resp_v_o),
    .lce_tr_resp_ready_i(lce_lce_tr_resp_ready_i)
  );


  itlb_vaddr_width_p56_paddr_width_p22_eaddr_width_p64_btb_indx_width_p9_bht_indx_width_p5_ras_addr_width_p22_asid_width_p10_ppn_start_bit_p12_tag_width_p10
  itlb_1
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .fe_itlb_i(bp_fe_cmd_i),
    .fe_itlb_v_i(bp_fe_cmd_v_i),
    .fe_itlb_ready_o(fe_itlb_ready),
    .pc_gen_itlb_i(pc_gen_itlb),
    .pc_gen_itlb_v_i(pc_gen_itlb_v),
    .pc_gen_itlb_ready_o(pc_gen_itlb_ready),
    .itlb_icache_o(itlb_icache),
    .itlb_icache_data_resp_v_o(itlb_icache_data_resp_v),
    .itlb_icache_data_resp_ready_i(itlb_icache_data_resp_ready),
    .itlb_fe_o(itlb_fe_queue),
    .itlb_fe_v_o(itlb_fe_v),
    .itlb_fe_ready_i(bp_fe_queue_ready_i)
  );

  assign N4 = ~bp_fe_cmd_i[108];
  assign N5 = bp_fe_cmd_i[107] | N4;
  assign N6 = bp_fe_cmd_i[106] | N5;
  assign N7 = ~N6;
  assign N8 = ~bp_fe_cmd_i[106];
  assign N9 = bp_fe_cmd_i[107] | bp_fe_cmd_i[108];
  assign N10 = N8 | N9;
  assign N11 = ~N10;
  assign N12 = ~bp_fe_cmd_i[41];
  assign N13 = bp_fe_cmd_i[40] | N12;
  assign N14 = bp_fe_cmd_i[39] | N13;
  assign N15 = ~N14;
  assign N16 = ~bp_fe_cmd_i[107];
  assign N17 = ~bp_fe_cmd_i[106];
  assign N18 = N16 | bp_fe_cmd_i[108];
  assign N19 = N17 | N18;
  assign N20 = ~N19;
  assign N21 = ~bp_fe_cmd_i[106];
  assign N22 = bp_fe_cmd_i[107] | bp_fe_cmd_i[108];
  assign N23 = N21 | N22;
  assign N24 = ~N23;
  assign N25 = ~bp_fe_cmd_i[108];
  assign N26 = bp_fe_cmd_i[107] | N25;
  assign N27 = bp_fe_cmd_i[106] | N26;
  assign N28 = ~N27;
  assign { fe_pc_gen_branch_metadata_fwd__35_, fe_pc_gen_branch_metadata_fwd__34_, fe_pc_gen_branch_metadata_fwd__33_, fe_pc_gen_branch_metadata_fwd__32_, fe_pc_gen_branch_metadata_fwd__31_, fe_pc_gen_branch_metadata_fwd__30_, fe_pc_gen_branch_metadata_fwd__29_, fe_pc_gen_branch_metadata_fwd__28_, fe_pc_gen_branch_metadata_fwd__27_, fe_pc_gen_branch_metadata_fwd__26_, fe_pc_gen_branch_metadata_fwd__25_, fe_pc_gen_branch_metadata_fwd__24_, fe_pc_gen_branch_metadata_fwd__23_, fe_pc_gen_branch_metadata_fwd__22_, fe_pc_gen_branch_metadata_fwd__21_, fe_pc_gen_branch_metadata_fwd__20_, fe_pc_gen_branch_metadata_fwd__19_, fe_pc_gen_branch_metadata_fwd__18_, fe_pc_gen_branch_metadata_fwd__17_, fe_pc_gen_branch_metadata_fwd__16_, fe_pc_gen_branch_metadata_fwd__15_, fe_pc_gen_branch_metadata_fwd__14_, fe_pc_gen_branch_metadata_fwd__13_, fe_pc_gen_branch_metadata_fwd__12_, fe_pc_gen_branch_metadata_fwd__11_, fe_pc_gen_branch_metadata_fwd__10_, fe_pc_gen_branch_metadata_fwd__9_, fe_pc_gen_branch_metadata_fwd__8_, fe_pc_gen_branch_metadata_fwd__7_, fe_pc_gen_branch_metadata_fwd__6_, fe_pc_gen_branch_metadata_fwd__5_, fe_pc_gen_branch_metadata_fwd__4_, fe_pc_gen_branch_metadata_fwd__3_, fe_pc_gen_branch_metadata_fwd__2_, fe_pc_gen_branch_metadata_fwd__1_, fe_pc_gen_branch_metadata_fwd__0_ } = (N0)? bp_fe_cmd_i[41:6] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N1)? bp_fe_cmd_i[38:3] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N28;
  assign N1 = N24;
  assign fe_pc_gen_pc_redirect_valid_ = N11 & N15;
  assign N2 = N24 | N28;
  assign N3 = ~N2;
  assign poison = cache_miss & N20;

endmodule

