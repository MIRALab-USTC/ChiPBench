VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MACRO bsg_mem_p570
  FOREIGN bsg_mem_p570 0 0 ;
  CLASS BLOCK ;
  SIZE 161.495 BY 81.75 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 79.715 160.36 79.885 ;
        RECT  1.14 76.915 160.36 77.085 ;
        RECT  1.14 74.115 160.36 74.285 ;
        RECT  1.14 71.315 160.36 71.485 ;
        RECT  1.14 68.515 160.36 68.685 ;
        RECT  1.14 65.715 160.36 65.885 ;
        RECT  1.14 62.915 160.36 63.085 ;
        RECT  1.14 60.115 160.36 60.285 ;
        RECT  1.14 57.315 160.36 57.485 ;
        RECT  1.14 54.515 160.36 54.685 ;
        RECT  1.14 51.715 160.36 51.885 ;
        RECT  1.14 48.915 160.36 49.085 ;
        RECT  1.14 46.115 160.36 46.285 ;
        RECT  1.14 43.315 160.36 43.485 ;
        RECT  1.14 40.515 160.36 40.685 ;
        RECT  1.14 37.715 160.36 37.885 ;
        RECT  1.14 34.915 160.36 35.085 ;
        RECT  1.14 32.115 160.36 32.285 ;
        RECT  1.14 29.315 160.36 29.485 ;
        RECT  1.14 26.515 160.36 26.685 ;
        RECT  1.14 23.715 160.36 23.885 ;
        RECT  1.14 20.915 160.36 21.085 ;
        RECT  1.14 18.115 160.36 18.285 ;
        RECT  1.14 15.315 160.36 15.485 ;
        RECT  1.14 12.515 160.36 12.685 ;
        RECT  1.14 9.715 160.36 9.885 ;
        RECT  1.14 6.915 160.36 7.085 ;
        RECT  1.14 4.115 160.36 4.285 ;
        RECT  1.14 1.315 160.36 1.485 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 78.315 160.36 78.485 ;
        RECT  1.14 75.515 160.36 75.685 ;
        RECT  1.14 72.715 160.36 72.885 ;
        RECT  1.14 69.915 160.36 70.085 ;
        RECT  1.14 67.115 160.36 67.285 ;
        RECT  1.14 64.315 160.36 64.485 ;
        RECT  1.14 61.515 160.36 61.685 ;
        RECT  1.14 58.715 160.36 58.885 ;
        RECT  1.14 55.915 160.36 56.085 ;
        RECT  1.14 53.115 160.36 53.285 ;
        RECT  1.14 50.315 160.36 50.485 ;
        RECT  1.14 47.515 160.36 47.685 ;
        RECT  1.14 44.715 160.36 44.885 ;
        RECT  1.14 41.915 160.36 42.085 ;
        RECT  1.14 39.115 160.36 39.285 ;
        RECT  1.14 36.315 160.36 36.485 ;
        RECT  1.14 33.515 160.36 33.685 ;
        RECT  1.14 30.715 160.36 30.885 ;
        RECT  1.14 27.915 160.36 28.085 ;
        RECT  1.14 25.115 160.36 25.285 ;
        RECT  1.14 22.315 160.36 22.485 ;
        RECT  1.14 19.515 160.36 19.685 ;
        RECT  1.14 16.715 160.36 16.885 ;
        RECT  1.14 13.915 160.36 14.085 ;
        RECT  1.14 11.115 160.36 11.285 ;
        RECT  1.14 8.315 160.36 8.485 ;
        RECT  1.14 5.515 160.36 5.685 ;
        RECT  1.14 2.715 160.36 2.885 ;
    END
  END VDD
  PIN r_addr_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 38.675 0.07 38.745 ;
    END
  END r_addr_i
  PIN r_data_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  132.185 0 132.325 0.14 ;
    END
  END r_data_o[0]
  PIN r_data_o[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  38.105 81.61 38.245 81.75 ;
    END
  END r_data_o[100]
  PIN r_data_o[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 77.875 0.07 77.945 ;
    END
  END r_data_o[101]
  PIN r_data_o[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  106.425 81.61 106.565 81.75 ;
    END
  END r_data_o[102]
  PIN r_data_o[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  15.705 81.61 15.845 81.75 ;
    END
  END r_data_o[103]
  PIN r_data_o[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 22.435 161.495 22.505 ;
    END
  END r_data_o[104]
  PIN r_data_o[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 52.955 0.07 53.025 ;
    END
  END r_data_o[105]
  PIN r_data_o[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  28.025 0 28.165 0.14 ;
    END
  END r_data_o[106]
  PIN r_data_o[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 3.395 0.07 3.465 ;
    END
  END r_data_o[107]
  PIN r_data_o[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 11.515 0.07 11.585 ;
    END
  END r_data_o[108]
  PIN r_data_o[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  89.625 0 89.765 0.14 ;
    END
  END r_data_o[109]
  PIN r_data_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 71.435 0.07 71.505 ;
    END
  END r_data_o[10]
  PIN r_data_o[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  48.745 81.61 48.885 81.75 ;
    END
  END r_data_o[110]
  PIN r_data_o[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 28.595 0.07 28.665 ;
    END
  END r_data_o[111]
  PIN r_data_o[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 46.235 161.495 46.305 ;
    END
  END r_data_o[112]
  PIN r_data_o[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 70.875 0.07 70.945 ;
    END
  END r_data_o[113]
  PIN r_data_o[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 61.635 0.07 61.705 ;
    END
  END r_data_o[114]
  PIN r_data_o[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 1.435 0.07 1.505 ;
    END
  END r_data_o[115]
  PIN r_data_o[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  48.185 0 48.325 0.14 ;
    END
  END r_data_o[116]
  PIN r_data_o[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 62.475 161.495 62.545 ;
    END
  END r_data_o[117]
  PIN r_data_o[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 6.755 0.07 6.825 ;
    END
  END r_data_o[118]
  PIN r_data_o[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 55.755 0.07 55.825 ;
    END
  END r_data_o[119]
  PIN r_data_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  86.265 0 86.405 0.14 ;
    END
  END r_data_o[11]
  PIN r_data_o[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 71.995 161.495 72.065 ;
    END
  END r_data_o[120]
  PIN r_data_o[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.665 0 10.805 0.14 ;
    END
  END r_data_o[121]
  PIN r_data_o[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  40.905 0 41.045 0.14 ;
    END
  END r_data_o[122]
  PIN r_data_o[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  117.625 81.61 117.765 81.75 ;
    END
  END r_data_o[123]
  PIN r_data_o[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 24.395 0.07 24.465 ;
    END
  END r_data_o[124]
  PIN r_data_o[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  70.585 0 70.725 0.14 ;
    END
  END r_data_o[125]
  PIN r_data_o[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 55.475 161.495 55.545 ;
    END
  END r_data_o[126]
  PIN r_data_o[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 71.155 0.07 71.225 ;
    END
  END r_data_o[127]
  PIN r_data_o[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 13.755 0.07 13.825 ;
    END
  END r_data_o[128]
  PIN r_data_o[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  81.225 0 81.365 0.14 ;
    END
  END r_data_o[129]
  PIN r_data_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  109.785 0 109.925 0.14 ;
    END
  END r_data_o[12]
  PIN r_data_o[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 78.995 0.07 79.065 ;
    END
  END r_data_o[130]
  PIN r_data_o[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  22.425 81.61 22.565 81.75 ;
    END
  END r_data_o[131]
  PIN r_data_o[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 0.875 161.495 0.945 ;
    END
  END r_data_o[132]
  PIN r_data_o[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  150.665 81.61 150.805 81.75 ;
    END
  END r_data_o[133]
  PIN r_data_o[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  48.185 81.61 48.325 81.75 ;
    END
  END r_data_o[134]
  PIN r_data_o[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 40.075 0.07 40.145 ;
    END
  END r_data_o[135]
  PIN r_data_o[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 69.755 0.07 69.825 ;
    END
  END r_data_o[136]
  PIN r_data_o[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  78.985 0 79.125 0.14 ;
    END
  END r_data_o[137]
  PIN r_data_o[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  35.305 81.61 35.445 81.75 ;
    END
  END r_data_o[138]
  PIN r_data_o[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 50.155 0.07 50.225 ;
    END
  END r_data_o[139]
  PIN r_data_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 14.035 0.07 14.105 ;
    END
  END r_data_o[13]
  PIN r_data_o[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 37.275 0.07 37.345 ;
    END
  END r_data_o[140]
  PIN r_data_o[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 79.275 161.495 79.345 ;
    END
  END r_data_o[141]
  PIN r_data_o[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 24.115 0.07 24.185 ;
    END
  END r_data_o[142]
  PIN r_data_o[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  30.265 81.61 30.405 81.75 ;
    END
  END r_data_o[143]
  PIN r_data_o[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 44.555 161.495 44.625 ;
    END
  END r_data_o[144]
  PIN r_data_o[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  106.985 81.61 107.125 81.75 ;
    END
  END r_data_o[145]
  PIN r_data_o[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 64.155 161.495 64.225 ;
    END
  END r_data_o[146]
  PIN r_data_o[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  78.425 81.61 78.565 81.75 ;
    END
  END r_data_o[147]
  PIN r_data_o[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 79.555 0.07 79.625 ;
    END
  END r_data_o[148]
  PIN r_data_o[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  87.945 81.61 88.085 81.75 ;
    END
  END r_data_o[149]
  PIN r_data_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  143.945 81.61 144.085 81.75 ;
    END
  END r_data_o[14]
  PIN r_data_o[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 10.115 161.495 10.185 ;
    END
  END r_data_o[150]
  PIN r_data_o[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  86.265 81.61 86.405 81.75 ;
    END
  END r_data_o[151]
  PIN r_data_o[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  77.305 81.61 77.445 81.75 ;
    END
  END r_data_o[152]
  PIN r_data_o[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 68.355 0.07 68.425 ;
    END
  END r_data_o[153]
  PIN r_data_o[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  61.625 81.61 61.765 81.75 ;
    END
  END r_data_o[154]
  PIN r_data_o[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  154.025 81.61 154.165 81.75 ;
    END
  END r_data_o[155]
  PIN r_data_o[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 4.795 0.07 4.865 ;
    END
  END r_data_o[156]
  PIN r_data_o[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 76.475 161.495 76.545 ;
    END
  END r_data_o[157]
  PIN r_data_o[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 57.155 0.07 57.225 ;
    END
  END r_data_o[158]
  PIN r_data_o[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  159.065 81.61 159.205 81.75 ;
    END
  END r_data_o[159]
  PIN r_data_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 42.035 0.07 42.105 ;
    END
  END r_data_o[15]
  PIN r_data_o[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  67.785 81.61 67.925 81.75 ;
    END
  END r_data_o[160]
  PIN r_data_o[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  104.745 0 104.885 0.14 ;
    END
  END r_data_o[161]
  PIN r_data_o[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 64.995 161.495 65.065 ;
    END
  END r_data_o[162]
  PIN r_data_o[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 21.595 161.495 21.665 ;
    END
  END r_data_o[163]
  PIN r_data_o[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 36.715 161.495 36.785 ;
    END
  END r_data_o[164]
  PIN r_data_o[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  54.905 0 55.045 0.14 ;
    END
  END r_data_o[165]
  PIN r_data_o[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  108.665 81.61 108.805 81.75 ;
    END
  END r_data_o[166]
  PIN r_data_o[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  128.265 81.61 128.405 81.75 ;
    END
  END r_data_o[167]
  PIN r_data_o[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.075 0.07 12.145 ;
    END
  END r_data_o[168]
  PIN r_data_o[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  131.625 0 131.765 0.14 ;
    END
  END r_data_o[169]
  PIN r_data_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  45.385 81.61 45.525 81.75 ;
    END
  END r_data_o[16]
  PIN r_data_o[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  53.785 0 53.925 0.14 ;
    END
  END r_data_o[170]
  PIN r_data_o[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 31.115 161.495 31.185 ;
    END
  END r_data_o[171]
  PIN r_data_o[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  45.945 0 46.085 0.14 ;
    END
  END r_data_o[172]
  PIN r_data_o[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  11.785 81.61 11.925 81.75 ;
    END
  END r_data_o[173]
  PIN r_data_o[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 70.595 0.07 70.665 ;
    END
  END r_data_o[174]
  PIN r_data_o[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 28.315 161.495 28.385 ;
    END
  END r_data_o[175]
  PIN r_data_o[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  39.225 0 39.365 0.14 ;
    END
  END r_data_o[176]
  PIN r_data_o[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  87.945 0 88.085 0.14 ;
    END
  END r_data_o[177]
  PIN r_data_o[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 56.035 161.495 56.105 ;
    END
  END r_data_o[178]
  PIN r_data_o[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 12.635 161.495 12.705 ;
    END
  END r_data_o[179]
  PIN r_data_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 45.115 161.495 45.185 ;
    END
  END r_data_o[17]
  PIN r_data_o[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  1.145 0 1.285 0.14 ;
    END
  END r_data_o[180]
  PIN r_data_o[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 8.995 0.07 9.065 ;
    END
  END r_data_o[181]
  PIN r_data_o[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 9.555 0.07 9.625 ;
    END
  END r_data_o[182]
  PIN r_data_o[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 4.235 161.495 4.305 ;
    END
  END r_data_o[183]
  PIN r_data_o[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  150.105 81.61 150.245 81.75 ;
    END
  END r_data_o[184]
  PIN r_data_o[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 17.955 161.495 18.025 ;
    END
  END r_data_o[185]
  PIN r_data_o[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 57.715 0.07 57.785 ;
    END
  END r_data_o[186]
  PIN r_data_o[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 76.195 161.495 76.265 ;
    END
  END r_data_o[187]
  PIN r_data_o[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 78.435 0.07 78.505 ;
    END
  END r_data_o[188]
  PIN r_data_o[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  76.185 81.61 76.325 81.75 ;
    END
  END r_data_o[189]
  PIN r_data_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  36.425 81.61 36.565 81.75 ;
    END
  END r_data_o[18]
  PIN r_data_o[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  105.305 0 105.445 0.14 ;
    END
  END r_data_o[190]
  PIN r_data_o[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 78.995 161.495 79.065 ;
    END
  END r_data_o[191]
  PIN r_data_o[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  42.025 81.61 42.165 81.75 ;
    END
  END r_data_o[192]
  PIN r_data_o[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 47.915 0.07 47.985 ;
    END
  END r_data_o[193]
  PIN r_data_o[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 64.155 0.07 64.225 ;
    END
  END r_data_o[194]
  PIN r_data_o[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  85.145 81.61 85.285 81.75 ;
    END
  END r_data_o[195]
  PIN r_data_o[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 67.795 0.07 67.865 ;
    END
  END r_data_o[196]
  PIN r_data_o[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  60.505 0 60.645 0.14 ;
    END
  END r_data_o[197]
  PIN r_data_o[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 66.675 161.495 66.745 ;
    END
  END r_data_o[198]
  PIN r_data_o[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 53.235 0.07 53.305 ;
    END
  END r_data_o[199]
  PIN r_data_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 60.515 0.07 60.585 ;
    END
  END r_data_o[19]
  PIN r_data_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 47.635 161.495 47.705 ;
    END
  END r_data_o[1]
  PIN r_data_o[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  24.105 0 24.245 0.14 ;
    END
  END r_data_o[200]
  PIN r_data_o[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 61.635 161.495 61.705 ;
    END
  END r_data_o[201]
  PIN r_data_o[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 19.915 161.495 19.985 ;
    END
  END r_data_o[202]
  PIN r_data_o[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 32.235 161.495 32.305 ;
    END
  END r_data_o[203]
  PIN r_data_o[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 41.195 0.07 41.265 ;
    END
  END r_data_o[204]
  PIN r_data_o[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  73.945 81.61 74.085 81.75 ;
    END
  END r_data_o[205]
  PIN r_data_o[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  58.265 0 58.405 0.14 ;
    END
  END r_data_o[206]
  PIN r_data_o[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 53.795 0.07 53.865 ;
    END
  END r_data_o[207]
  PIN r_data_o[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 60.235 161.495 60.305 ;
    END
  END r_data_o[208]
  PIN r_data_o[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 42.595 161.495 42.665 ;
    END
  END r_data_o[209]
  PIN r_data_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.915 0.07 12.985 ;
    END
  END r_data_o[20]
  PIN r_data_o[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 45.115 0.07 45.185 ;
    END
  END r_data_o[210]
  PIN r_data_o[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  57.145 81.61 57.285 81.75 ;
    END
  END r_data_o[211]
  PIN r_data_o[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 54.635 0.07 54.705 ;
    END
  END r_data_o[212]
  PIN r_data_o[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 17.675 0.07 17.745 ;
    END
  END r_data_o[213]
  PIN r_data_o[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  159.625 0 159.765 0.14 ;
    END
  END r_data_o[214]
  PIN r_data_o[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 71.435 161.495 71.505 ;
    END
  END r_data_o[215]
  PIN r_data_o[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  69.465 0 69.605 0.14 ;
    END
  END r_data_o[216]
  PIN r_data_o[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  142.825 0 142.965 0.14 ;
    END
  END r_data_o[217]
  PIN r_data_o[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  113.705 81.61 113.845 81.75 ;
    END
  END r_data_o[218]
  PIN r_data_o[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 20.475 161.495 20.545 ;
    END
  END r_data_o[219]
  PIN r_data_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 54.915 161.495 54.985 ;
    END
  END r_data_o[21]
  PIN r_data_o[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  148.985 0 149.125 0.14 ;
    END
  END r_data_o[220]
  PIN r_data_o[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 47.075 161.495 47.145 ;
    END
  END r_data_o[221]
  PIN r_data_o[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  82.345 81.61 82.485 81.75 ;
    END
  END r_data_o[222]
  PIN r_data_o[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  138.905 81.61 139.045 81.75 ;
    END
  END r_data_o[223]
  PIN r_data_o[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 3.955 0.07 4.025 ;
    END
  END r_data_o[224]
  PIN r_data_o[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  32.505 0 32.645 0.14 ;
    END
  END r_data_o[225]
  PIN r_data_o[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  64.425 81.61 64.565 81.75 ;
    END
  END r_data_o[226]
  PIN r_data_o[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 17.675 161.495 17.745 ;
    END
  END r_data_o[227]
  PIN r_data_o[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  43.705 0 43.845 0.14 ;
    END
  END r_data_o[228]
  PIN r_data_o[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  2.825 0 2.965 0.14 ;
    END
  END r_data_o[229]
  PIN r_data_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 80.115 161.495 80.185 ;
    END
  END r_data_o[22]
  PIN r_data_o[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 24.395 161.495 24.465 ;
    END
  END r_data_o[230]
  PIN r_data_o[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 72.275 0.07 72.345 ;
    END
  END r_data_o[231]
  PIN r_data_o[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 54.355 0.07 54.425 ;
    END
  END r_data_o[232]
  PIN r_data_o[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 72.835 0.07 72.905 ;
    END
  END r_data_o[233]
  PIN r_data_o[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 80.115 0.07 80.185 ;
    END
  END r_data_o[234]
  PIN r_data_o[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 65.275 161.495 65.345 ;
    END
  END r_data_o[235]
  PIN r_data_o[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  37.545 81.61 37.685 81.75 ;
    END
  END r_data_o[236]
  PIN r_data_o[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  50.425 0 50.565 0.14 ;
    END
  END r_data_o[237]
  PIN r_data_o[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 17.115 161.495 17.185 ;
    END
  END r_data_o[238]
  PIN r_data_o[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 10.955 0.07 11.025 ;
    END
  END r_data_o[239]
  PIN r_data_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 59.395 161.495 59.465 ;
    END
  END r_data_o[23]
  PIN r_data_o[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 69.475 0.07 69.545 ;
    END
  END r_data_o[240]
  PIN r_data_o[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  122.665 81.61 122.805 81.75 ;
    END
  END r_data_o[241]
  PIN r_data_o[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 42.875 161.495 42.945 ;
    END
  END r_data_o[242]
  PIN r_data_o[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  127.705 0 127.845 0.14 ;
    END
  END r_data_o[243]
  PIN r_data_o[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 53.795 161.495 53.865 ;
    END
  END r_data_o[244]
  PIN r_data_o[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  44.825 81.61 44.965 81.75 ;
    END
  END r_data_o[245]
  PIN r_data_o[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 75.355 161.495 75.425 ;
    END
  END r_data_o[246]
  PIN r_data_o[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 61.355 0.07 61.425 ;
    END
  END r_data_o[247]
  PIN r_data_o[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 38.955 0.07 39.025 ;
    END
  END r_data_o[248]
  PIN r_data_o[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 6.755 161.495 6.825 ;
    END
  END r_data_o[249]
  PIN r_data_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  141.705 0 141.845 0.14 ;
    END
  END r_data_o[24]
  PIN r_data_o[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 29.995 161.495 30.065 ;
    END
  END r_data_o[250]
  PIN r_data_o[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  78.985 81.61 79.125 81.75 ;
    END
  END r_data_o[251]
  PIN r_data_o[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 79.835 161.495 79.905 ;
    END
  END r_data_o[252]
  PIN r_data_o[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 25.795 0.07 25.865 ;
    END
  END r_data_o[253]
  PIN r_data_o[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  98.585 0 98.725 0.14 ;
    END
  END r_data_o[254]
  PIN r_data_o[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 33.355 161.495 33.425 ;
    END
  END r_data_o[255]
  PIN r_data_o[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 9.835 161.495 9.905 ;
    END
  END r_data_o[256]
  PIN r_data_o[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 49.595 0.07 49.665 ;
    END
  END r_data_o[257]
  PIN r_data_o[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  38.665 0 38.805 0.14 ;
    END
  END r_data_o[258]
  PIN r_data_o[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 77.035 0.07 77.105 ;
    END
  END r_data_o[259]
  PIN r_data_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  70.025 0 70.165 0.14 ;
    END
  END r_data_o[25]
  PIN r_data_o[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  123.785 81.61 123.925 81.75 ;
    END
  END r_data_o[260]
  PIN r_data_o[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  101.385 0 101.525 0.14 ;
    END
  END r_data_o[261]
  PIN r_data_o[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 17.395 161.495 17.465 ;
    END
  END r_data_o[262]
  PIN r_data_o[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  30.265 0 30.405 0.14 ;
    END
  END r_data_o[263]
  PIN r_data_o[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.675 0.07 31.745 ;
    END
  END r_data_o[264]
  PIN r_data_o[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 36.715 0.07 36.785 ;
    END
  END r_data_o[265]
  PIN r_data_o[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 46.515 161.495 46.585 ;
    END
  END r_data_o[266]
  PIN r_data_o[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  2.265 81.61 2.405 81.75 ;
    END
  END r_data_o[267]
  PIN r_data_o[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 56.035 0.07 56.105 ;
    END
  END r_data_o[268]
  PIN r_data_o[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 56.595 161.495 56.665 ;
    END
  END r_data_o[269]
  PIN r_data_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 55.755 161.495 55.825 ;
    END
  END r_data_o[26]
  PIN r_data_o[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 67.515 161.495 67.585 ;
    END
  END r_data_o[270]
  PIN r_data_o[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  59.945 0 60.085 0.14 ;
    END
  END r_data_o[271]
  PIN r_data_o[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  146.745 81.61 146.885 81.75 ;
    END
  END r_data_o[272]
  PIN r_data_o[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 71.715 161.495 71.785 ;
    END
  END r_data_o[273]
  PIN r_data_o[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 20.195 0.07 20.265 ;
    END
  END r_data_o[274]
  PIN r_data_o[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  109.225 0 109.365 0.14 ;
    END
  END r_data_o[275]
  PIN r_data_o[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 50.715 0.07 50.785 ;
    END
  END r_data_o[276]
  PIN r_data_o[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 43.435 0.07 43.505 ;
    END
  END r_data_o[277]
  PIN r_data_o[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 77.035 161.495 77.105 ;
    END
  END r_data_o[278]
  PIN r_data_o[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  141.705 81.61 141.845 81.75 ;
    END
  END r_data_o[279]
  PIN r_data_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  36.425 0 36.565 0.14 ;
    END
  END r_data_o[27]
  PIN r_data_o[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 65.835 161.495 65.905 ;
    END
  END r_data_o[280]
  PIN r_data_o[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 34.755 161.495 34.825 ;
    END
  END r_data_o[281]
  PIN r_data_o[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  40.345 81.61 40.485 81.75 ;
    END
  END r_data_o[282]
  PIN r_data_o[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  116.505 0 116.645 0.14 ;
    END
  END r_data_o[283]
  PIN r_data_o[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 69.195 0.07 69.265 ;
    END
  END r_data_o[284]
  PIN r_data_o[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  93.545 0 93.685 0.14 ;
    END
  END r_data_o[285]
  PIN r_data_o[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 12.915 161.495 12.985 ;
    END
  END r_data_o[286]
  PIN r_data_o[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 61.075 161.495 61.145 ;
    END
  END r_data_o[287]
  PIN r_data_o[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 59.115 161.495 59.185 ;
    END
  END r_data_o[288]
  PIN r_data_o[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  62.745 0 62.885 0.14 ;
    END
  END r_data_o[289]
  PIN r_data_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 18.235 0.07 18.305 ;
    END
  END r_data_o[28]
  PIN r_data_o[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 75.355 0.07 75.425 ;
    END
  END r_data_o[290]
  PIN r_data_o[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  58.825 81.61 58.965 81.75 ;
    END
  END r_data_o[291]
  PIN r_data_o[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  158.505 0 158.645 0.14 ;
    END
  END r_data_o[292]
  PIN r_data_o[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  29.145 81.61 29.285 81.75 ;
    END
  END r_data_o[293]
  PIN r_data_o[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  48.745 0 48.885 0.14 ;
    END
  END r_data_o[294]
  PIN r_data_o[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 26.075 0.07 26.145 ;
    END
  END r_data_o[295]
  PIN r_data_o[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  29.705 0 29.845 0.14 ;
    END
  END r_data_o[296]
  PIN r_data_o[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  72.265 0 72.405 0.14 ;
    END
  END r_data_o[297]
  PIN r_data_o[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 29.995 0.07 30.065 ;
    END
  END r_data_o[298]
  PIN r_data_o[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  90.745 81.61 90.885 81.75 ;
    END
  END r_data_o[299]
  PIN r_data_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  54.905 81.61 55.045 81.75 ;
    END
  END r_data_o[29]
  PIN r_data_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  81.785 0 81.925 0.14 ;
    END
  END r_data_o[2]
  PIN r_data_o[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  110.905 81.61 111.045 81.75 ;
    END
  END r_data_o[300]
  PIN r_data_o[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  33.625 81.61 33.765 81.75 ;
    END
  END r_data_o[301]
  PIN r_data_o[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  157.945 0 158.085 0.14 ;
    END
  END r_data_o[302]
  PIN r_data_o[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 2.555 0.07 2.625 ;
    END
  END r_data_o[303]
  PIN r_data_o[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 32.515 0.07 32.585 ;
    END
  END r_data_o[304]
  PIN r_data_o[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  80.665 81.61 80.805 81.75 ;
    END
  END r_data_o[305]
  PIN r_data_o[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 9.835 0.07 9.905 ;
    END
  END r_data_o[306]
  PIN r_data_o[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 38.955 161.495 39.025 ;
    END
  END r_data_o[307]
  PIN r_data_o[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  140.025 0 140.165 0.14 ;
    END
  END r_data_o[308]
  PIN r_data_o[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  1.705 0 1.845 0.14 ;
    END
  END r_data_o[309]
  PIN r_data_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  81.785 81.61 81.925 81.75 ;
    END
  END r_data_o[30]
  PIN r_data_o[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 11.795 161.495 11.865 ;
    END
  END r_data_o[310]
  PIN r_data_o[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 43.155 161.495 43.225 ;
    END
  END r_data_o[311]
  PIN r_data_o[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 20.475 0.07 20.545 ;
    END
  END r_data_o[312]
  PIN r_data_o[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  44.265 0 44.405 0.14 ;
    END
  END r_data_o[313]
  PIN r_data_o[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 60.795 0.07 60.865 ;
    END
  END r_data_o[314]
  PIN r_data_o[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  33.625 0 33.765 0.14 ;
    END
  END r_data_o[315]
  PIN r_data_o[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 7.595 161.495 7.665 ;
    END
  END r_data_o[316]
  PIN r_data_o[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 74.515 161.495 74.585 ;
    END
  END r_data_o[317]
  PIN r_data_o[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  76.745 0 76.885 0.14 ;
    END
  END r_data_o[318]
  PIN r_data_o[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 8.155 161.495 8.225 ;
    END
  END r_data_o[319]
  PIN r_data_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 28.595 161.495 28.665 ;
    END
  END r_data_o[31]
  PIN r_data_o[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  155.145 0 155.285 0.14 ;
    END
  END r_data_o[320]
  PIN r_data_o[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 46.795 161.495 46.865 ;
    END
  END r_data_o[321]
  PIN r_data_o[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  99.145 0 99.285 0.14 ;
    END
  END r_data_o[322]
  PIN r_data_o[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  53.225 0 53.365 0.14 ;
    END
  END r_data_o[323]
  PIN r_data_o[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 34.195 161.495 34.265 ;
    END
  END r_data_o[324]
  PIN r_data_o[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  104.745 81.61 104.885 81.75 ;
    END
  END r_data_o[325]
  PIN r_data_o[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  84.025 0 84.165 0.14 ;
    END
  END r_data_o[326]
  PIN r_data_o[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  126.585 81.61 126.725 81.75 ;
    END
  END r_data_o[327]
  PIN r_data_o[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 10.955 161.495 11.025 ;
    END
  END r_data_o[328]
  PIN r_data_o[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  147.305 81.61 147.445 81.75 ;
    END
  END r_data_o[329]
  PIN r_data_o[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.185 0 34.325 0.14 ;
    END
  END r_data_o[32]
  PIN r_data_o[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 23.555 161.495 23.625 ;
    END
  END r_data_o[330]
  PIN r_data_o[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 23.835 0.07 23.905 ;
    END
  END r_data_o[331]
  PIN r_data_o[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  21.865 81.61 22.005 81.75 ;
    END
  END r_data_o[332]
  PIN r_data_o[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 16.835 0.07 16.905 ;
    END
  END r_data_o[333]
  PIN r_data_o[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  55.465 0 55.605 0.14 ;
    END
  END r_data_o[334]
  PIN r_data_o[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 30.835 161.495 30.905 ;
    END
  END r_data_o[335]
  PIN r_data_o[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 40.355 0.07 40.425 ;
    END
  END r_data_o[336]
  PIN r_data_o[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 40.915 161.495 40.985 ;
    END
  END r_data_o[337]
  PIN r_data_o[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.905 0 13.045 0.14 ;
    END
  END r_data_o[338]
  PIN r_data_o[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  77.305 0 77.445 0.14 ;
    END
  END r_data_o[339]
  PIN r_data_o[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 22.155 0.07 22.225 ;
    END
  END r_data_o[33]
  PIN r_data_o[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  22.425 0 22.565 0.14 ;
    END
  END r_data_o[340]
  PIN r_data_o[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 16.555 0.07 16.625 ;
    END
  END r_data_o[341]
  PIN r_data_o[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  135.545 0 135.685 0.14 ;
    END
  END r_data_o[342]
  PIN r_data_o[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  132.745 81.61 132.885 81.75 ;
    END
  END r_data_o[343]
  PIN r_data_o[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.955 0.07 32.025 ;
    END
  END r_data_o[344]
  PIN r_data_o[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 59.675 161.495 59.745 ;
    END
  END r_data_o[345]
  PIN r_data_o[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  130.505 81.61 130.645 81.75 ;
    END
  END r_data_o[346]
  PIN r_data_o[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 68.635 161.495 68.705 ;
    END
  END r_data_o[347]
  PIN r_data_o[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  108.105 81.61 108.245 81.75 ;
    END
  END r_data_o[348]
  PIN r_data_o[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 52.675 0.07 52.745 ;
    END
  END r_data_o[349]
  PIN r_data_o[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  152.345 81.61 152.485 81.75 ;
    END
  END r_data_o[34]
  PIN r_data_o[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 71.715 0.07 71.785 ;
    END
  END r_data_o[350]
  PIN r_data_o[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 39.235 161.495 39.305 ;
    END
  END r_data_o[351]
  PIN r_data_o[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  91.865 81.61 92.005 81.75 ;
    END
  END r_data_o[352]
  PIN r_data_o[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.305 81.61 7.445 81.75 ;
    END
  END r_data_o[353]
  PIN r_data_o[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  115.385 81.61 115.525 81.75 ;
    END
  END r_data_o[354]
  PIN r_data_o[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 74.235 0.07 74.305 ;
    END
  END r_data_o[355]
  PIN r_data_o[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 73.395 0.07 73.465 ;
    END
  END r_data_o[356]
  PIN r_data_o[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 26.635 0.07 26.705 ;
    END
  END r_data_o[357]
  PIN r_data_o[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  42.585 81.61 42.725 81.75 ;
    END
  END r_data_o[358]
  PIN r_data_o[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 8.715 0.07 8.785 ;
    END
  END r_data_o[359]
  PIN r_data_o[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 29.155 161.495 29.225 ;
    END
  END r_data_o[35]
  PIN r_data_o[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  89.065 0 89.205 0.14 ;
    END
  END r_data_o[360]
  PIN r_data_o[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  145.625 0 145.765 0.14 ;
    END
  END r_data_o[361]
  PIN r_data_o[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  120.985 0 121.125 0.14 ;
    END
  END r_data_o[362]
  PIN r_data_o[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 66.675 0.07 66.745 ;
    END
  END r_data_o[363]
  PIN r_data_o[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  155.705 81.61 155.845 81.75 ;
    END
  END r_data_o[364]
  PIN r_data_o[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  91.305 0 91.445 0.14 ;
    END
  END r_data_o[365]
  PIN r_data_o[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 3.115 161.495 3.185 ;
    END
  END r_data_o[366]
  PIN r_data_o[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  11.225 81.61 11.365 81.75 ;
    END
  END r_data_o[367]
  PIN r_data_o[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 46.515 0.07 46.585 ;
    END
  END r_data_o[368]
  PIN r_data_o[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 63.035 0.07 63.105 ;
    END
  END r_data_o[369]
  PIN r_data_o[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 15.435 161.495 15.505 ;
    END
  END r_data_o[36]
  PIN r_data_o[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  15.705 0 15.845 0.14 ;
    END
  END r_data_o[370]
  PIN r_data_o[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  19.625 0 19.765 0.14 ;
    END
  END r_data_o[371]
  PIN r_data_o[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  88.505 81.61 88.645 81.75 ;
    END
  END r_data_o[372]
  PIN r_data_o[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 18.515 161.495 18.585 ;
    END
  END r_data_o[373]
  PIN r_data_o[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  136.105 0 136.245 0.14 ;
    END
  END r_data_o[374]
  PIN r_data_o[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 62.195 0.07 62.265 ;
    END
  END r_data_o[375]
  PIN r_data_o[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  129.945 0 130.085 0.14 ;
    END
  END r_data_o[376]
  PIN r_data_o[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  89.065 81.61 89.205 81.75 ;
    END
  END r_data_o[377]
  PIN r_data_o[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  111.465 81.61 111.605 81.75 ;
    END
  END r_data_o[378]
  PIN r_data_o[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 38.115 161.495 38.185 ;
    END
  END r_data_o[379]
  PIN r_data_o[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 56.315 0.07 56.385 ;
    END
  END r_data_o[37]
  PIN r_data_o[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 27.755 0.07 27.825 ;
    END
  END r_data_o[380]
  PIN r_data_o[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  52.105 0 52.245 0.14 ;
    END
  END r_data_o[381]
  PIN r_data_o[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 66.955 0.07 67.025 ;
    END
  END r_data_o[382]
  PIN r_data_o[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 45.395 0.07 45.465 ;
    END
  END r_data_o[383]
  PIN r_data_o[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  15.145 0 15.285 0.14 ;
    END
  END r_data_o[384]
  PIN r_data_o[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  8.425 81.61 8.565 81.75 ;
    END
  END r_data_o[385]
  PIN r_data_o[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 50.995 0.07 51.065 ;
    END
  END r_data_o[386]
  PIN r_data_o[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 74.235 161.495 74.305 ;
    END
  END r_data_o[387]
  PIN r_data_o[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 75.915 0.07 75.985 ;
    END
  END r_data_o[388]
  PIN r_data_o[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  38.665 81.61 38.805 81.75 ;
    END
  END r_data_o[389]
  PIN r_data_o[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  39.785 81.61 39.925 81.75 ;
    END
  END r_data_o[38]
  PIN r_data_o[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  16.825 81.61 16.965 81.75 ;
    END
  END r_data_o[390]
  PIN r_data_o[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 15.715 0.07 15.785 ;
    END
  END r_data_o[391]
  PIN r_data_o[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.595 0.07 21.665 ;
    END
  END r_data_o[392]
  PIN r_data_o[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  65.545 0 65.685 0.14 ;
    END
  END r_data_o[393]
  PIN r_data_o[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  47.625 81.61 47.765 81.75 ;
    END
  END r_data_o[394]
  PIN r_data_o[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 65.275 0.07 65.345 ;
    END
  END r_data_o[395]
  PIN r_data_o[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 48.755 161.495 48.825 ;
    END
  END r_data_o[396]
  PIN r_data_o[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 29.435 161.495 29.505 ;
    END
  END r_data_o[397]
  PIN r_data_o[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  147.865 81.61 148.005 81.75 ;
    END
  END r_data_o[398]
  PIN r_data_o[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 17.395 0.07 17.465 ;
    END
  END r_data_o[399]
  PIN r_data_o[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  72.825 0 72.965 0.14 ;
    END
  END r_data_o[39]
  PIN r_data_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  21.305 81.61 21.445 81.75 ;
    END
  END r_data_o[3]
  PIN r_data_o[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 57.995 161.495 58.065 ;
    END
  END r_data_o[400]
  PIN r_data_o[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  56.585 0 56.725 0.14 ;
    END
  END r_data_o[401]
  PIN r_data_o[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  60.505 81.61 60.645 81.75 ;
    END
  END r_data_o[402]
  PIN r_data_o[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 54.915 0.07 54.985 ;
    END
  END r_data_o[403]
  PIN r_data_o[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 42.315 161.495 42.385 ;
    END
  END r_data_o[404]
  PIN r_data_o[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  66.105 81.61 66.245 81.75 ;
    END
  END r_data_o[405]
  PIN r_data_o[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  123.225 81.61 123.365 81.75 ;
    END
  END r_data_o[406]
  PIN r_data_o[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 24.675 0.07 24.745 ;
    END
  END r_data_o[407]
  PIN r_data_o[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 67.235 0.07 67.305 ;
    END
  END r_data_o[408]
  PIN r_data_o[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 48.755 0.07 48.825 ;
    END
  END r_data_o[409]
  PIN r_data_o[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  20.185 0 20.325 0.14 ;
    END
  END r_data_o[40]
  PIN r_data_o[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  77.865 81.61 78.005 81.75 ;
    END
  END r_data_o[410]
  PIN r_data_o[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  5.625 81.61 5.765 81.75 ;
    END
  END r_data_o[411]
  PIN r_data_o[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 81.61 0.725 81.75 ;
    END
  END r_data_o[412]
  PIN r_data_o[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  147.305 0 147.445 0.14 ;
    END
  END r_data_o[413]
  PIN r_data_o[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 44.275 161.495 44.345 ;
    END
  END r_data_o[414]
  PIN r_data_o[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 38.395 0.07 38.465 ;
    END
  END r_data_o[415]
  PIN r_data_o[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 24.955 0.07 25.025 ;
    END
  END r_data_o[416]
  PIN r_data_o[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 45.955 0.07 46.025 ;
    END
  END r_data_o[417]
  PIN r_data_o[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 75.635 161.495 75.705 ;
    END
  END r_data_o[418]
  PIN r_data_o[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 60.795 161.495 60.865 ;
    END
  END r_data_o[419]
  PIN r_data_o[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 7.035 161.495 7.105 ;
    END
  END r_data_o[41]
  PIN r_data_o[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 62.755 0.07 62.825 ;
    END
  END r_data_o[420]
  PIN r_data_o[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  117.065 0 117.205 0.14 ;
    END
  END r_data_o[421]
  PIN r_data_o[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  156.825 0 156.965 0.14 ;
    END
  END r_data_o[422]
  PIN r_data_o[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  50.985 0 51.125 0.14 ;
    END
  END r_data_o[423]
  PIN r_data_o[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  75.625 81.61 75.765 81.75 ;
    END
  END r_data_o[424]
  PIN r_data_o[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 35.875 0.07 35.945 ;
    END
  END r_data_o[425]
  PIN r_data_o[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  119.305 81.61 119.445 81.75 ;
    END
  END r_data_o[426]
  PIN r_data_o[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 60.235 0.07 60.305 ;
    END
  END r_data_o[427]
  PIN r_data_o[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 25.235 161.495 25.305 ;
    END
  END r_data_o[428]
  PIN r_data_o[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  58.265 81.61 58.405 81.75 ;
    END
  END r_data_o[429]
  PIN r_data_o[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 57.995 0.07 58.065 ;
    END
  END r_data_o[42]
  PIN r_data_o[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 1.715 0.07 1.785 ;
    END
  END r_data_o[430]
  PIN r_data_o[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 5.075 0.07 5.145 ;
    END
  END r_data_o[431]
  PIN r_data_o[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 25.795 161.495 25.865 ;
    END
  END r_data_o[432]
  PIN r_data_o[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  37.545 0 37.685 0.14 ;
    END
  END r_data_o[433]
  PIN r_data_o[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 70.315 0.07 70.385 ;
    END
  END r_data_o[434]
  PIN r_data_o[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 72.835 161.495 72.905 ;
    END
  END r_data_o[435]
  PIN r_data_o[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 21.875 161.495 21.945 ;
    END
  END r_data_o[436]
  PIN r_data_o[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  62.745 81.61 62.885 81.75 ;
    END
  END r_data_o[437]
  PIN r_data_o[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.115 0.07 31.185 ;
    END
  END r_data_o[438]
  PIN r_data_o[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 61.915 161.495 61.985 ;
    END
  END r_data_o[439]
  PIN r_data_o[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 41.475 0.07 41.545 ;
    END
  END r_data_o[43]
  PIN r_data_o[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 13.755 161.495 13.825 ;
    END
  END r_data_o[440]
  PIN r_data_o[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 50.995 161.495 51.065 ;
    END
  END r_data_o[441]
  PIN r_data_o[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  134.985 0 135.125 0.14 ;
    END
  END r_data_o[442]
  PIN r_data_o[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 67.235 161.495 67.305 ;
    END
  END r_data_o[443]
  PIN r_data_o[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 30.275 161.495 30.345 ;
    END
  END r_data_o[444]
  PIN r_data_o[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 49.875 0.07 49.945 ;
    END
  END r_data_o[445]
  PIN r_data_o[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 63.315 161.495 63.385 ;
    END
  END r_data_o[446]
  PIN r_data_o[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 76.755 0.07 76.825 ;
    END
  END r_data_o[447]
  PIN r_data_o[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  61.625 0 61.765 0.14 ;
    END
  END r_data_o[448]
  PIN r_data_o[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  57.145 0 57.285 0.14 ;
    END
  END r_data_o[449]
  PIN r_data_o[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 48.475 0.07 48.545 ;
    END
  END r_data_o[44]
  PIN r_data_o[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  75.065 0 75.205 0.14 ;
    END
  END r_data_o[450]
  PIN r_data_o[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  5.625 0 5.765 0.14 ;
    END
  END r_data_o[451]
  PIN r_data_o[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.105 81.61 10.245 81.75 ;
    END
  END r_data_o[452]
  PIN r_data_o[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 52.395 161.495 52.465 ;
    END
  END r_data_o[453]
  PIN r_data_o[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 74.515 0.07 74.585 ;
    END
  END r_data_o[454]
  PIN r_data_o[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  79.545 81.61 79.685 81.75 ;
    END
  END r_data_o[455]
  PIN r_data_o[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 49.035 0.07 49.105 ;
    END
  END r_data_o[456]
  PIN r_data_o[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  50.985 81.61 51.125 81.75 ;
    END
  END r_data_o[457]
  PIN r_data_o[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  75.625 0 75.765 0.14 ;
    END
  END r_data_o[458]
  PIN r_data_o[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 58.555 161.495 58.625 ;
    END
  END r_data_o[459]
  PIN r_data_o[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.875 0.07 21.945 ;
    END
  END r_data_o[45]
  PIN r_data_o[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  21.305 0 21.445 0.14 ;
    END
  END r_data_o[460]
  PIN r_data_o[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 39.235 0.07 39.305 ;
    END
  END r_data_o[461]
  PIN r_data_o[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 10.675 0.07 10.745 ;
    END
  END r_data_o[462]
  PIN r_data_o[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  85.705 0 85.845 0.14 ;
    END
  END r_data_o[463]
  PIN r_data_o[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  22.985 0 23.125 0.14 ;
    END
  END r_data_o[464]
  PIN r_data_o[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  133.865 81.61 134.005 81.75 ;
    END
  END r_data_o[465]
  PIN r_data_o[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  54.345 81.61 54.485 81.75 ;
    END
  END r_data_o[466]
  PIN r_data_o[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  63.305 0 63.445 0.14 ;
    END
  END r_data_o[467]
  PIN r_data_o[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 42.595 0.07 42.665 ;
    END
  END r_data_o[468]
  PIN r_data_o[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  47.625 0 47.765 0.14 ;
    END
  END r_data_o[469]
  PIN r_data_o[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  148.985 81.61 149.125 81.75 ;
    END
  END r_data_o[46]
  PIN r_data_o[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  151.225 0 151.365 0.14 ;
    END
  END r_data_o[470]
  PIN r_data_o[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 31.675 161.495 31.745 ;
    END
  END r_data_o[471]
  PIN r_data_o[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 15.715 161.495 15.785 ;
    END
  END r_data_o[472]
  PIN r_data_o[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 15.995 0.07 16.065 ;
    END
  END r_data_o[473]
  PIN r_data_o[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  26.345 81.61 26.485 81.75 ;
    END
  END r_data_o[474]
  PIN r_data_o[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 41.755 0.07 41.825 ;
    END
  END r_data_o[475]
  PIN r_data_o[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  49.865 81.61 50.005 81.75 ;
    END
  END r_data_o[476]
  PIN r_data_o[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 50.715 161.495 50.785 ;
    END
  END r_data_o[477]
  PIN r_data_o[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 15.995 161.495 16.065 ;
    END
  END r_data_o[478]
  PIN r_data_o[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 28.315 0.07 28.385 ;
    END
  END r_data_o[479]
  PIN r_data_o[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  157.385 81.61 157.525 81.75 ;
    END
  END r_data_o[47]
  PIN r_data_o[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  94.665 81.61 94.805 81.75 ;
    END
  END r_data_o[480]
  PIN r_data_o[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  136.665 0 136.805 0.14 ;
    END
  END r_data_o[481]
  PIN r_data_o[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  92.985 0 93.125 0.14 ;
    END
  END r_data_o[482]
  PIN r_data_o[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 50.435 0.07 50.505 ;
    END
  END r_data_o[483]
  PIN r_data_o[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  138.345 0 138.485 0.14 ;
    END
  END r_data_o[484]
  PIN r_data_o[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  99.145 81.61 99.285 81.75 ;
    END
  END r_data_o[485]
  PIN r_data_o[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 33.635 161.495 33.705 ;
    END
  END r_data_o[486]
  PIN r_data_o[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  154.025 0 154.165 0.14 ;
    END
  END r_data_o[487]
  PIN r_data_o[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  157.945 81.61 158.085 81.75 ;
    END
  END r_data_o[488]
  PIN r_data_o[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 42.315 0.07 42.385 ;
    END
  END r_data_o[489]
  PIN r_data_o[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  6.745 0 6.885 0.14 ;
    END
  END r_data_o[48]
  PIN r_data_o[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  33.065 81.61 33.205 81.75 ;
    END
  END r_data_o[490]
  PIN r_data_o[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  68.905 81.61 69.045 81.75 ;
    END
  END r_data_o[491]
  PIN r_data_o[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 35.875 161.495 35.945 ;
    END
  END r_data_o[492]
  PIN r_data_o[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.385 0 17.525 0.14 ;
    END
  END r_data_o[493]
  PIN r_data_o[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  151.785 0 151.925 0.14 ;
    END
  END r_data_o[494]
  PIN r_data_o[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  8.985 81.61 9.125 81.75 ;
    END
  END r_data_o[495]
  PIN r_data_o[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 4.795 161.495 4.865 ;
    END
  END r_data_o[496]
  PIN r_data_o[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 1.995 161.495 2.065 ;
    END
  END r_data_o[497]
  PIN r_data_o[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  133.865 0 134.005 0.14 ;
    END
  END r_data_o[498]
  PIN r_data_o[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 69.475 161.495 69.545 ;
    END
  END r_data_o[499]
  PIN r_data_o[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 29.715 0.07 29.785 ;
    END
  END r_data_o[49]
  PIN r_data_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  126.025 0 126.165 0.14 ;
    END
  END r_data_o[4]
  PIN r_data_o[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 65.555 0.07 65.625 ;
    END
  END r_data_o[500]
  PIN r_data_o[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 10.115 0.07 10.185 ;
    END
  END r_data_o[501]
  PIN r_data_o[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  49.305 81.61 49.445 81.75 ;
    END
  END r_data_o[502]
  PIN r_data_o[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  94.665 0 94.805 0.14 ;
    END
  END r_data_o[503]
  PIN r_data_o[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  74.505 81.61 74.645 81.75 ;
    END
  END r_data_o[504]
  PIN r_data_o[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 63.875 0.07 63.945 ;
    END
  END r_data_o[505]
  PIN r_data_o[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 32.795 161.495 32.865 ;
    END
  END r_data_o[506]
  PIN r_data_o[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 1.155 161.495 1.225 ;
    END
  END r_data_o[507]
  PIN r_data_o[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 41.195 161.495 41.265 ;
    END
  END r_data_o[508]
  PIN r_data_o[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 58.835 0.07 58.905 ;
    END
  END r_data_o[509]
  PIN r_data_o[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 79.555 161.495 79.625 ;
    END
  END r_data_o[50]
  PIN r_data_o[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  135.545 81.61 135.685 81.75 ;
    END
  END r_data_o[510]
  PIN r_data_o[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 28.035 0.07 28.105 ;
    END
  END r_data_o[511]
  PIN r_data_o[512]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  136.665 81.61 136.805 81.75 ;
    END
  END r_data_o[512]
  PIN r_data_o[513]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  113.145 81.61 113.285 81.75 ;
    END
  END r_data_o[513]
  PIN r_data_o[514]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  45.385 0 45.525 0.14 ;
    END
  END r_data_o[514]
  PIN r_data_o[515]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  90.185 0 90.325 0.14 ;
    END
  END r_data_o[515]
  PIN r_data_o[516]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  140.585 81.61 140.725 81.75 ;
    END
  END r_data_o[516]
  PIN r_data_o[517]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.345 81.61 12.485 81.75 ;
    END
  END r_data_o[517]
  PIN r_data_o[518]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  128.825 0 128.965 0.14 ;
    END
  END r_data_o[518]
  PIN r_data_o[519]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  89.625 81.61 89.765 81.75 ;
    END
  END r_data_o[519]
  PIN r_data_o[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  25.785 0 25.925 0.14 ;
    END
  END r_data_o[51]
  PIN r_data_o[520]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  5.065 0 5.205 0.14 ;
    END
  END r_data_o[520]
  PIN r_data_o[521]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  124.905 0 125.045 0.14 ;
    END
  END r_data_o[521]
  PIN r_data_o[522]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  46.505 0 46.645 0.14 ;
    END
  END r_data_o[522]
  PIN r_data_o[523]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 13.475 161.495 13.545 ;
    END
  END r_data_o[523]
  PIN r_data_o[524]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 50.155 161.495 50.225 ;
    END
  END r_data_o[524]
  PIN r_data_o[525]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 33.915 161.495 33.985 ;
    END
  END r_data_o[525]
  PIN r_data_o[526]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 76.195 0.07 76.265 ;
    END
  END r_data_o[526]
  PIN r_data_o[527]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  11.225 0 11.365 0.14 ;
    END
  END r_data_o[527]
  PIN r_data_o[528]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  129.945 81.61 130.085 81.75 ;
    END
  END r_data_o[528]
  PIN r_data_o[529]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 58.275 0.07 58.345 ;
    END
  END r_data_o[529]
  PIN r_data_o[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  6.185 81.61 6.325 81.75 ;
    END
  END r_data_o[52]
  PIN r_data_o[530]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.385 0 31.525 0.14 ;
    END
  END r_data_o[530]
  PIN r_data_o[531]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  92.425 0 92.565 0.14 ;
    END
  END r_data_o[531]
  PIN r_data_o[532]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  70.025 81.61 70.165 81.75 ;
    END
  END r_data_o[532]
  PIN r_data_o[533]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  33.065 0 33.205 0.14 ;
    END
  END r_data_o[533]
  PIN r_data_o[534]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 22.995 161.495 23.065 ;
    END
  END r_data_o[534]
  PIN r_data_o[535]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 26.355 0.07 26.425 ;
    END
  END r_data_o[535]
  PIN r_data_o[536]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  97.465 0 97.605 0.14 ;
    END
  END r_data_o[536]
  PIN r_data_o[537]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 69.755 161.495 69.825 ;
    END
  END r_data_o[537]
  PIN r_data_o[538]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  67.785 0 67.925 0.14 ;
    END
  END r_data_o[538]
  PIN r_data_o[539]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 6.475 0.07 6.545 ;
    END
  END r_data_o[539]
  PIN r_data_o[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  115.385 0 115.525 0.14 ;
    END
  END r_data_o[53]
  PIN r_data_o[540]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 20.755 161.495 20.825 ;
    END
  END r_data_o[540]
  PIN r_data_o[541]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 76.755 161.495 76.825 ;
    END
  END r_data_o[541]
  PIN r_data_o[542]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 75.635 0.07 75.705 ;
    END
  END r_data_o[542]
  PIN r_data_o[543]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 65.835 0.07 65.905 ;
    END
  END r_data_o[543]
  PIN r_data_o[544]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 11.515 161.495 11.585 ;
    END
  END r_data_o[544]
  PIN r_data_o[545]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 22.715 161.495 22.785 ;
    END
  END r_data_o[545]
  PIN r_data_o[546]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  57.705 81.61 57.845 81.75 ;
    END
  END r_data_o[546]
  PIN r_data_o[547]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 53.515 161.495 53.585 ;
    END
  END r_data_o[547]
  PIN r_data_o[548]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 9.555 161.495 9.625 ;
    END
  END r_data_o[548]
  PIN r_data_o[549]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  78.425 0 78.565 0.14 ;
    END
  END r_data_o[549]
  PIN r_data_o[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 51.555 161.495 51.625 ;
    END
  END r_data_o[54]
  PIN r_data_o[550]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 13.195 161.495 13.265 ;
    END
  END r_data_o[550]
  PIN r_data_o[551]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 32.235 0.07 32.305 ;
    END
  END r_data_o[551]
  PIN r_data_o[552]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  24.665 81.61 24.805 81.75 ;
    END
  END r_data_o[552]
  PIN r_data_o[553]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  26.905 0 27.045 0.14 ;
    END
  END r_data_o[553]
  PIN r_data_o[554]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 35.035 0.07 35.105 ;
    END
  END r_data_o[554]
  PIN r_data_o[555]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  68.345 0 68.485 0.14 ;
    END
  END r_data_o[555]
  PIN r_data_o[556]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  82.905 81.61 83.045 81.75 ;
    END
  END r_data_o[556]
  PIN r_data_o[557]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  126.585 0 126.725 0.14 ;
    END
  END r_data_o[557]
  PIN r_data_o[558]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  44.825 0 44.965 0.14 ;
    END
  END r_data_o[558]
  PIN r_data_o[559]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  152.905 81.61 153.045 81.75 ;
    END
  END r_data_o[559]
  PIN r_data_o[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 80.675 161.495 80.745 ;
    END
  END r_data_o[55]
  PIN r_data_o[560]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  117.065 81.61 117.205 81.75 ;
    END
  END r_data_o[560]
  PIN r_data_o[561]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.395 0.07 31.465 ;
    END
  END r_data_o[561]
  PIN r_data_o[562]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  126.025 81.61 126.165 81.75 ;
    END
  END r_data_o[562]
  PIN r_data_o[563]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  129.385 81.61 129.525 81.75 ;
    END
  END r_data_o[563]
  PIN r_data_o[564]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 42.875 0.07 42.945 ;
    END
  END r_data_o[564]
  PIN r_data_o[565]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  140.025 81.61 140.165 81.75 ;
    END
  END r_data_o[565]
  PIN r_data_o[566]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 70.315 161.495 70.385 ;
    END
  END r_data_o[566]
  PIN r_data_o[567]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  44.265 81.61 44.405 81.75 ;
    END
  END r_data_o[567]
  PIN r_data_o[568]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 64.995 0.07 65.065 ;
    END
  END r_data_o[568]
  PIN r_data_o[569]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.945 81.61 32.085 81.75 ;
    END
  END r_data_o[569]
  PIN r_data_o[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  73.945 0 74.085 0.14 ;
    END
  END r_data_o[56]
  PIN r_data_o[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  151.225 81.61 151.365 81.75 ;
    END
  END r_data_o[57]
  PIN r_data_o[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 70.875 161.495 70.945 ;
    END
  END r_data_o[58]
  PIN r_data_o[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  129.385 0 129.525 0.14 ;
    END
  END r_data_o[59]
  PIN r_data_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  3.385 81.61 3.525 81.75 ;
    END
  END r_data_o[5]
  PIN r_data_o[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 37.835 0.07 37.905 ;
    END
  END r_data_o[60]
  PIN r_data_o[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  118.185 0 118.325 0.14 ;
    END
  END r_data_o[61]
  PIN r_data_o[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 38.395 161.495 38.465 ;
    END
  END r_data_o[62]
  PIN r_data_o[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 77.875 161.495 77.945 ;
    END
  END r_data_o[63]
  PIN r_data_o[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  96.345 0 96.485 0.14 ;
    END
  END r_data_o[64]
  PIN r_data_o[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 26.915 161.495 26.985 ;
    END
  END r_data_o[65]
  PIN r_data_o[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  154.585 0 154.725 0.14 ;
    END
  END r_data_o[66]
  PIN r_data_o[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  154.585 81.61 154.725 81.75 ;
    END
  END r_data_o[67]
  PIN r_data_o[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 66.955 161.495 67.025 ;
    END
  END r_data_o[68]
  PIN r_data_o[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  53.225 81.61 53.365 81.75 ;
    END
  END r_data_o[69]
  PIN r_data_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 29.715 161.495 29.785 ;
    END
  END r_data_o[6]
  PIN r_data_o[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 6.195 0.07 6.265 ;
    END
  END r_data_o[70]
  PIN r_data_o[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 16.835 161.495 16.905 ;
    END
  END r_data_o[71]
  PIN r_data_o[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 26.355 161.495 26.425 ;
    END
  END r_data_o[72]
  PIN r_data_o[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 2.555 161.495 2.625 ;
    END
  END r_data_o[73]
  PIN r_data_o[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  133.305 81.61 133.445 81.75 ;
    END
  END r_data_o[74]
  PIN r_data_o[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 1.435 161.495 1.505 ;
    END
  END r_data_o[75]
  PIN r_data_o[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 74.795 0.07 74.865 ;
    END
  END r_data_o[76]
  PIN r_data_o[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  6.745 81.61 6.885 81.75 ;
    END
  END r_data_o[77]
  PIN r_data_o[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 49.315 161.495 49.385 ;
    END
  END r_data_o[78]
  PIN r_data_o[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 33.355 0.07 33.425 ;
    END
  END r_data_o[79]
  PIN r_data_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  141.145 0 141.285 0.14 ;
    END
  END r_data_o[7]
  PIN r_data_o[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 16.275 161.495 16.345 ;
    END
  END r_data_o[80]
  PIN r_data_o[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  72.825 81.61 72.965 81.75 ;
    END
  END r_data_o[81]
  PIN r_data_o[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  66.665 81.61 66.805 81.75 ;
    END
  END r_data_o[82]
  PIN r_data_o[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  84.585 0 84.725 0.14 ;
    END
  END r_data_o[83]
  PIN r_data_o[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 39.795 0.07 39.865 ;
    END
  END r_data_o[84]
  PIN r_data_o[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 49.035 161.495 49.105 ;
    END
  END r_data_o[85]
  PIN r_data_o[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 1.715 161.495 1.785 ;
    END
  END r_data_o[86]
  PIN r_data_o[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.185 81.61 34.325 81.75 ;
    END
  END r_data_o[87]
  PIN r_data_o[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 18.795 0.07 18.865 ;
    END
  END r_data_o[88]
  PIN r_data_o[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 38.115 0.07 38.185 ;
    END
  END r_data_o[89]
  PIN r_data_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  113.145 0 113.285 0.14 ;
    END
  END r_data_o[8]
  PIN r_data_o[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 66.395 0.07 66.465 ;
    END
  END r_data_o[90]
  PIN r_data_o[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  13.465 81.61 13.605 81.75 ;
    END
  END r_data_o[91]
  PIN r_data_o[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 78.155 161.495 78.225 ;
    END
  END r_data_o[92]
  PIN r_data_o[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.345 0 12.485 0.14 ;
    END
  END r_data_o[93]
  PIN r_data_o[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  79.545 0 79.685 0.14 ;
    END
  END r_data_o[94]
  PIN r_data_o[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.035 0.07 7.105 ;
    END
  END r_data_o[95]
  PIN r_data_o[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 77.315 0.07 77.385 ;
    END
  END r_data_o[96]
  PIN r_data_o[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 14.315 161.495 14.385 ;
    END
  END r_data_o[97]
  PIN r_data_o[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  29.705 81.61 29.845 81.75 ;
    END
  END r_data_o[98]
  PIN r_data_o[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  43.705 81.61 43.845 81.75 ;
    END
  END r_data_o[99]
  PIN r_data_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  4.505 81.61 4.645 81.75 ;
    END
  END r_data_o[9]
  PIN r_v_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  124.345 81.61 124.485 81.75 ;
    END
  END r_v_i
  PIN w_addr_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  43.145 81.61 43.285 81.75 ;
    END
  END w_addr_i
  PIN w_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  150.105 0 150.245 0.14 ;
    END
  END w_clk_i
  PIN w_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  105.865 0 106.005 0.14 ;
    END
  END w_data_i[0]
  PIN w_data_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  11.785 0 11.925 0.14 ;
    END
  END w_data_i[100]
  PIN w_data_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  20.185 81.61 20.325 81.75 ;
    END
  END w_data_i[101]
  PIN w_data_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 5.355 0.07 5.425 ;
    END
  END w_data_i[102]
  PIN w_data_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  143.385 81.61 143.525 81.75 ;
    END
  END w_data_i[103]
  PIN w_data_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  30.825 0 30.965 0.14 ;
    END
  END w_data_i[104]
  PIN w_data_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  114.825 81.61 114.965 81.75 ;
    END
  END w_data_i[105]
  PIN w_data_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 27.475 0.07 27.545 ;
    END
  END w_data_i[106]
  PIN w_data_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  56.025 81.61 56.165 81.75 ;
    END
  END w_data_i[107]
  PIN w_data_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  120.985 81.61 121.125 81.75 ;
    END
  END w_data_i[108]
  PIN w_data_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 65.555 161.495 65.625 ;
    END
  END w_data_i[109]
  PIN w_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  85.705 81.61 85.845 81.75 ;
    END
  END w_data_i[10]
  PIN w_data_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  23.545 81.61 23.685 81.75 ;
    END
  END w_data_i[110]
  PIN w_data_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 51.275 161.495 51.345 ;
    END
  END w_data_i[111]
  PIN w_data_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 59.675 0.07 59.745 ;
    END
  END w_data_i[112]
  PIN w_data_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 25.235 0.07 25.305 ;
    END
  END w_data_i[113]
  PIN w_data_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  23.545 0 23.685 0.14 ;
    END
  END w_data_i[114]
  PIN w_data_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  131.625 81.61 131.765 81.75 ;
    END
  END w_data_i[115]
  PIN w_data_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 51.275 0.07 51.345 ;
    END
  END w_data_i[116]
  PIN w_data_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 53.235 161.495 53.305 ;
    END
  END w_data_i[117]
  PIN w_data_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 24.955 161.495 25.025 ;
    END
  END w_data_i[118]
  PIN w_data_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  55.465 81.61 55.605 81.75 ;
    END
  END w_data_i[119]
  PIN w_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 22.995 0.07 23.065 ;
    END
  END w_data_i[11]
  PIN w_data_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 5.915 161.495 5.985 ;
    END
  END w_data_i[120]
  PIN w_data_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  119.865 81.61 120.005 81.75 ;
    END
  END w_data_i[121]
  PIN w_data_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  59.945 81.61 60.085 81.75 ;
    END
  END w_data_i[122]
  PIN w_data_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 23.275 161.495 23.345 ;
    END
  END w_data_i[123]
  PIN w_data_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  137.785 81.61 137.925 81.75 ;
    END
  END w_data_i[124]
  PIN w_data_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.635 0.07 12.705 ;
    END
  END w_data_i[125]
  PIN w_data_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 67.515 0.07 67.585 ;
    END
  END w_data_i[126]
  PIN w_data_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  142.265 0 142.405 0.14 ;
    END
  END w_data_i[127]
  PIN w_data_i[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 57.715 161.495 57.785 ;
    END
  END w_data_i[128]
  PIN w_data_i[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  100.825 0 100.965 0.14 ;
    END
  END w_data_i[129]
  PIN w_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  100.265 0 100.405 0.14 ;
    END
  END w_data_i[12]
  PIN w_data_i[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  61.065 81.61 61.205 81.75 ;
    END
  END w_data_i[130]
  PIN w_data_i[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  123.225 0 123.365 0.14 ;
    END
  END w_data_i[131]
  PIN w_data_i[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 41.755 161.495 41.825 ;
    END
  END w_data_i[132]
  PIN w_data_i[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 73.955 0.07 74.025 ;
    END
  END w_data_i[133]
  PIN w_data_i[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  47.065 0 47.205 0.14 ;
    END
  END w_data_i[134]
  PIN w_data_i[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  69.465 81.61 69.605 81.75 ;
    END
  END w_data_i[135]
  PIN w_data_i[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  20.745 81.61 20.885 81.75 ;
    END
  END w_data_i[136]
  PIN w_data_i[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 48.195 161.495 48.265 ;
    END
  END w_data_i[137]
  PIN w_data_i[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 1.155 0.07 1.225 ;
    END
  END w_data_i[138]
  PIN w_data_i[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  45.945 81.61 46.085 81.75 ;
    END
  END w_data_i[139]
  PIN w_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  102.505 0 102.645 0.14 ;
    END
  END w_data_i[13]
  PIN w_data_i[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 68.915 0.07 68.985 ;
    END
  END w_data_i[140]
  PIN w_data_i[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  88.505 0 88.645 0.14 ;
    END
  END w_data_i[141]
  PIN w_data_i[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  49.305 0 49.445 0.14 ;
    END
  END w_data_i[142]
  PIN w_data_i[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  125.465 0 125.605 0.14 ;
    END
  END w_data_i[143]
  PIN w_data_i[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 19.635 0.07 19.705 ;
    END
  END w_data_i[144]
  PIN w_data_i[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 37.835 161.495 37.905 ;
    END
  END w_data_i[145]
  PIN w_data_i[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  105.305 81.61 105.445 81.75 ;
    END
  END w_data_i[146]
  PIN w_data_i[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 59.395 0.07 59.465 ;
    END
  END w_data_i[147]
  PIN w_data_i[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.745 0 34.885 0.14 ;
    END
  END w_data_i[148]
  PIN w_data_i[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  25.225 0 25.365 0.14 ;
    END
  END w_data_i[149]
  PIN w_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 21.035 161.495 21.105 ;
    END
  END w_data_i[14]
  PIN w_data_i[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  94.105 81.61 94.245 81.75 ;
    END
  END w_data_i[150]
  PIN w_data_i[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  22.985 81.61 23.125 81.75 ;
    END
  END w_data_i[151]
  PIN w_data_i[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 70.035 161.495 70.105 ;
    END
  END w_data_i[152]
  PIN w_data_i[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  149.545 81.61 149.685 81.75 ;
    END
  END w_data_i[153]
  PIN w_data_i[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  140.585 0 140.725 0.14 ;
    END
  END w_data_i[154]
  PIN w_data_i[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 33.635 0.07 33.705 ;
    END
  END w_data_i[155]
  PIN w_data_i[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 29.155 0.07 29.225 ;
    END
  END w_data_i[156]
  PIN w_data_i[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  40.905 81.61 41.045 81.75 ;
    END
  END w_data_i[157]
  PIN w_data_i[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 7.315 161.495 7.385 ;
    END
  END w_data_i[158]
  PIN w_data_i[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 1.995 0.07 2.065 ;
    END
  END w_data_i[159]
  PIN w_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  96.905 0 97.045 0.14 ;
    END
  END w_data_i[15]
  PIN w_data_i[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  30.825 81.61 30.965 81.75 ;
    END
  END w_data_i[160]
  PIN w_data_i[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  25.785 81.61 25.925 81.75 ;
    END
  END w_data_i[161]
  PIN w_data_i[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  139.465 0 139.605 0.14 ;
    END
  END w_data_i[162]
  PIN w_data_i[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.385 81.61 17.525 81.75 ;
    END
  END w_data_i[163]
  PIN w_data_i[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  106.985 0 107.125 0.14 ;
    END
  END w_data_i[164]
  PIN w_data_i[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  27.465 0 27.605 0.14 ;
    END
  END w_data_i[165]
  PIN w_data_i[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 35.315 0.07 35.385 ;
    END
  END w_data_i[166]
  PIN w_data_i[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  125.465 81.61 125.605 81.75 ;
    END
  END w_data_i[167]
  PIN w_data_i[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  114.265 81.61 114.405 81.75 ;
    END
  END w_data_i[168]
  PIN w_data_i[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 24.675 161.495 24.745 ;
    END
  END w_data_i[169]
  PIN w_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  128.825 81.61 128.965 81.75 ;
    END
  END w_data_i[16]
  PIN w_data_i[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 21.315 161.495 21.385 ;
    END
  END w_data_i[170]
  PIN w_data_i[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 28.875 0.07 28.945 ;
    END
  END w_data_i[171]
  PIN w_data_i[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  121.545 0 121.685 0.14 ;
    END
  END w_data_i[172]
  PIN w_data_i[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  141.145 81.61 141.285 81.75 ;
    END
  END w_data_i[173]
  PIN w_data_i[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  62.185 81.61 62.325 81.75 ;
    END
  END w_data_i[174]
  PIN w_data_i[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  6.185 0 6.325 0.14 ;
    END
  END w_data_i[175]
  PIN w_data_i[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 58.275 161.495 58.345 ;
    END
  END w_data_i[176]
  PIN w_data_i[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 63.595 0.07 63.665 ;
    END
  END w_data_i[177]
  PIN w_data_i[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  36.985 81.61 37.125 81.75 ;
    END
  END w_data_i[178]
  PIN w_data_i[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  142.825 81.61 142.965 81.75 ;
    END
  END w_data_i[179]
  PIN w_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  91.305 81.61 91.445 81.75 ;
    END
  END w_data_i[17]
  PIN w_data_i[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  64.985 81.61 65.125 81.75 ;
    END
  END w_data_i[180]
  PIN w_data_i[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 7.875 161.495 7.945 ;
    END
  END w_data_i[181]
  PIN w_data_i[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  131.065 81.61 131.205 81.75 ;
    END
  END w_data_i[182]
  PIN w_data_i[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  63.865 81.61 64.005 81.75 ;
    END
  END w_data_i[183]
  PIN w_data_i[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  66.665 0 66.805 0.14 ;
    END
  END w_data_i[184]
  PIN w_data_i[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 56.875 0.07 56.945 ;
    END
  END w_data_i[185]
  PIN w_data_i[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 41.475 161.495 41.545 ;
    END
  END w_data_i[186]
  PIN w_data_i[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 64.715 161.495 64.785 ;
    END
  END w_data_i[187]
  PIN w_data_i[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  9.545 0 9.685 0.14 ;
    END
  END w_data_i[188]
  PIN w_data_i[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 28.035 161.495 28.105 ;
    END
  END w_data_i[189]
  PIN w_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 30.555 0.07 30.625 ;
    END
  END w_data_i[18]
  PIN w_data_i[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  95.225 81.61 95.365 81.75 ;
    END
  END w_data_i[190]
  PIN w_data_i[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 57.155 161.495 57.225 ;
    END
  END w_data_i[191]
  PIN w_data_i[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  87.385 0 87.525 0.14 ;
    END
  END w_data_i[192]
  PIN w_data_i[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  74.505 0 74.645 0.14 ;
    END
  END w_data_i[193]
  PIN w_data_i[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  153.465 81.61 153.605 81.75 ;
    END
  END w_data_i[194]
  PIN w_data_i[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 33.915 0.07 33.985 ;
    END
  END w_data_i[195]
  PIN w_data_i[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 47.915 161.495 47.985 ;
    END
  END w_data_i[196]
  PIN w_data_i[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 30.555 161.495 30.625 ;
    END
  END w_data_i[197]
  PIN w_data_i[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 43.715 161.495 43.785 ;
    END
  END w_data_i[198]
  PIN w_data_i[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 16.555 161.495 16.625 ;
    END
  END w_data_i[199]
  PIN w_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  134.425 0 134.565 0.14 ;
    END
  END w_data_i[19]
  PIN w_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 73.115 161.495 73.185 ;
    END
  END w_data_i[1]
  PIN w_data_i[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 3.955 161.495 4.025 ;
    END
  END w_data_i[200]
  PIN w_data_i[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 42.035 161.495 42.105 ;
    END
  END w_data_i[201]
  PIN w_data_i[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  132.185 81.61 132.325 81.75 ;
    END
  END w_data_i[202]
  PIN w_data_i[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  137.225 81.61 137.365 81.75 ;
    END
  END w_data_i[203]
  PIN w_data_i[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 14.595 161.495 14.665 ;
    END
  END w_data_i[204]
  PIN w_data_i[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  152.905 0 153.045 0.14 ;
    END
  END w_data_i[205]
  PIN w_data_i[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  101.945 81.61 102.085 81.75 ;
    END
  END w_data_i[206]
  PIN w_data_i[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  103.625 81.61 103.765 81.75 ;
    END
  END w_data_i[207]
  PIN w_data_i[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  39.225 81.61 39.365 81.75 ;
    END
  END w_data_i[208]
  PIN w_data_i[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  81.225 81.61 81.365 81.75 ;
    END
  END w_data_i[209]
  PIN w_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  98.025 0 98.165 0.14 ;
    END
  END w_data_i[20]
  PIN w_data_i[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 71.995 0.07 72.065 ;
    END
  END w_data_i[210]
  PIN w_data_i[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 44.835 161.495 44.905 ;
    END
  END w_data_i[211]
  PIN w_data_i[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 22.435 0.07 22.505 ;
    END
  END w_data_i[212]
  PIN w_data_i[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 20.195 161.495 20.265 ;
    END
  END w_data_i[213]
  PIN w_data_i[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 4.235 0.07 4.305 ;
    END
  END w_data_i[214]
  PIN w_data_i[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 27.195 161.495 27.265 ;
    END
  END w_data_i[215]
  PIN w_data_i[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 32.515 161.495 32.585 ;
    END
  END w_data_i[216]
  PIN w_data_i[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 79.835 0.07 79.905 ;
    END
  END w_data_i[217]
  PIN w_data_i[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 50.435 161.495 50.505 ;
    END
  END w_data_i[218]
  PIN w_data_i[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 63.035 161.495 63.105 ;
    END
  END w_data_i[219]
  PIN w_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 43.715 0.07 43.785 ;
    END
  END w_data_i[21]
  PIN w_data_i[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 68.075 161.495 68.145 ;
    END
  END w_data_i[220]
  PIN w_data_i[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 49.595 161.495 49.665 ;
    END
  END w_data_i[221]
  PIN w_data_i[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  146.185 0 146.325 0.14 ;
    END
  END w_data_i[222]
  PIN w_data_i[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 39.515 0.07 39.585 ;
    END
  END w_data_i[223]
  PIN w_data_i[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  1.145 81.61 1.285 81.75 ;
    END
  END w_data_i[224]
  PIN w_data_i[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  130.505 0 130.645 0.14 ;
    END
  END w_data_i[225]
  PIN w_data_i[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 19.355 161.495 19.425 ;
    END
  END w_data_i[226]
  PIN w_data_i[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  95.225 0 95.365 0.14 ;
    END
  END w_data_i[227]
  PIN w_data_i[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.305 0 7.445 0.14 ;
    END
  END w_data_i[228]
  PIN w_data_i[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 63.595 161.495 63.665 ;
    END
  END w_data_i[229]
  PIN w_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  71.145 0 71.285 0.14 ;
    END
  END w_data_i[22]
  PIN w_data_i[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 5.635 0.07 5.705 ;
    END
  END w_data_i[230]
  PIN w_data_i[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  80.105 81.61 80.245 81.75 ;
    END
  END w_data_i[231]
  PIN w_data_i[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 22.715 0.07 22.785 ;
    END
  END w_data_i[232]
  PIN w_data_i[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 46.795 0.07 46.865 ;
    END
  END w_data_i[233]
  PIN w_data_i[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 14.315 0.07 14.385 ;
    END
  END w_data_i[234]
  PIN w_data_i[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 19.075 161.495 19.145 ;
    END
  END w_data_i[235]
  PIN w_data_i[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  50.425 81.61 50.565 81.75 ;
    END
  END w_data_i[236]
  PIN w_data_i[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  124.345 0 124.485 0.14 ;
    END
  END w_data_i[237]
  PIN w_data_i[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  66.105 0 66.245 0.14 ;
    END
  END w_data_i[238]
  PIN w_data_i[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  115.945 0 116.085 0.14 ;
    END
  END w_data_i[239]
  PIN w_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  2.265 0 2.405 0.14 ;
    END
  END w_data_i[23]
  PIN w_data_i[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  83.465 81.61 83.605 81.75 ;
    END
  END w_data_i[240]
  PIN w_data_i[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 56.315 161.495 56.385 ;
    END
  END w_data_i[241]
  PIN w_data_i[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  95.785 81.61 95.925 81.75 ;
    END
  END w_data_i[242]
  PIN w_data_i[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  42.025 0 42.165 0.14 ;
    END
  END w_data_i[243]
  PIN w_data_i[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 25.515 0.07 25.585 ;
    END
  END w_data_i[244]
  PIN w_data_i[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 2.275 0.07 2.345 ;
    END
  END w_data_i[245]
  PIN w_data_i[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 40.075 161.495 40.145 ;
    END
  END w_data_i[246]
  PIN w_data_i[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.875 0.07 7.945 ;
    END
  END w_data_i[247]
  PIN w_data_i[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.585 81.61 14.725 81.75 ;
    END
  END w_data_i[248]
  PIN w_data_i[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  19.065 81.61 19.205 81.75 ;
    END
  END w_data_i[249]
  PIN w_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 44.275 0.07 44.345 ;
    END
  END w_data_i[24]
  PIN w_data_i[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  67.225 0 67.365 0.14 ;
    END
  END w_data_i[250]
  PIN w_data_i[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  92.425 81.61 92.565 81.75 ;
    END
  END w_data_i[251]
  PIN w_data_i[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 47.355 0.07 47.425 ;
    END
  END w_data_i[252]
  PIN w_data_i[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  16.265 81.61 16.405 81.75 ;
    END
  END w_data_i[253]
  PIN w_data_i[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 58.555 0.07 58.625 ;
    END
  END w_data_i[254]
  PIN w_data_i[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  110.345 81.61 110.485 81.75 ;
    END
  END w_data_i[255]
  PIN w_data_i[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 10.395 0.07 10.465 ;
    END
  END w_data_i[256]
  PIN w_data_i[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 5.075 161.495 5.145 ;
    END
  END w_data_i[257]
  PIN w_data_i[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  109.225 81.61 109.365 81.75 ;
    END
  END w_data_i[258]
  PIN w_data_i[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 44.835 0.07 44.905 ;
    END
  END w_data_i[259]
  PIN w_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  104.185 81.61 104.325 81.75 ;
    END
  END w_data_i[25]
  PIN w_data_i[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  124.905 81.61 125.045 81.75 ;
    END
  END w_data_i[260]
  PIN w_data_i[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 27.195 0.07 27.265 ;
    END
  END w_data_i[261]
  PIN w_data_i[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 68.355 161.495 68.425 ;
    END
  END w_data_i[262]
  PIN w_data_i[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  148.425 0 148.565 0.14 ;
    END
  END w_data_i[263]
  PIN w_data_i[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  118.745 0 118.885 0.14 ;
    END
  END w_data_i[264]
  PIN w_data_i[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  143.945 0 144.085 0.14 ;
    END
  END w_data_i[265]
  PIN w_data_i[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  80.665 0 80.805 0.14 ;
    END
  END w_data_i[266]
  PIN w_data_i[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 55.195 161.495 55.265 ;
    END
  END w_data_i[267]
  PIN w_data_i[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  105.865 81.61 106.005 81.75 ;
    END
  END w_data_i[268]
  PIN w_data_i[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  97.465 81.61 97.605 81.75 ;
    END
  END w_data_i[269]
  PIN w_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 39.515 161.495 39.585 ;
    END
  END w_data_i[26]
  PIN w_data_i[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  98.025 81.61 98.165 81.75 ;
    END
  END w_data_i[270]
  PIN w_data_i[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 53.515 0.07 53.585 ;
    END
  END w_data_i[271]
  PIN w_data_i[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 61.915 0.07 61.985 ;
    END
  END w_data_i[272]
  PIN w_data_i[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  53.785 81.61 53.925 81.75 ;
    END
  END w_data_i[273]
  PIN w_data_i[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  104.185 0 104.325 0.14 ;
    END
  END w_data_i[274]
  PIN w_data_i[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  46.505 81.61 46.645 81.75 ;
    END
  END w_data_i[275]
  PIN w_data_i[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 55.195 0.07 55.265 ;
    END
  END w_data_i[276]
  PIN w_data_i[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 34.475 0.07 34.545 ;
    END
  END w_data_i[277]
  PIN w_data_i[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 51.555 0.07 51.625 ;
    END
  END w_data_i[278]
  PIN w_data_i[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  56.585 81.61 56.725 81.75 ;
    END
  END w_data_i[279]
  PIN w_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  127.705 81.61 127.845 81.75 ;
    END
  END w_data_i[27]
  PIN w_data_i[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  76.185 0 76.325 0.14 ;
    END
  END w_data_i[280]
  PIN w_data_i[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 63.875 161.495 63.945 ;
    END
  END w_data_i[281]
  PIN w_data_i[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.385 81.61 31.525 81.75 ;
    END
  END w_data_i[282]
  PIN w_data_i[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.945 81.61 18.085 81.75 ;
    END
  END w_data_i[283]
  PIN w_data_i[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 72.275 161.495 72.345 ;
    END
  END w_data_i[284]
  PIN w_data_i[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  98.585 81.61 98.725 81.75 ;
    END
  END w_data_i[285]
  PIN w_data_i[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 38.675 161.495 38.745 ;
    END
  END w_data_i[286]
  PIN w_data_i[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  76.745 81.61 76.885 81.75 ;
    END
  END w_data_i[287]
  PIN w_data_i[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  91.865 0 92.005 0.14 ;
    END
  END w_data_i[288]
  PIN w_data_i[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  49.865 0 50.005 0.14 ;
    END
  END w_data_i[289]
  PIN w_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  158.505 81.61 158.645 81.75 ;
    END
  END w_data_i[28]
  PIN w_data_i[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 62.475 0.07 62.545 ;
    END
  END w_data_i[290]
  PIN w_data_i[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 69.195 161.495 69.265 ;
    END
  END w_data_i[291]
  PIN w_data_i[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  61.065 0 61.205 0.14 ;
    END
  END w_data_i[292]
  PIN w_data_i[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  112.025 81.61 112.165 81.75 ;
    END
  END w_data_i[293]
  PIN w_data_i[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  67.225 81.61 67.365 81.75 ;
    END
  END w_data_i[294]
  PIN w_data_i[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 35.035 161.495 35.105 ;
    END
  END w_data_i[295]
  PIN w_data_i[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 6.195 161.495 6.265 ;
    END
  END w_data_i[296]
  PIN w_data_i[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 8.715 161.495 8.785 ;
    END
  END w_data_i[297]
  PIN w_data_i[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 73.955 161.495 74.025 ;
    END
  END w_data_i[298]
  PIN w_data_i[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  63.305 81.61 63.445 81.75 ;
    END
  END w_data_i[299]
  PIN w_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  77.865 0 78.005 0.14 ;
    END
  END w_data_i[29]
  PIN w_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  43.145 0 43.285 0.14 ;
    END
  END w_data_i[2]
  PIN w_data_i[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 64.435 161.495 64.505 ;
    END
  END w_data_i[300]
  PIN w_data_i[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  156.265 0 156.405 0.14 ;
    END
  END w_data_i[301]
  PIN w_data_i[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  101.945 0 102.085 0.14 ;
    END
  END w_data_i[302]
  PIN w_data_i[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  118.745 81.61 118.885 81.75 ;
    END
  END w_data_i[303]
  PIN w_data_i[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 35.315 161.495 35.385 ;
    END
  END w_data_i[304]
  PIN w_data_i[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 80.395 161.495 80.465 ;
    END
  END w_data_i[305]
  PIN w_data_i[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.865 0 8.005 0.14 ;
    END
  END w_data_i[306]
  PIN w_data_i[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 3.675 0.07 3.745 ;
    END
  END w_data_i[307]
  PIN w_data_i[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 73.395 161.495 73.465 ;
    END
  END w_data_i[308]
  PIN w_data_i[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  147.865 0 148.005 0.14 ;
    END
  END w_data_i[309]
  PIN w_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 54.075 161.495 54.145 ;
    END
  END w_data_i[30]
  PIN w_data_i[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  92.985 81.61 93.125 81.75 ;
    END
  END w_data_i[310]
  PIN w_data_i[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  19.065 0 19.205 0.14 ;
    END
  END w_data_i[311]
  PIN w_data_i[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 78.435 161.495 78.505 ;
    END
  END w_data_i[312]
  PIN w_data_i[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  85.145 0 85.285 0.14 ;
    END
  END w_data_i[313]
  PIN w_data_i[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 36.155 161.495 36.225 ;
    END
  END w_data_i[314]
  PIN w_data_i[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  146.745 0 146.885 0.14 ;
    END
  END w_data_i[315]
  PIN w_data_i[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.665 81.61 10.805 81.75 ;
    END
  END w_data_i[316]
  PIN w_data_i[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  100.265 81.61 100.405 81.75 ;
    END
  END w_data_i[317]
  PIN w_data_i[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  116.505 81.61 116.645 81.75 ;
    END
  END w_data_i[318]
  PIN w_data_i[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 43.995 0.07 44.065 ;
    END
  END w_data_i[319]
  PIN w_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  107.545 81.61 107.685 81.75 ;
    END
  END w_data_i[31]
  PIN w_data_i[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 43.435 161.495 43.505 ;
    END
  END w_data_i[320]
  PIN w_data_i[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.035 0.07 21.105 ;
    END
  END w_data_i[321]
  PIN w_data_i[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  3.945 81.61 4.085 81.75 ;
    END
  END w_data_i[322]
  PIN w_data_i[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 29.435 0.07 29.505 ;
    END
  END w_data_i[323]
  PIN w_data_i[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 66.395 161.495 66.465 ;
    END
  END w_data_i[324]
  PIN w_data_i[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 28.875 161.495 28.945 ;
    END
  END w_data_i[325]
  PIN w_data_i[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 5.355 161.495 5.425 ;
    END
  END w_data_i[326]
  PIN w_data_i[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  109.785 81.61 109.925 81.75 ;
    END
  END w_data_i[327]
  PIN w_data_i[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  144.505 81.61 144.645 81.75 ;
    END
  END w_data_i[328]
  PIN w_data_i[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  112.585 0 112.725 0.14 ;
    END
  END w_data_i[329]
  PIN w_data_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  110.905 0 111.045 0.14 ;
    END
  END w_data_i[32]
  PIN w_data_i[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 6.475 161.495 6.545 ;
    END
  END w_data_i[330]
  PIN w_data_i[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  127.145 81.61 127.285 81.75 ;
    END
  END w_data_i[331]
  PIN w_data_i[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  38.105 0 38.245 0.14 ;
    END
  END w_data_i[332]
  PIN w_data_i[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 77.315 161.495 77.385 ;
    END
  END w_data_i[333]
  PIN w_data_i[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 58.835 161.495 58.905 ;
    END
  END w_data_i[334]
  PIN w_data_i[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 34.195 0.07 34.265 ;
    END
  END w_data_i[335]
  PIN w_data_i[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 49.875 161.495 49.945 ;
    END
  END w_data_i[336]
  PIN w_data_i[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  19.625 81.61 19.765 81.75 ;
    END
  END w_data_i[337]
  PIN w_data_i[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 25.515 161.495 25.585 ;
    END
  END w_data_i[338]
  PIN w_data_i[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 19.915 0.07 19.985 ;
    END
  END w_data_i[339]
  PIN w_data_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 45.395 161.495 45.465 ;
    END
  END w_data_i[33]
  PIN w_data_i[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  68.905 0 69.045 0.14 ;
    END
  END w_data_i[340]
  PIN w_data_i[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  160.745 81.61 160.885 81.75 ;
    END
  END w_data_i[341]
  PIN w_data_i[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 32.795 0.07 32.865 ;
    END
  END w_data_i[342]
  PIN w_data_i[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 33.075 0.07 33.145 ;
    END
  END w_data_i[343]
  PIN w_data_i[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  51.545 81.61 51.685 81.75 ;
    END
  END w_data_i[344]
  PIN w_data_i[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 2.275 161.495 2.345 ;
    END
  END w_data_i[345]
  PIN w_data_i[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  132.745 0 132.885 0.14 ;
    END
  END w_data_i[346]
  PIN w_data_i[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  16.265 0 16.405 0.14 ;
    END
  END w_data_i[347]
  PIN w_data_i[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  24.665 0 24.805 0.14 ;
    END
  END w_data_i[348]
  PIN w_data_i[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 18.235 161.495 18.305 ;
    END
  END w_data_i[349]
  PIN w_data_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 80.395 0.07 80.465 ;
    END
  END w_data_i[34]
  PIN w_data_i[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 79.275 0.07 79.345 ;
    END
  END w_data_i[350]
  PIN w_data_i[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 4.515 0.07 4.585 ;
    END
  END w_data_i[351]
  PIN w_data_i[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  128.265 0 128.405 0.14 ;
    END
  END w_data_i[352]
  PIN w_data_i[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.945 0 18.085 0.14 ;
    END
  END w_data_i[353]
  PIN w_data_i[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  2.825 81.61 2.965 81.75 ;
    END
  END w_data_i[354]
  PIN w_data_i[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 70.035 0.07 70.105 ;
    END
  END w_data_i[355]
  PIN w_data_i[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  71.705 0 71.845 0.14 ;
    END
  END w_data_i[356]
  PIN w_data_i[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  145.065 0 145.205 0.14 ;
    END
  END w_data_i[357]
  PIN w_data_i[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 77.595 0.07 77.665 ;
    END
  END w_data_i[358]
  PIN w_data_i[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 40.355 161.495 40.425 ;
    END
  END w_data_i[359]
  PIN w_data_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 57.435 0.07 57.505 ;
    END
  END w_data_i[35]
  PIN w_data_i[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  122.105 0 122.245 0.14 ;
    END
  END w_data_i[360]
  PIN w_data_i[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  119.865 0 120.005 0.14 ;
    END
  END w_data_i[361]
  PIN w_data_i[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  15.145 81.61 15.285 81.75 ;
    END
  END w_data_i[362]
  PIN w_data_i[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  123.785 0 123.925 0.14 ;
    END
  END w_data_i[363]
  PIN w_data_i[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  9.545 81.61 9.685 81.75 ;
    END
  END w_data_i[364]
  PIN w_data_i[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.945 0 32.085 0.14 ;
    END
  END w_data_i[365]
  PIN w_data_i[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 8.995 161.495 9.065 ;
    END
  END w_data_i[366]
  PIN w_data_i[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 18.795 161.495 18.865 ;
    END
  END w_data_i[367]
  PIN w_data_i[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 36.435 0.07 36.505 ;
    END
  END w_data_i[368]
  PIN w_data_i[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 18.515 0.07 18.585 ;
    END
  END w_data_i[369]
  PIN w_data_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 73.115 0.07 73.185 ;
    END
  END w_data_i[36]
  PIN w_data_i[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 56.595 0.07 56.665 ;
    END
  END w_data_i[370]
  PIN w_data_i[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  159.065 0 159.205 0.14 ;
    END
  END w_data_i[371]
  PIN w_data_i[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  82.905 0 83.045 0.14 ;
    END
  END w_data_i[372]
  PIN w_data_i[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  18.505 81.61 18.645 81.75 ;
    END
  END w_data_i[373]
  PIN w_data_i[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  120.425 0 120.565 0.14 ;
    END
  END w_data_i[374]
  PIN w_data_i[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 3.675 161.495 3.745 ;
    END
  END w_data_i[375]
  PIN w_data_i[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 8.155 0.07 8.225 ;
    END
  END w_data_i[376]
  PIN w_data_i[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 55.475 0.07 55.545 ;
    END
  END w_data_i[377]
  PIN w_data_i[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  139.465 81.61 139.605 81.75 ;
    END
  END w_data_i[378]
  PIN w_data_i[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  110.345 0 110.485 0.14 ;
    END
  END w_data_i[379]
  PIN w_data_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 0.875 0.07 0.945 ;
    END
  END w_data_i[37]
  PIN w_data_i[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 23.835 161.495 23.905 ;
    END
  END w_data_i[380]
  PIN w_data_i[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 52.955 161.495 53.025 ;
    END
  END w_data_i[381]
  PIN w_data_i[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 47.355 161.495 47.425 ;
    END
  END w_data_i[382]
  PIN w_data_i[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  82.345 0 82.485 0.14 ;
    END
  END w_data_i[383]
  PIN w_data_i[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  3.945 0 4.085 0.14 ;
    END
  END w_data_i[384]
  PIN w_data_i[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 64.435 0.07 64.505 ;
    END
  END w_data_i[385]
  PIN w_data_i[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  52.105 81.61 52.245 81.75 ;
    END
  END w_data_i[386]
  PIN w_data_i[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 8.435 161.495 8.505 ;
    END
  END w_data_i[387]
  PIN w_data_i[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 68.075 0.07 68.145 ;
    END
  END w_data_i[388]
  PIN w_data_i[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 8.435 0.07 8.505 ;
    END
  END w_data_i[389]
  PIN w_data_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 27.475 161.495 27.545 ;
    END
  END w_data_i[38]
  PIN w_data_i[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 11.795 0.07 11.865 ;
    END
  END w_data_i[390]
  PIN w_data_i[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 9.275 0.07 9.345 ;
    END
  END w_data_i[391]
  PIN w_data_i[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  137.225 0 137.365 0.14 ;
    END
  END w_data_i[392]
  PIN w_data_i[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 14.595 0.07 14.665 ;
    END
  END w_data_i[393]
  PIN w_data_i[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 30.835 0.07 30.905 ;
    END
  END w_data_i[394]
  PIN w_data_i[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  160.745 0 160.885 0.14 ;
    END
  END w_data_i[395]
  PIN w_data_i[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 13.195 0.07 13.265 ;
    END
  END w_data_i[396]
  PIN w_data_i[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.315 0.07 7.385 ;
    END
  END w_data_i[397]
  PIN w_data_i[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  62.185 0 62.325 0.14 ;
    END
  END w_data_i[398]
  PIN w_data_i[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 52.395 0.07 52.465 ;
    END
  END w_data_i[399]
  PIN w_data_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 40.915 0.07 40.985 ;
    END
  END w_data_i[39]
  PIN w_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 57.435 161.495 57.505 ;
    END
  END w_data_i[3]
  PIN w_data_i[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  32.505 81.61 32.645 81.75 ;
    END
  END w_data_i[400]
  PIN w_data_i[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 63.315 0.07 63.385 ;
    END
  END w_data_i[401]
  PIN w_data_i[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 26.635 161.495 26.705 ;
    END
  END w_data_i[402]
  PIN w_data_i[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  95.785 0 95.925 0.14 ;
    END
  END w_data_i[403]
  PIN w_data_i[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 40.635 0.07 40.705 ;
    END
  END w_data_i[404]
  PIN w_data_i[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  70.585 81.61 70.725 81.75 ;
    END
  END w_data_i[405]
  PIN w_data_i[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 37.275 161.495 37.345 ;
    END
  END w_data_i[406]
  PIN w_data_i[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 5.915 0.07 5.985 ;
    END
  END w_data_i[407]
  PIN w_data_i[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  54.345 0 54.485 0.14 ;
    END
  END w_data_i[408]
  PIN w_data_i[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  156.265 81.61 156.405 81.75 ;
    END
  END w_data_i[409]
  PIN w_data_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  152.345 0 152.485 0.14 ;
    END
  END w_data_i[40]
  PIN w_data_i[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  65.545 81.61 65.685 81.75 ;
    END
  END w_data_i[410]
  PIN w_data_i[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 49.315 0.07 49.385 ;
    END
  END w_data_i[411]
  PIN w_data_i[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  1.705 81.61 1.845 81.75 ;
    END
  END w_data_i[412]
  PIN w_data_i[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  26.905 81.61 27.045 81.75 ;
    END
  END w_data_i[413]
  PIN w_data_i[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  83.465 0 83.605 0.14 ;
    END
  END w_data_i[414]
  PIN w_data_i[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  122.105 81.61 122.245 81.75 ;
    END
  END w_data_i[415]
  PIN w_data_i[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  150.665 0 150.805 0.14 ;
    END
  END w_data_i[416]
  PIN w_data_i[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 75.915 161.495 75.985 ;
    END
  END w_data_i[417]
  PIN w_data_i[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  40.345 0 40.485 0.14 ;
    END
  END w_data_i[418]
  PIN w_data_i[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 76.475 0.07 76.545 ;
    END
  END w_data_i[419]
  PIN w_data_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  119.305 0 119.445 0.14 ;
    END
  END w_data_i[41]
  PIN w_data_i[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  106.425 0 106.565 0.14 ;
    END
  END w_data_i[420]
  PIN w_data_i[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  87.385 81.61 87.525 81.75 ;
    END
  END w_data_i[421]
  PIN w_data_i[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 61.355 161.495 61.425 ;
    END
  END w_data_i[422]
  PIN w_data_i[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 27.755 161.495 27.825 ;
    END
  END w_data_i[423]
  PIN w_data_i[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 78.715 161.495 78.785 ;
    END
  END w_data_i[424]
  PIN w_data_i[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  131.065 0 131.205 0.14 ;
    END
  END w_data_i[425]
  PIN w_data_i[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 23.275 0.07 23.345 ;
    END
  END w_data_i[426]
  PIN w_data_i[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 45.675 0.07 45.745 ;
    END
  END w_data_i[427]
  PIN w_data_i[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 48.195 0.07 48.265 ;
    END
  END w_data_i[428]
  PIN w_data_i[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 54.355 161.495 54.425 ;
    END
  END w_data_i[429]
  PIN w_data_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 68.915 161.495 68.985 ;
    END
  END w_data_i[42]
  PIN w_data_i[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 3.395 161.495 3.465 ;
    END
  END w_data_i[430]
  PIN w_data_i[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 45.955 161.495 46.025 ;
    END
  END w_data_i[431]
  PIN w_data_i[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  145.625 81.61 145.765 81.75 ;
    END
  END w_data_i[432]
  PIN w_data_i[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 35.595 0.07 35.665 ;
    END
  END w_data_i[433]
  PIN w_data_i[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  16.825 0 16.965 0.14 ;
    END
  END w_data_i[434]
  PIN w_data_i[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  107.545 0 107.685 0.14 ;
    END
  END w_data_i[435]
  PIN w_data_i[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  57.705 0 57.845 0.14 ;
    END
  END w_data_i[436]
  PIN w_data_i[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 36.995 161.495 37.065 ;
    END
  END w_data_i[437]
  PIN w_data_i[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.025 0 14.165 0.14 ;
    END
  END w_data_i[438]
  PIN w_data_i[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  59.385 0 59.525 0.14 ;
    END
  END w_data_i[439]
  PIN w_data_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 34.475 161.495 34.545 ;
    END
  END w_data_i[43]
  PIN w_data_i[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 15.155 0.07 15.225 ;
    END
  END w_data_i[440]
  PIN w_data_i[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 59.955 161.495 60.025 ;
    END
  END w_data_i[441]
  PIN w_data_i[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  21.865 0 22.005 0.14 ;
    END
  END w_data_i[442]
  PIN w_data_i[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 52.675 161.495 52.745 ;
    END
  END w_data_i[443]
  PIN w_data_i[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  137.785 0 137.925 0.14 ;
    END
  END w_data_i[444]
  PIN w_data_i[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 17.955 0.07 18.025 ;
    END
  END w_data_i[445]
  PIN w_data_i[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  127.145 0 127.285 0.14 ;
    END
  END w_data_i[446]
  PIN w_data_i[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 71.155 161.495 71.225 ;
    END
  END w_data_i[447]
  PIN w_data_i[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  93.545 81.61 93.685 81.75 ;
    END
  END w_data_i[448]
  PIN w_data_i[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  72.265 81.61 72.405 81.75 ;
    END
  END w_data_i[449]
  PIN w_data_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  24.105 81.61 24.245 81.75 ;
    END
  END w_data_i[44]
  PIN w_data_i[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  96.905 81.61 97.045 81.75 ;
    END
  END w_data_i[450]
  PIN w_data_i[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 59.115 0.07 59.185 ;
    END
  END w_data_i[451]
  PIN w_data_i[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  64.985 0 65.125 0.14 ;
    END
  END w_data_i[452]
  PIN w_data_i[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 24.115 161.495 24.185 ;
    END
  END w_data_i[453]
  PIN w_data_i[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 48.475 161.495 48.545 ;
    END
  END w_data_i[454]
  PIN w_data_i[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 72.555 161.495 72.625 ;
    END
  END w_data_i[455]
  PIN w_data_i[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 14.875 0.07 14.945 ;
    END
  END w_data_i[456]
  PIN w_data_i[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  149.545 0 149.685 0.14 ;
    END
  END w_data_i[457]
  PIN w_data_i[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  134.985 81.61 135.125 81.75 ;
    END
  END w_data_i[458]
  PIN w_data_i[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  159.625 81.61 159.765 81.75 ;
    END
  END w_data_i[459]
  PIN w_data_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  84.025 81.61 84.165 81.75 ;
    END
  END w_data_i[45]
  PIN w_data_i[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 23.555 0.07 23.625 ;
    END
  END w_data_i[460]
  PIN w_data_i[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 9.275 161.495 9.345 ;
    END
  END w_data_i[461]
  PIN w_data_i[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  115.945 81.61 116.085 81.75 ;
    END
  END w_data_i[462]
  PIN w_data_i[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 5.635 161.495 5.705 ;
    END
  END w_data_i[463]
  PIN w_data_i[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 36.155 0.07 36.225 ;
    END
  END w_data_i[464]
  PIN w_data_i[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  35.305 0 35.445 0.14 ;
    END
  END w_data_i[465]
  PIN w_data_i[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  52.665 0 52.805 0.14 ;
    END
  END w_data_i[466]
  PIN w_data_i[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 11.235 161.495 11.305 ;
    END
  END w_data_i[467]
  PIN w_data_i[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.355 0.07 12.425 ;
    END
  END w_data_i[468]
  PIN w_data_i[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  138.345 81.61 138.485 81.75 ;
    END
  END w_data_i[469]
  PIN w_data_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.905 81.61 13.045 81.75 ;
    END
  END w_data_i[46]
  PIN w_data_i[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  5.065 81.61 5.205 81.75 ;
    END
  END w_data_i[470]
  PIN w_data_i[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 68.635 0.07 68.705 ;
    END
  END w_data_i[471]
  PIN w_data_i[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  64.425 0 64.565 0.14 ;
    END
  END w_data_i[472]
  PIN w_data_i[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  121.545 81.61 121.685 81.75 ;
    END
  END w_data_i[473]
  PIN w_data_i[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 19.635 161.495 19.705 ;
    END
  END w_data_i[474]
  PIN w_data_i[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 64.715 0.07 64.785 ;
    END
  END w_data_i[475]
  PIN w_data_i[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  41.465 0 41.605 0.14 ;
    END
  END w_data_i[476]
  PIN w_data_i[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  145.065 81.61 145.205 81.75 ;
    END
  END w_data_i[477]
  PIN w_data_i[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 19.355 0.07 19.425 ;
    END
  END w_data_i[478]
  PIN w_data_i[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  41.465 81.61 41.605 81.75 ;
    END
  END w_data_i[479]
  PIN w_data_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  75.065 81.61 75.205 81.75 ;
    END
  END w_data_i[47]
  PIN w_data_i[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  84.585 81.61 84.725 81.75 ;
    END
  END w_data_i[480]
  PIN w_data_i[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  86.825 81.61 86.965 81.75 ;
    END
  END w_data_i[481]
  PIN w_data_i[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  111.465 0 111.605 0.14 ;
    END
  END w_data_i[482]
  PIN w_data_i[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  25.225 81.61 25.365 81.75 ;
    END
  END w_data_i[483]
  PIN w_data_i[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 19.075 0.07 19.145 ;
    END
  END w_data_i[484]
  PIN w_data_i[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  3.385 0 3.525 0.14 ;
    END
  END w_data_i[485]
  PIN w_data_i[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 2.835 161.495 2.905 ;
    END
  END w_data_i[486]
  PIN w_data_i[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  112.025 0 112.165 0.14 ;
    END
  END w_data_i[487]
  PIN w_data_i[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 31.395 161.495 31.465 ;
    END
  END w_data_i[488]
  PIN w_data_i[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  47.065 81.61 47.205 81.75 ;
    END
  END w_data_i[489]
  PIN w_data_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 39.795 161.495 39.865 ;
    END
  END w_data_i[48]
  PIN w_data_i[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 43.155 0.07 43.225 ;
    END
  END w_data_i[490]
  PIN w_data_i[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  8.985 0 9.125 0.14 ;
    END
  END w_data_i[491]
  PIN w_data_i[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  42.585 0 42.725 0.14 ;
    END
  END w_data_i[492]
  PIN w_data_i[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  94.105 0 94.245 0.14 ;
    END
  END w_data_i[493]
  PIN w_data_i[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  27.465 81.61 27.605 81.75 ;
    END
  END w_data_i[494]
  PIN w_data_i[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 4.515 161.495 4.585 ;
    END
  END w_data_i[495]
  PIN w_data_i[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  80.105 0 80.245 0.14 ;
    END
  END w_data_i[496]
  PIN w_data_i[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  157.385 0 157.525 0.14 ;
    END
  END w_data_i[497]
  PIN w_data_i[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 74.795 161.495 74.865 ;
    END
  END w_data_i[498]
  PIN w_data_i[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  136.105 81.61 136.245 81.75 ;
    END
  END w_data_i[499]
  PIN w_data_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  160.185 0 160.325 0.14 ;
    END
  END w_data_i[49]
  PIN w_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 46.235 0.07 46.305 ;
    END
  END w_data_i[4]
  PIN w_data_i[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 22.155 161.495 22.225 ;
    END
  END w_data_i[500]
  PIN w_data_i[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  146.185 81.61 146.325 81.75 ;
    END
  END w_data_i[501]
  PIN w_data_i[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.865 81.61 8.005 81.75 ;
    END
  END w_data_i[502]
  PIN w_data_i[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 75.075 161.495 75.145 ;
    END
  END w_data_i[503]
  PIN w_data_i[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  155.705 0 155.845 0.14 ;
    END
  END w_data_i[504]
  PIN w_data_i[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  52.665 81.61 52.805 81.75 ;
    END
  END w_data_i[505]
  PIN w_data_i[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 31.955 161.495 32.025 ;
    END
  END w_data_i[506]
  PIN w_data_i[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 78.715 0.07 78.785 ;
    END
  END w_data_i[507]
  PIN w_data_i[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 14.035 161.495 14.105 ;
    END
  END w_data_i[508]
  PIN w_data_i[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 44.555 0.07 44.625 ;
    END
  END w_data_i[509]
  PIN w_data_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  26.345 0 26.485 0.14 ;
    END
  END w_data_i[50]
  PIN w_data_i[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 70.595 161.495 70.665 ;
    END
  END w_data_i[510]
  PIN w_data_i[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  113.705 0 113.845 0.14 ;
    END
  END w_data_i[511]
  PIN w_data_i[512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  151.785 81.61 151.925 81.75 ;
    END
  END w_data_i[512]
  PIN w_data_i[513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  51.545 0 51.685 0.14 ;
    END
  END w_data_i[513]
  PIN w_data_i[514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 14.875 161.495 14.945 ;
    END
  END w_data_i[514]
  PIN w_data_i[515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 54.075 0.07 54.145 ;
    END
  END w_data_i[515]
  PIN w_data_i[516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  59.385 81.61 59.525 81.75 ;
    END
  END w_data_i[516]
  PIN w_data_i[517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  134.425 81.61 134.565 81.75 ;
    END
  END w_data_i[517]
  PIN w_data_i[518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 52.115 0.07 52.185 ;
    END
  END w_data_i[518]
  PIN w_data_i[519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 61.075 0.07 61.145 ;
    END
  END w_data_i[519]
  PIN w_data_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 35.595 161.495 35.665 ;
    END
  END w_data_i[51]
  PIN w_data_i[520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 47.635 0.07 47.705 ;
    END
  END w_data_i[520]
  PIN w_data_i[521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 51.835 161.495 51.905 ;
    END
  END w_data_i[521]
  PIN w_data_i[522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  28.585 81.61 28.725 81.75 ;
    END
  END w_data_i[522]
  PIN w_data_i[523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 75.075 0.07 75.145 ;
    END
  END w_data_i[523]
  PIN w_data_i[524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 37.555 0.07 37.625 ;
    END
  END w_data_i[524]
  PIN w_data_i[525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  18.505 0 18.645 0.14 ;
    END
  END w_data_i[525]
  PIN w_data_i[526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  108.665 0 108.805 0.14 ;
    END
  END w_data_i[526]
  PIN w_data_i[527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  148.425 81.61 148.565 81.75 ;
    END
  END w_data_i[527]
  PIN w_data_i[528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  160.185 81.61 160.325 81.75 ;
    END
  END w_data_i[528]
  PIN w_data_i[529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 15.435 0.07 15.505 ;
    END
  END w_data_i[529]
  PIN w_data_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 73.675 161.495 73.745 ;
    END
  END w_data_i[52]
  PIN w_data_i[530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 45.675 161.495 45.745 ;
    END
  END w_data_i[530]
  PIN w_data_i[531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 12.355 161.495 12.425 ;
    END
  END w_data_i[531]
  PIN w_data_i[532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  35.865 81.61 36.005 81.75 ;
    END
  END w_data_i[532]
  PIN w_data_i[533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  90.185 81.61 90.325 81.75 ;
    END
  END w_data_i[533]
  PIN w_data_i[534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  108.105 0 108.245 0.14 ;
    END
  END w_data_i[534]
  PIN w_data_i[535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  153.465 0 153.605 0.14 ;
    END
  END w_data_i[535]
  PIN w_data_i[536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 20.755 0.07 20.825 ;
    END
  END w_data_i[536]
  PIN w_data_i[537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 51.835 0.07 51.905 ;
    END
  END w_data_i[537]
  PIN w_data_i[538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  103.065 0 103.205 0.14 ;
    END
  END w_data_i[538]
  PIN w_data_i[539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  20.745 0 20.885 0.14 ;
    END
  END w_data_i[539]
  PIN w_data_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 73.675 0.07 73.745 ;
    END
  END w_data_i[53]
  PIN w_data_i[540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 67.795 161.495 67.865 ;
    END
  END w_data_i[540]
  PIN w_data_i[541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  118.185 81.61 118.325 81.75 ;
    END
  END w_data_i[541]
  PIN w_data_i[542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  73.385 0 73.525 0.14 ;
    END
  END w_data_i[542]
  PIN w_data_i[543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  73.385 81.61 73.525 81.75 ;
    END
  END w_data_i[543]
  PIN w_data_i[544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 52.115 161.495 52.185 ;
    END
  END w_data_i[544]
  PIN w_data_i[545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  144.505 0 144.645 0.14 ;
    END
  END w_data_i[545]
  PIN w_data_i[546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  71.705 81.61 71.845 81.75 ;
    END
  END w_data_i[546]
  PIN w_data_i[547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  138.905 0 139.045 0.14 ;
    END
  END w_data_i[547]
  PIN w_data_i[548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  58.825 0 58.965 0.14 ;
    END
  END w_data_i[548]
  PIN w_data_i[549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.105 0 10.245 0.14 ;
    END
  END w_data_i[549]
  PIN w_data_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 12.075 161.495 12.145 ;
    END
  END w_data_i[54]
  PIN w_data_i[550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 36.435 161.495 36.505 ;
    END
  END w_data_i[550]
  PIN w_data_i[551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 78.155 0.07 78.225 ;
    END
  END w_data_i[551]
  PIN w_data_i[552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  142.265 81.61 142.405 81.75 ;
    END
  END w_data_i[552]
  PIN w_data_i[553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 30.275 0.07 30.345 ;
    END
  END w_data_i[553]
  PIN w_data_i[554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 36.995 0.07 37.065 ;
    END
  END w_data_i[554]
  PIN w_data_i[555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 34.755 0.07 34.825 ;
    END
  END w_data_i[555]
  PIN w_data_i[556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  8.425 0 8.565 0.14 ;
    END
  END w_data_i[556]
  PIN w_data_i[557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  39.785 0 39.925 0.14 ;
    END
  END w_data_i[557]
  PIN w_data_i[558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 56.875 161.495 56.945 ;
    END
  END w_data_i[558]
  PIN w_data_i[559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  103.625 0 103.765 0.14 ;
    END
  END w_data_i[559]
  PIN w_data_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  68.345 81.61 68.485 81.75 ;
    END
  END w_data_i[55]
  PIN w_data_i[560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  112.585 81.61 112.725 81.75 ;
    END
  END w_data_i[560]
  PIN w_data_i[561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.595 0.07 7.665 ;
    END
  END w_data_i[561]
  PIN w_data_i[562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  28.585 0 28.725 0.14 ;
    END
  END w_data_i[562]
  PIN w_data_i[563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 62.755 161.495 62.825 ;
    END
  END w_data_i[563]
  PIN w_data_i[564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  120.425 81.61 120.565 81.75 ;
    END
  END w_data_i[564]
  PIN w_data_i[565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 13.475 0.07 13.545 ;
    END
  END w_data_i[565]
  PIN w_data_i[566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 77.595 161.495 77.665 ;
    END
  END w_data_i[566]
  PIN w_data_i[567]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 37.555 161.495 37.625 ;
    END
  END w_data_i[567]
  PIN w_data_i[568]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  122.665 0 122.805 0.14 ;
    END
  END w_data_i[568]
  PIN w_data_i[569]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  102.505 81.61 102.645 81.75 ;
    END
  END w_data_i[569]
  PIN w_data_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 80.675 0.07 80.745 ;
    END
  END w_data_i[56]
  PIN w_data_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  56.025 0 56.165 0.14 ;
    END
  END w_data_i[57]
  PIN w_data_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 60.515 161.495 60.585 ;
    END
  END w_data_i[58]
  PIN w_data_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  143.385 0 143.525 0.14 ;
    END
  END w_data_i[59]
  PIN w_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 33.075 161.495 33.145 ;
    END
  END w_data_i[5]
  PIN w_data_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.315 0.07 21.385 ;
    END
  END w_data_i[60]
  PIN w_data_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 10.395 161.495 10.465 ;
    END
  END w_data_i[61]
  PIN w_data_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  29.145 0 29.285 0.14 ;
    END
  END w_data_i[62]
  PIN w_data_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  86.825 0 86.965 0.14 ;
    END
  END w_data_i[63]
  PIN w_data_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 43.995 161.495 44.065 ;
    END
  END w_data_i[64]
  PIN w_data_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  103.065 81.61 103.205 81.75 ;
    END
  END w_data_i[65]
  PIN w_data_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  156.825 81.61 156.965 81.75 ;
    END
  END w_data_i[66]
  PIN w_data_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 10.675 161.495 10.745 ;
    END
  END w_data_i[67]
  PIN w_data_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.585 0 14.725 0.14 ;
    END
  END w_data_i[68]
  PIN w_data_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 54.635 161.495 54.705 ;
    END
  END w_data_i[69]
  PIN w_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  4.505 0 4.645 0.14 ;
    END
  END w_data_i[6]
  PIN w_data_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  155.145 81.61 155.285 81.75 ;
    END
  END w_data_i[70]
  PIN w_data_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  100.825 81.61 100.965 81.75 ;
    END
  END w_data_i[71]
  PIN w_data_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 15.155 161.495 15.225 ;
    END
  END w_data_i[72]
  PIN w_data_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  96.345 81.61 96.485 81.75 ;
    END
  END w_data_i[73]
  PIN w_data_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  114.825 0 114.965 0.14 ;
    END
  END w_data_i[74]
  PIN w_data_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 11.235 0.07 11.305 ;
    END
  END w_data_i[75]
  PIN w_data_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  114.265 0 114.405 0.14 ;
    END
  END w_data_i[76]
  PIN w_data_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END w_data_i[77]
  PIN w_data_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  133.305 0 133.445 0.14 ;
    END
  END w_data_i[78]
  PIN w_data_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 26.915 0.07 26.985 ;
    END
  END w_data_i[79]
  PIN w_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 59.955 0.07 60.025 ;
    END
  END w_data_i[7]
  PIN w_data_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  28.025 81.61 28.165 81.75 ;
    END
  END w_data_i[80]
  PIN w_data_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 16.275 0.07 16.345 ;
    END
  END w_data_i[81]
  PIN w_data_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  35.865 0 36.005 0.14 ;
    END
  END w_data_i[82]
  PIN w_data_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  13.465 0 13.605 0.14 ;
    END
  END w_data_i[83]
  PIN w_data_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  71.145 81.61 71.285 81.75 ;
    END
  END w_data_i[84]
  PIN w_data_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.745 81.61 34.885 81.75 ;
    END
  END w_data_i[85]
  PIN w_data_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  90.745 0 90.885 0.14 ;
    END
  END w_data_i[86]
  PIN w_data_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 2.835 0.07 2.905 ;
    END
  END w_data_i[87]
  PIN w_data_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 26.075 161.495 26.145 ;
    END
  END w_data_i[88]
  PIN w_data_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 47.075 0.07 47.145 ;
    END
  END w_data_i[89]
  PIN w_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 66.115 161.495 66.185 ;
    END
  END w_data_i[8]
  PIN w_data_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  36.985 0 37.125 0.14 ;
    END
  END w_data_i[90]
  PIN w_data_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  63.865 0 64.005 0.14 ;
    END
  END w_data_i[91]
  PIN w_data_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 3.115 0.07 3.185 ;
    END
  END w_data_i[92]
  PIN w_data_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 62.195 161.495 62.265 ;
    END
  END w_data_i[93]
  PIN w_data_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  99.705 0 99.845 0.14 ;
    END
  END w_data_i[94]
  PIN w_data_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  101.385 81.61 101.525 81.75 ;
    END
  END w_data_i[95]
  PIN w_data_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  99.705 81.61 99.845 81.75 ;
    END
  END w_data_i[96]
  PIN w_data_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 72.555 0.07 72.625 ;
    END
  END w_data_i[97]
  PIN w_data_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.025 81.61 14.165 81.75 ;
    END
  END w_data_i[98]
  PIN w_data_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  117.625 0 117.765 0.14 ;
    END
  END w_data_i[99]
  PIN w_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 17.115 0.07 17.185 ;
    END
  END w_data_i[9]
  PIN w_reset_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 66.115 0.07 66.185 ;
    END
  END w_reset_i
  PIN w_v_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  161.425 40.635 161.495 40.705 ;
    END
  END w_v_i
  OBS
    LAYER metal1 ;
     RECT  0 -0.085 3.23 81.75 ;
     RECT  3.23 0 161.495 81.75 ;
    LAYER metal2 ;
     RECT  0 0 161.495 81.75 ;
    LAYER metal3 ;
     RECT  0 0 161.495 81.75 ;
    LAYER metal4 ;
     RECT  0 0 161.495 81.75 ;
  END
END bsg_mem_p570
END LIBRARY
