VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MACRO bsg_mem_p540
  FOREIGN bsg_mem_p540 0 0 ;
  CLASS BLOCK ;
  SIZE 146.865 BY 190.32 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 188.915 145.73 189.085 ;
        RECT  1.14 186.115 145.73 186.285 ;
        RECT  1.14 183.315 145.73 183.485 ;
        RECT  1.14 180.515 145.73 180.685 ;
        RECT  1.14 177.715 145.73 177.885 ;
        RECT  1.14 174.915 145.73 175.085 ;
        RECT  1.14 172.115 145.73 172.285 ;
        RECT  1.14 169.315 145.73 169.485 ;
        RECT  1.14 166.515 145.73 166.685 ;
        RECT  1.14 163.715 145.73 163.885 ;
        RECT  1.14 160.915 145.73 161.085 ;
        RECT  1.14 158.115 145.73 158.285 ;
        RECT  1.14 155.315 145.73 155.485 ;
        RECT  1.14 152.515 145.73 152.685 ;
        RECT  1.14 149.715 145.73 149.885 ;
        RECT  1.14 146.915 145.73 147.085 ;
        RECT  1.14 144.115 145.73 144.285 ;
        RECT  1.14 141.315 145.73 141.485 ;
        RECT  1.14 138.515 145.73 138.685 ;
        RECT  1.14 135.715 145.73 135.885 ;
        RECT  1.14 132.915 145.73 133.085 ;
        RECT  1.14 130.115 145.73 130.285 ;
        RECT  1.14 127.315 145.73 127.485 ;
        RECT  1.14 124.515 145.73 124.685 ;
        RECT  1.14 121.715 145.73 121.885 ;
        RECT  1.14 118.915 145.73 119.085 ;
        RECT  1.14 116.115 145.73 116.285 ;
        RECT  1.14 113.315 145.73 113.485 ;
        RECT  1.14 110.515 145.73 110.685 ;
        RECT  1.14 107.715 145.73 107.885 ;
        RECT  1.14 104.915 145.73 105.085 ;
        RECT  1.14 102.115 145.73 102.285 ;
        RECT  1.14 99.315 145.73 99.485 ;
        RECT  1.14 96.515 145.73 96.685 ;
        RECT  1.14 93.715 145.73 93.885 ;
        RECT  1.14 90.915 145.73 91.085 ;
        RECT  1.14 88.115 145.73 88.285 ;
        RECT  1.14 85.315 145.73 85.485 ;
        RECT  1.14 82.515 145.73 82.685 ;
        RECT  1.14 79.715 145.73 79.885 ;
        RECT  1.14 76.915 145.73 77.085 ;
        RECT  1.14 74.115 145.73 74.285 ;
        RECT  1.14 71.315 145.73 71.485 ;
        RECT  1.14 68.515 145.73 68.685 ;
        RECT  1.14 65.715 145.73 65.885 ;
        RECT  1.14 62.915 145.73 63.085 ;
        RECT  1.14 60.115 145.73 60.285 ;
        RECT  1.14 57.315 145.73 57.485 ;
        RECT  1.14 54.515 145.73 54.685 ;
        RECT  1.14 51.715 145.73 51.885 ;
        RECT  1.14 48.915 145.73 49.085 ;
        RECT  1.14 46.115 145.73 46.285 ;
        RECT  1.14 43.315 145.73 43.485 ;
        RECT  1.14 40.515 145.73 40.685 ;
        RECT  1.14 37.715 145.73 37.885 ;
        RECT  1.14 34.915 145.73 35.085 ;
        RECT  1.14 32.115 145.73 32.285 ;
        RECT  1.14 29.315 145.73 29.485 ;
        RECT  1.14 26.515 145.73 26.685 ;
        RECT  1.14 23.715 145.73 23.885 ;
        RECT  1.14 20.915 145.73 21.085 ;
        RECT  1.14 18.115 145.73 18.285 ;
        RECT  1.14 15.315 145.73 15.485 ;
        RECT  1.14 12.515 145.73 12.685 ;
        RECT  1.14 9.715 145.73 9.885 ;
        RECT  1.14 6.915 145.73 7.085 ;
        RECT  1.14 4.115 145.73 4.285 ;
        RECT  1.14 1.315 145.73 1.485 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 187.515 145.73 187.685 ;
        RECT  1.14 184.715 145.73 184.885 ;
        RECT  1.14 181.915 145.73 182.085 ;
        RECT  1.14 179.115 145.73 179.285 ;
        RECT  1.14 176.315 145.73 176.485 ;
        RECT  1.14 173.515 145.73 173.685 ;
        RECT  1.14 170.715 145.73 170.885 ;
        RECT  1.14 167.915 145.73 168.085 ;
        RECT  1.14 165.115 145.73 165.285 ;
        RECT  1.14 162.315 145.73 162.485 ;
        RECT  1.14 159.515 145.73 159.685 ;
        RECT  1.14 156.715 145.73 156.885 ;
        RECT  1.14 153.915 145.73 154.085 ;
        RECT  1.14 151.115 145.73 151.285 ;
        RECT  1.14 148.315 145.73 148.485 ;
        RECT  1.14 145.515 145.73 145.685 ;
        RECT  1.14 142.715 145.73 142.885 ;
        RECT  1.14 139.915 145.73 140.085 ;
        RECT  1.14 137.115 145.73 137.285 ;
        RECT  1.14 134.315 145.73 134.485 ;
        RECT  1.14 131.515 145.73 131.685 ;
        RECT  1.14 128.715 145.73 128.885 ;
        RECT  1.14 125.915 145.73 126.085 ;
        RECT  1.14 123.115 145.73 123.285 ;
        RECT  1.14 120.315 145.73 120.485 ;
        RECT  1.14 117.515 145.73 117.685 ;
        RECT  1.14 114.715 145.73 114.885 ;
        RECT  1.14 111.915 145.73 112.085 ;
        RECT  1.14 109.115 145.73 109.285 ;
        RECT  1.14 106.315 145.73 106.485 ;
        RECT  1.14 103.515 145.73 103.685 ;
        RECT  1.14 100.715 145.73 100.885 ;
        RECT  1.14 97.915 145.73 98.085 ;
        RECT  1.14 95.115 145.73 95.285 ;
        RECT  1.14 92.315 145.73 92.485 ;
        RECT  1.14 89.515 145.73 89.685 ;
        RECT  1.14 86.715 145.73 86.885 ;
        RECT  1.14 83.915 145.73 84.085 ;
        RECT  1.14 81.115 145.73 81.285 ;
        RECT  1.14 78.315 145.73 78.485 ;
        RECT  1.14 75.515 145.73 75.685 ;
        RECT  1.14 72.715 145.73 72.885 ;
        RECT  1.14 69.915 145.73 70.085 ;
        RECT  1.14 67.115 145.73 67.285 ;
        RECT  1.14 64.315 145.73 64.485 ;
        RECT  1.14 61.515 145.73 61.685 ;
        RECT  1.14 58.715 145.73 58.885 ;
        RECT  1.14 55.915 145.73 56.085 ;
        RECT  1.14 53.115 145.73 53.285 ;
        RECT  1.14 50.315 145.73 50.485 ;
        RECT  1.14 47.515 145.73 47.685 ;
        RECT  1.14 44.715 145.73 44.885 ;
        RECT  1.14 41.915 145.73 42.085 ;
        RECT  1.14 39.115 145.73 39.285 ;
        RECT  1.14 36.315 145.73 36.485 ;
        RECT  1.14 33.515 145.73 33.685 ;
        RECT  1.14 30.715 145.73 30.885 ;
        RECT  1.14 27.915 145.73 28.085 ;
        RECT  1.14 25.115 145.73 25.285 ;
        RECT  1.14 22.315 145.73 22.485 ;
        RECT  1.14 19.515 145.73 19.685 ;
        RECT  1.14 16.715 145.73 16.885 ;
        RECT  1.14 13.915 145.73 14.085 ;
        RECT  1.14 11.115 145.73 11.285 ;
        RECT  1.14 8.315 145.73 8.485 ;
        RECT  1.14 5.515 145.73 5.685 ;
        RECT  1.14 2.715 145.73 2.885 ;
    END
  END VDD
  PIN r_addr_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  54.345 0 54.485 0.14 ;
    END
  END r_addr_i
  PIN r_data_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  24.665 190.18 24.805 190.32 ;
    END
  END r_data_o[0]
  PIN r_data_o[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 28.035 146.865 28.105 ;
    END
  END r_data_o[100]
  PIN r_data_o[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.105 0 10.245 0.14 ;
    END
  END r_data_o[101]
  PIN r_data_o[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 39.235 0.07 39.305 ;
    END
  END r_data_o[102]
  PIN r_data_o[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 3.115 146.865 3.185 ;
    END
  END r_data_o[103]
  PIN r_data_o[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 145.075 146.865 145.145 ;
    END
  END r_data_o[104]
  PIN r_data_o[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 117.635 0.07 117.705 ;
    END
  END r_data_o[105]
  PIN r_data_o[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 136.955 146.865 137.025 ;
    END
  END r_data_o[106]
  PIN r_data_o[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.185 0 34.325 0.14 ;
    END
  END r_data_o[107]
  PIN r_data_o[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 182.875 0.07 182.945 ;
    END
  END r_data_o[108]
  PIN r_data_o[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 115.395 146.865 115.465 ;
    END
  END r_data_o[109]
  PIN r_data_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 49.315 0.07 49.385 ;
    END
  END r_data_o[10]
  PIN r_data_o[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  86.265 0 86.405 0.14 ;
    END
  END r_data_o[110]
  PIN r_data_o[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 168.875 0.07 168.945 ;
    END
  END r_data_o[111]
  PIN r_data_o[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 180.915 146.865 180.985 ;
    END
  END r_data_o[112]
  PIN r_data_o[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  114.825 0 114.965 0.14 ;
    END
  END r_data_o[113]
  PIN r_data_o[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  80.105 0 80.245 0.14 ;
    END
  END r_data_o[114]
  PIN r_data_o[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 112.315 146.865 112.385 ;
    END
  END r_data_o[115]
  PIN r_data_o[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.355 0.07 12.425 ;
    END
  END r_data_o[116]
  PIN r_data_o[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  70.585 190.18 70.725 190.32 ;
    END
  END r_data_o[117]
  PIN r_data_o[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 72.555 0.07 72.625 ;
    END
  END r_data_o[118]
  PIN r_data_o[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 155.715 0.07 155.785 ;
    END
  END r_data_o[119]
  PIN r_data_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 131.635 146.865 131.705 ;
    END
  END r_data_o[11]
  PIN r_data_o[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 102.795 146.865 102.865 ;
    END
  END r_data_o[120]
  PIN r_data_o[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 56.035 146.865 56.105 ;
    END
  END r_data_o[121]
  PIN r_data_o[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  95.785 0 95.925 0.14 ;
    END
  END r_data_o[122]
  PIN r_data_o[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  43.705 190.18 43.845 190.32 ;
    END
  END r_data_o[123]
  PIN r_data_o[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 52.395 0.07 52.465 ;
    END
  END r_data_o[124]
  PIN r_data_o[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  67.785 190.18 67.925 190.32 ;
    END
  END r_data_o[125]
  PIN r_data_o[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 122.115 0.07 122.185 ;
    END
  END r_data_o[126]
  PIN r_data_o[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.865 0 8.005 0.14 ;
    END
  END r_data_o[127]
  PIN r_data_o[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  3.945 0 4.085 0.14 ;
    END
  END r_data_o[128]
  PIN r_data_o[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  66.105 190.18 66.245 190.32 ;
    END
  END r_data_o[129]
  PIN r_data_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 110.915 0.07 110.985 ;
    END
  END r_data_o[12]
  PIN r_data_o[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 35.035 0.07 35.105 ;
    END
  END r_data_o[130]
  PIN r_data_o[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  125.465 190.18 125.605 190.32 ;
    END
  END r_data_o[131]
  PIN r_data_o[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.105 190.18 10.245 190.32 ;
    END
  END r_data_o[132]
  PIN r_data_o[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  56.585 190.18 56.725 190.32 ;
    END
  END r_data_o[133]
  PIN r_data_o[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  77.305 190.18 77.445 190.32 ;
    END
  END r_data_o[134]
  PIN r_data_o[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 150.395 146.865 150.465 ;
    END
  END r_data_o[135]
  PIN r_data_o[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 59.955 0.07 60.025 ;
    END
  END r_data_o[136]
  PIN r_data_o[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 1.715 146.865 1.785 ;
    END
  END r_data_o[137]
  PIN r_data_o[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 27.755 146.865 27.825 ;
    END
  END r_data_o[138]
  PIN r_data_o[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 90.195 0.07 90.265 ;
    END
  END r_data_o[139]
  PIN r_data_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 64.715 0.07 64.785 ;
    END
  END r_data_o[13]
  PIN r_data_o[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 173.635 0.07 173.705 ;
    END
  END r_data_o[140]
  PIN r_data_o[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 126.315 0.07 126.385 ;
    END
  END r_data_o[141]
  PIN r_data_o[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  101.385 0 101.525 0.14 ;
    END
  END r_data_o[142]
  PIN r_data_o[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  54.345 190.18 54.485 190.32 ;
    END
  END r_data_o[143]
  PIN r_data_o[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 31.955 146.865 32.025 ;
    END
  END r_data_o[144]
  PIN r_data_o[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.905 190.18 13.045 190.32 ;
    END
  END r_data_o[145]
  PIN r_data_o[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 141.715 146.865 141.785 ;
    END
  END r_data_o[146]
  PIN r_data_o[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 75.355 146.865 75.425 ;
    END
  END r_data_o[147]
  PIN r_data_o[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 87.955 146.865 88.025 ;
    END
  END r_data_o[148]
  PIN r_data_o[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.315 0.07 21.385 ;
    END
  END r_data_o[149]
  PIN r_data_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 136.395 146.865 136.465 ;
    END
  END r_data_o[14]
  PIN r_data_o[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 181.475 0.07 181.545 ;
    END
  END r_data_o[150]
  PIN r_data_o[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 167.475 0.07 167.545 ;
    END
  END r_data_o[151]
  PIN r_data_o[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  49.305 0 49.445 0.14 ;
    END
  END r_data_o[152]
  PIN r_data_o[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 43.995 0.07 44.065 ;
    END
  END r_data_o[153]
  PIN r_data_o[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 172.795 0.07 172.865 ;
    END
  END r_data_o[154]
  PIN r_data_o[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 128.835 0.07 128.905 ;
    END
  END r_data_o[155]
  PIN r_data_o[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 86.275 146.865 86.345 ;
    END
  END r_data_o[156]
  PIN r_data_o[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  25.225 190.18 25.365 190.32 ;
    END
  END r_data_o[157]
  PIN r_data_o[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  101.385 190.18 101.525 190.32 ;
    END
  END r_data_o[158]
  PIN r_data_o[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 73.395 146.865 73.465 ;
    END
  END r_data_o[159]
  PIN r_data_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  47.625 0 47.765 0.14 ;
    END
  END r_data_o[15]
  PIN r_data_o[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.385 190.18 31.525 190.32 ;
    END
  END r_data_o[160]
  PIN r_data_o[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  105.305 190.18 105.445 190.32 ;
    END
  END r_data_o[161]
  PIN r_data_o[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 43.715 0.07 43.785 ;
    END
  END r_data_o[162]
  PIN r_data_o[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 53.235 0.07 53.305 ;
    END
  END r_data_o[163]
  PIN r_data_o[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 160.755 0.07 160.825 ;
    END
  END r_data_o[164]
  PIN r_data_o[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  47.625 190.18 47.765 190.32 ;
    END
  END r_data_o[165]
  PIN r_data_o[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 7.875 146.865 7.945 ;
    END
  END r_data_o[166]
  PIN r_data_o[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 66.115 0.07 66.185 ;
    END
  END r_data_o[167]
  PIN r_data_o[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 52.675 0.07 52.745 ;
    END
  END r_data_o[168]
  PIN r_data_o[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  51.545 0 51.685 0.14 ;
    END
  END r_data_o[169]
  PIN r_data_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 180.355 146.865 180.425 ;
    END
  END r_data_o[16]
  PIN r_data_o[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 103.355 146.865 103.425 ;
    END
  END r_data_o[170]
  PIN r_data_o[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 185.675 0.07 185.745 ;
    END
  END r_data_o[171]
  PIN r_data_o[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 161.595 146.865 161.665 ;
    END
  END r_data_o[172]
  PIN r_data_o[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 173.915 146.865 173.985 ;
    END
  END r_data_o[173]
  PIN r_data_o[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 134.995 146.865 135.065 ;
    END
  END r_data_o[174]
  PIN r_data_o[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 78.715 0.07 78.785 ;
    END
  END r_data_o[175]
  PIN r_data_o[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  51.545 190.18 51.685 190.32 ;
    END
  END r_data_o[176]
  PIN r_data_o[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 75.915 0.07 75.985 ;
    END
  END r_data_o[177]
  PIN r_data_o[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 139.475 146.865 139.545 ;
    END
  END r_data_o[178]
  PIN r_data_o[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  97.465 190.18 97.605 190.32 ;
    END
  END r_data_o[179]
  PIN r_data_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 80.675 0.07 80.745 ;
    END
  END r_data_o[17]
  PIN r_data_o[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 182.595 146.865 182.665 ;
    END
  END r_data_o[180]
  PIN r_data_o[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 87.395 146.865 87.465 ;
    END
  END r_data_o[181]
  PIN r_data_o[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 118.755 0.07 118.825 ;
    END
  END r_data_o[182]
  PIN r_data_o[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  52.105 0 52.245 0.14 ;
    END
  END r_data_o[183]
  PIN r_data_o[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 153.475 0.07 153.545 ;
    END
  END r_data_o[184]
  PIN r_data_o[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  85.145 190.18 85.285 190.32 ;
    END
  END r_data_o[185]
  PIN r_data_o[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 119.035 146.865 119.105 ;
    END
  END r_data_o[186]
  PIN r_data_o[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 45.115 0.07 45.185 ;
    END
  END r_data_o[187]
  PIN r_data_o[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 151.515 0.07 151.585 ;
    END
  END r_data_o[188]
  PIN r_data_o[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 66.115 146.865 66.185 ;
    END
  END r_data_o[189]
  PIN r_data_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 62.195 146.865 62.265 ;
    END
  END r_data_o[18]
  PIN r_data_o[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  27.465 0 27.605 0.14 ;
    END
  END r_data_o[190]
  PIN r_data_o[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 156.835 146.865 156.905 ;
    END
  END r_data_o[191]
  PIN r_data_o[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  62.185 0 62.325 0.14 ;
    END
  END r_data_o[192]
  PIN r_data_o[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 149.835 146.865 149.905 ;
    END
  END r_data_o[193]
  PIN r_data_o[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 98.875 0.07 98.945 ;
    END
  END r_data_o[194]
  PIN r_data_o[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  40.905 0 41.045 0.14 ;
    END
  END r_data_o[195]
  PIN r_data_o[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  92.985 0 93.125 0.14 ;
    END
  END r_data_o[196]
  PIN r_data_o[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 131.355 0.07 131.425 ;
    END
  END r_data_o[197]
  PIN r_data_o[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 104.195 0.07 104.265 ;
    END
  END r_data_o[198]
  PIN r_data_o[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  133.305 190.18 133.445 190.32 ;
    END
  END r_data_o[199]
  PIN r_data_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  30.265 0 30.405 0.14 ;
    END
  END r_data_o[19]
  PIN r_data_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 46.515 146.865 46.585 ;
    END
  END r_data_o[1]
  PIN r_data_o[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 114.835 146.865 114.905 ;
    END
  END r_data_o[200]
  PIN r_data_o[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  23.545 190.18 23.685 190.32 ;
    END
  END r_data_o[201]
  PIN r_data_o[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  100.265 0 100.405 0.14 ;
    END
  END r_data_o[202]
  PIN r_data_o[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 53.795 0.07 53.865 ;
    END
  END r_data_o[203]
  PIN r_data_o[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 65.555 146.865 65.625 ;
    END
  END r_data_o[204]
  PIN r_data_o[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 148.715 0.07 148.785 ;
    END
  END r_data_o[205]
  PIN r_data_o[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 84.035 0.07 84.105 ;
    END
  END r_data_o[206]
  PIN r_data_o[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  145.065 190.18 145.205 190.32 ;
    END
  END r_data_o[207]
  PIN r_data_o[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 77.595 146.865 77.665 ;
    END
  END r_data_o[208]
  PIN r_data_o[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 150.955 146.865 151.025 ;
    END
  END r_data_o[209]
  PIN r_data_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 143.675 146.865 143.745 ;
    END
  END r_data_o[20]
  PIN r_data_o[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  138.345 190.18 138.485 190.32 ;
    END
  END r_data_o[210]
  PIN r_data_o[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  141.705 0 141.845 0.14 ;
    END
  END r_data_o[211]
  PIN r_data_o[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 171.675 0.07 171.745 ;
    END
  END r_data_o[212]
  PIN r_data_o[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 56.035 0.07 56.105 ;
    END
  END r_data_o[213]
  PIN r_data_o[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 98.035 146.865 98.105 ;
    END
  END r_data_o[214]
  PIN r_data_o[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 124.915 0.07 124.985 ;
    END
  END r_data_o[215]
  PIN r_data_o[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  87.945 0 88.085 0.14 ;
    END
  END r_data_o[216]
  PIN r_data_o[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  70.585 0 70.725 0.14 ;
    END
  END r_data_o[217]
  PIN r_data_o[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 57.995 146.865 58.065 ;
    END
  END r_data_o[218]
  PIN r_data_o[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  55.465 190.18 55.605 190.32 ;
    END
  END r_data_o[219]
  PIN r_data_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 181.755 146.865 181.825 ;
    END
  END r_data_o[21]
  PIN r_data_o[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 165.515 0.07 165.585 ;
    END
  END r_data_o[220]
  PIN r_data_o[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 38.675 146.865 38.745 ;
    END
  END r_data_o[221]
  PIN r_data_o[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  5.065 190.18 5.205 190.32 ;
    END
  END r_data_o[222]
  PIN r_data_o[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 147.595 146.865 147.665 ;
    END
  END r_data_o[223]
  PIN r_data_o[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  119.865 0 120.005 0.14 ;
    END
  END r_data_o[224]
  PIN r_data_o[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 150.115 0.07 150.185 ;
    END
  END r_data_o[225]
  PIN r_data_o[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 92.995 146.865 93.065 ;
    END
  END r_data_o[226]
  PIN r_data_o[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  145.065 0 145.205 0.14 ;
    END
  END r_data_o[227]
  PIN r_data_o[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 81.515 146.865 81.585 ;
    END
  END r_data_o[228]
  PIN r_data_o[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  136.105 0 136.245 0.14 ;
    END
  END r_data_o[229]
  PIN r_data_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 24.395 146.865 24.465 ;
    END
  END r_data_o[22]
  PIN r_data_o[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  113.145 0 113.285 0.14 ;
    END
  END r_data_o[230]
  PIN r_data_o[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 155.435 0.07 155.505 ;
    END
  END r_data_o[231]
  PIN r_data_o[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 184.275 0.07 184.345 ;
    END
  END r_data_o[232]
  PIN r_data_o[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.945 0 32.085 0.14 ;
    END
  END r_data_o[233]
  PIN r_data_o[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 174.475 146.865 174.545 ;
    END
  END r_data_o[234]
  PIN r_data_o[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 80.115 146.865 80.185 ;
    END
  END r_data_o[235]
  PIN r_data_o[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 96.915 146.865 96.985 ;
    END
  END r_data_o[236]
  PIN r_data_o[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 187.075 146.865 187.145 ;
    END
  END r_data_o[237]
  PIN r_data_o[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 122.955 146.865 123.025 ;
    END
  END r_data_o[238]
  PIN r_data_o[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 81.235 0.07 81.305 ;
    END
  END r_data_o[239]
  PIN r_data_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 152.075 0.07 152.145 ;
    END
  END r_data_o[23]
  PIN r_data_o[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 122.955 0.07 123.025 ;
    END
  END r_data_o[240]
  PIN r_data_o[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 148.435 146.865 148.505 ;
    END
  END r_data_o[241]
  PIN r_data_o[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 24.955 0.07 25.025 ;
    END
  END r_data_o[242]
  PIN r_data_o[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  105.305 0 105.445 0.14 ;
    END
  END r_data_o[243]
  PIN r_data_o[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  74.505 190.18 74.645 190.32 ;
    END
  END r_data_o[244]
  PIN r_data_o[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  117.065 0 117.205 0.14 ;
    END
  END r_data_o[245]
  PIN r_data_o[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 115.955 0.07 116.025 ;
    END
  END r_data_o[246]
  PIN r_data_o[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  130.505 0 130.645 0.14 ;
    END
  END r_data_o[247]
  PIN r_data_o[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 167.755 0.07 167.825 ;
    END
  END r_data_o[248]
  PIN r_data_o[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 169.715 0.07 169.785 ;
    END
  END r_data_o[249]
  PIN r_data_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 45.955 146.865 46.025 ;
    END
  END r_data_o[24]
  PIN r_data_o[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 84.595 0.07 84.665 ;
    END
  END r_data_o[250]
  PIN r_data_o[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 47.355 0.07 47.425 ;
    END
  END r_data_o[251]
  PIN r_data_o[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  102.505 190.18 102.645 190.32 ;
    END
  END r_data_o[252]
  PIN r_data_o[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 97.475 146.865 97.545 ;
    END
  END r_data_o[253]
  PIN r_data_o[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 144.235 146.865 144.305 ;
    END
  END r_data_o[254]
  PIN r_data_o[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  1.145 0 1.285 0.14 ;
    END
  END r_data_o[255]
  PIN r_data_o[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 91.875 0.07 91.945 ;
    END
  END r_data_o[256]
  PIN r_data_o[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 55.195 0.07 55.265 ;
    END
  END r_data_o[257]
  PIN r_data_o[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  73.385 0 73.525 0.14 ;
    END
  END r_data_o[258]
  PIN r_data_o[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  64.985 190.18 65.125 190.32 ;
    END
  END r_data_o[259]
  PIN r_data_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  57.145 0 57.285 0.14 ;
    END
  END r_data_o[25]
  PIN r_data_o[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 70.595 146.865 70.665 ;
    END
  END r_data_o[260]
  PIN r_data_o[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  43.705 0 43.845 0.14 ;
    END
  END r_data_o[261]
  PIN r_data_o[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  74.505 0 74.645 0.14 ;
    END
  END r_data_o[262]
  PIN r_data_o[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 122.675 0.07 122.745 ;
    END
  END r_data_o[263]
  PIN r_data_o[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  90.185 190.18 90.325 190.32 ;
    END
  END r_data_o[264]
  PIN r_data_o[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 101.395 146.865 101.465 ;
    END
  END r_data_o[265]
  PIN r_data_o[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 15.715 0.07 15.785 ;
    END
  END r_data_o[266]
  PIN r_data_o[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 111.475 0.07 111.545 ;
    END
  END r_data_o[267]
  PIN r_data_o[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 66.675 146.865 66.745 ;
    END
  END r_data_o[268]
  PIN r_data_o[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.595 0.07 7.665 ;
    END
  END r_data_o[269]
  PIN r_data_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  68.905 0 69.045 0.14 ;
    END
  END r_data_o[26]
  PIN r_data_o[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 158.235 146.865 158.305 ;
    END
  END r_data_o[270]
  PIN r_data_o[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  138.905 0 139.045 0.14 ;
    END
  END r_data_o[271]
  PIN r_data_o[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 50.715 146.865 50.785 ;
    END
  END r_data_o[272]
  PIN r_data_o[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 28.595 0.07 28.665 ;
    END
  END r_data_o[273]
  PIN r_data_o[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 54.075 146.865 54.145 ;
    END
  END r_data_o[274]
  PIN r_data_o[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 132.755 0.07 132.825 ;
    END
  END r_data_o[275]
  PIN r_data_o[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 102.235 146.865 102.305 ;
    END
  END r_data_o[276]
  PIN r_data_o[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  142.265 190.18 142.405 190.32 ;
    END
  END r_data_o[277]
  PIN r_data_o[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 2.275 0.07 2.345 ;
    END
  END r_data_o[278]
  PIN r_data_o[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  32.505 190.18 32.645 190.32 ;
    END
  END r_data_o[279]
  PIN r_data_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 71.435 146.865 71.505 ;
    END
  END r_data_o[27]
  PIN r_data_o[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 79.275 0.07 79.345 ;
    END
  END r_data_o[280]
  PIN r_data_o[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 175.035 146.865 175.105 ;
    END
  END r_data_o[281]
  PIN r_data_o[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 29.715 0.07 29.785 ;
    END
  END r_data_o[282]
  PIN r_data_o[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 31.115 146.865 31.185 ;
    END
  END r_data_o[283]
  PIN r_data_o[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 35.315 0.07 35.385 ;
    END
  END r_data_o[284]
  PIN r_data_o[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 59.395 146.865 59.465 ;
    END
  END r_data_o[285]
  PIN r_data_o[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 170.275 0.07 170.345 ;
    END
  END r_data_o[286]
  PIN r_data_o[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 77.875 0.07 77.945 ;
    END
  END r_data_o[287]
  PIN r_data_o[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 13.195 0.07 13.265 ;
    END
  END r_data_o[288]
  PIN r_data_o[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 136.115 146.865 136.185 ;
    END
  END r_data_o[289]
  PIN r_data_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.115 0.07 31.185 ;
    END
  END r_data_o[28]
  PIN r_data_o[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 55.475 146.865 55.545 ;
    END
  END r_data_o[290]
  PIN r_data_o[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 112.035 0.07 112.105 ;
    END
  END r_data_o[291]
  PIN r_data_o[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 29.155 0.07 29.225 ;
    END
  END r_data_o[292]
  PIN r_data_o[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 76.475 0.07 76.545 ;
    END
  END r_data_o[293]
  PIN r_data_o[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  98.585 190.18 98.725 190.32 ;
    END
  END r_data_o[294]
  PIN r_data_o[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  1.145 190.18 1.285 190.32 ;
    END
  END r_data_o[295]
  PIN r_data_o[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  111.465 190.18 111.605 190.32 ;
    END
  END r_data_o[296]
  PIN r_data_o[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 59.115 0.07 59.185 ;
    END
  END r_data_o[297]
  PIN r_data_o[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 62.755 0.07 62.825 ;
    END
  END r_data_o[298]
  PIN r_data_o[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 182.315 0.07 182.385 ;
    END
  END r_data_o[299]
  PIN r_data_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 105.035 146.865 105.105 ;
    END
  END r_data_o[29]
  PIN r_data_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 9.835 146.865 9.905 ;
    END
  END r_data_o[2]
  PIN r_data_o[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 1.995 146.865 2.065 ;
    END
  END r_data_o[300]
  PIN r_data_o[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 92.155 146.865 92.225 ;
    END
  END r_data_o[301]
  PIN r_data_o[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 144.795 0.07 144.865 ;
    END
  END r_data_o[302]
  PIN r_data_o[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 109.515 146.865 109.585 ;
    END
  END r_data_o[303]
  PIN r_data_o[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 5.355 146.865 5.425 ;
    END
  END r_data_o[304]
  PIN r_data_o[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  77.305 0 77.445 0.14 ;
    END
  END r_data_o[305]
  PIN r_data_o[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 93.555 0.07 93.625 ;
    END
  END r_data_o[306]
  PIN r_data_o[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 26.635 146.865 26.705 ;
    END
  END r_data_o[307]
  PIN r_data_o[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 78.155 146.865 78.225 ;
    END
  END r_data_o[308]
  PIN r_data_o[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 147.035 0.07 147.105 ;
    END
  END r_data_o[309]
  PIN r_data_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 42.035 146.865 42.105 ;
    END
  END r_data_o[30]
  PIN r_data_o[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 88.795 146.865 88.865 ;
    END
  END r_data_o[310]
  PIN r_data_o[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 106.155 146.865 106.225 ;
    END
  END r_data_o[311]
  PIN r_data_o[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 61.915 0.07 61.985 ;
    END
  END r_data_o[312]
  PIN r_data_o[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 176.995 146.865 177.065 ;
    END
  END r_data_o[313]
  PIN r_data_o[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  123.785 190.18 123.925 190.32 ;
    END
  END r_data_o[314]
  PIN r_data_o[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 42.595 0.07 42.665 ;
    END
  END r_data_o[315]
  PIN r_data_o[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 95.515 0.07 95.585 ;
    END
  END r_data_o[316]
  PIN r_data_o[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 116.235 0.07 116.305 ;
    END
  END r_data_o[317]
  PIN r_data_o[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 112.875 146.865 112.945 ;
    END
  END r_data_o[318]
  PIN r_data_o[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 122.115 146.865 122.185 ;
    END
  END r_data_o[319]
  PIN r_data_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 113.435 146.865 113.505 ;
    END
  END r_data_o[31]
  PIN r_data_o[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 187.075 0.07 187.145 ;
    END
  END r_data_o[320]
  PIN r_data_o[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 68.075 0.07 68.145 ;
    END
  END r_data_o[321]
  PIN r_data_o[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 134.715 0.07 134.785 ;
    END
  END r_data_o[322]
  PIN r_data_o[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 175.595 146.865 175.665 ;
    END
  END r_data_o[323]
  PIN r_data_o[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  133.305 0 133.445 0.14 ;
    END
  END r_data_o[324]
  PIN r_data_o[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 105.595 0.07 105.665 ;
    END
  END r_data_o[325]
  PIN r_data_o[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  135.545 190.18 135.685 190.32 ;
    END
  END r_data_o[326]
  PIN r_data_o[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 94.675 146.865 94.745 ;
    END
  END r_data_o[327]
  PIN r_data_o[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  22.425 0 22.565 0.14 ;
    END
  END r_data_o[328]
  PIN r_data_o[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 179.515 0.07 179.585 ;
    END
  END r_data_o[329]
  PIN r_data_o[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 10.955 0.07 11.025 ;
    END
  END r_data_o[32]
  PIN r_data_o[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 123.515 0.07 123.585 ;
    END
  END r_data_o[330]
  PIN r_data_o[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  122.665 0 122.805 0.14 ;
    END
  END r_data_o[331]
  PIN r_data_o[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  143.945 0 144.085 0.14 ;
    END
  END r_data_o[332]
  PIN r_data_o[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 117.635 146.865 117.705 ;
    END
  END r_data_o[333]
  PIN r_data_o[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 47.915 146.865 47.985 ;
    END
  END r_data_o[334]
  PIN r_data_o[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 179.795 146.865 179.865 ;
    END
  END r_data_o[335]
  PIN r_data_o[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 112.875 0.07 112.945 ;
    END
  END r_data_o[336]
  PIN r_data_o[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 79.555 146.865 79.625 ;
    END
  END r_data_o[337]
  PIN r_data_o[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 156.275 146.865 156.345 ;
    END
  END r_data_o[338]
  PIN r_data_o[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 161.035 146.865 161.105 ;
    END
  END r_data_o[339]
  PIN r_data_o[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 41.195 0.07 41.265 ;
    END
  END r_data_o[33]
  PIN r_data_o[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 63.875 0.07 63.945 ;
    END
  END r_data_o[340]
  PIN r_data_o[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  76.745 190.18 76.885 190.32 ;
    END
  END r_data_o[341]
  PIN r_data_o[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  118.745 190.18 118.885 190.32 ;
    END
  END r_data_o[342]
  PIN r_data_o[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.305 190.18 7.445 190.32 ;
    END
  END r_data_o[343]
  PIN r_data_o[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 119.315 0.07 119.385 ;
    END
  END r_data_o[344]
  PIN r_data_o[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 172.515 146.865 172.585 ;
    END
  END r_data_o[345]
  PIN r_data_o[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 97.475 0.07 97.545 ;
    END
  END r_data_o[346]
  PIN r_data_o[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 174.475 0.07 174.545 ;
    END
  END r_data_o[347]
  PIN r_data_o[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 175.595 0.07 175.665 ;
    END
  END r_data_o[348]
  PIN r_data_o[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  15.705 190.18 15.845 190.32 ;
    END
  END r_data_o[349]
  PIN r_data_o[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 87.955 0.07 88.025 ;
    END
  END r_data_o[34]
  PIN r_data_o[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 39.235 146.865 39.305 ;
    END
  END r_data_o[350]
  PIN r_data_o[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 121.555 146.865 121.625 ;
    END
  END r_data_o[351]
  PIN r_data_o[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 8.995 0.07 9.065 ;
    END
  END r_data_o[352]
  PIN r_data_o[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 132.755 146.865 132.825 ;
    END
  END r_data_o[353]
  PIN r_data_o[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 51.275 146.865 51.345 ;
    END
  END r_data_o[354]
  PIN r_data_o[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 180.915 0.07 180.985 ;
    END
  END r_data_o[355]
  PIN r_data_o[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 101.395 0.07 101.465 ;
    END
  END r_data_o[356]
  PIN r_data_o[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 96.075 146.865 96.145 ;
    END
  END r_data_o[357]
  PIN r_data_o[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 55.755 0.07 55.825 ;
    END
  END r_data_o[358]
  PIN r_data_o[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 30.555 146.865 30.625 ;
    END
  END r_data_o[359]
  PIN r_data_o[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 106.715 146.865 106.785 ;
    END
  END r_data_o[35]
  PIN r_data_o[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 19.915 0.07 19.985 ;
    END
  END r_data_o[360]
  PIN r_data_o[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 158.515 146.865 158.585 ;
    END
  END r_data_o[361]
  PIN r_data_o[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  70.025 190.18 70.165 190.32 ;
    END
  END r_data_o[362]
  PIN r_data_o[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 49.315 146.865 49.385 ;
    END
  END r_data_o[363]
  PIN r_data_o[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  95.785 190.18 95.925 190.32 ;
    END
  END r_data_o[364]
  PIN r_data_o[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  117.065 190.18 117.205 190.32 ;
    END
  END r_data_o[365]
  PIN r_data_o[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  4.505 190.18 4.645 190.32 ;
    END
  END r_data_o[366]
  PIN r_data_o[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  97.465 0 97.605 0.14 ;
    END
  END r_data_o[367]
  PIN r_data_o[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 126.875 0.07 126.945 ;
    END
  END r_data_o[368]
  PIN r_data_o[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 45.395 0.07 45.465 ;
    END
  END r_data_o[369]
  PIN r_data_o[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 17.675 0.07 17.745 ;
    END
  END r_data_o[36]
  PIN r_data_o[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  29.145 190.18 29.285 190.32 ;
    END
  END r_data_o[370]
  PIN r_data_o[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 143.395 0.07 143.465 ;
    END
  END r_data_o[371]
  PIN r_data_o[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 179.795 0.07 179.865 ;
    END
  END r_data_o[372]
  PIN r_data_o[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 99.435 146.865 99.505 ;
    END
  END r_data_o[373]
  PIN r_data_o[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  141.145 190.18 141.285 190.32 ;
    END
  END r_data_o[374]
  PIN r_data_o[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 104.755 0.07 104.825 ;
    END
  END r_data_o[375]
  PIN r_data_o[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 104.195 146.865 104.265 ;
    END
  END r_data_o[376]
  PIN r_data_o[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 12.355 146.865 12.425 ;
    END
  END r_data_o[377]
  PIN r_data_o[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 91.315 146.865 91.385 ;
    END
  END r_data_o[378]
  PIN r_data_o[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 187.635 0.07 187.705 ;
    END
  END r_data_o[379]
  PIN r_data_o[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  122.665 190.18 122.805 190.32 ;
    END
  END r_data_o[37]
  PIN r_data_o[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 183.155 0.07 183.225 ;
    END
  END r_data_o[380]
  PIN r_data_o[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  85.145 0 85.285 0.14 ;
    END
  END r_data_o[381]
  PIN r_data_o[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 22.435 0.07 22.505 ;
    END
  END r_data_o[382]
  PIN r_data_o[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 124.075 0.07 124.145 ;
    END
  END r_data_o[383]
  PIN r_data_o[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  127.705 0 127.845 0.14 ;
    END
  END r_data_o[384]
  PIN r_data_o[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 68.635 0.07 68.705 ;
    END
  END r_data_o[385]
  PIN r_data_o[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 165.795 0.07 165.865 ;
    END
  END r_data_o[386]
  PIN r_data_o[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 138.915 146.865 138.985 ;
    END
  END r_data_o[387]
  PIN r_data_o[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 170.835 0.07 170.905 ;
    END
  END r_data_o[388]
  PIN r_data_o[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 4.235 0.07 4.305 ;
    END
  END r_data_o[389]
  PIN r_data_o[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 187.915 146.865 187.985 ;
    END
  END r_data_o[38]
  PIN r_data_o[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  86.265 190.18 86.405 190.32 ;
    END
  END r_data_o[390]
  PIN r_data_o[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 171.675 146.865 171.745 ;
    END
  END r_data_o[391]
  PIN r_data_o[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 138.355 146.865 138.425 ;
    END
  END r_data_o[392]
  PIN r_data_o[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 99.995 0.07 100.065 ;
    END
  END r_data_o[393]
  PIN r_data_o[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 119.595 0.07 119.665 ;
    END
  END r_data_o[394]
  PIN r_data_o[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  82.345 0 82.485 0.14 ;
    END
  END r_data_o[395]
  PIN r_data_o[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 167.755 146.865 167.825 ;
    END
  END r_data_o[396]
  PIN r_data_o[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  92.985 190.18 93.125 190.32 ;
    END
  END r_data_o[397]
  PIN r_data_o[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 124.355 146.865 124.425 ;
    END
  END r_data_o[398]
  PIN r_data_o[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  115.945 190.18 116.085 190.32 ;
    END
  END r_data_o[399]
  PIN r_data_o[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 65.275 0.07 65.345 ;
    END
  END r_data_o[39]
  PIN r_data_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 148.155 0.07 148.225 ;
    END
  END r_data_o[3]
  PIN r_data_o[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 142.835 146.865 142.905 ;
    END
  END r_data_o[400]
  PIN r_data_o[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 33.915 146.865 33.985 ;
    END
  END r_data_o[401]
  PIN r_data_o[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 105.595 146.865 105.665 ;
    END
  END r_data_o[402]
  PIN r_data_o[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  110.345 0 110.485 0.14 ;
    END
  END r_data_o[403]
  PIN r_data_o[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 39.795 146.865 39.865 ;
    END
  END r_data_o[404]
  PIN r_data_o[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 29.155 146.865 29.225 ;
    END
  END r_data_o[405]
  PIN r_data_o[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.385 0 31.525 0.14 ;
    END
  END r_data_o[406]
  PIN r_data_o[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 71.155 0.07 71.225 ;
    END
  END r_data_o[407]
  PIN r_data_o[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 130.795 146.865 130.865 ;
    END
  END r_data_o[408]
  PIN r_data_o[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  125.465 0 125.605 0.14 ;
    END
  END r_data_o[409]
  PIN r_data_o[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 41.755 0.07 41.825 ;
    END
  END r_data_o[40]
  PIN r_data_o[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  71.705 0 71.845 0.14 ;
    END
  END r_data_o[410]
  PIN r_data_o[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 15.155 0.07 15.225 ;
    END
  END r_data_o[411]
  PIN r_data_o[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 96.635 0.07 96.705 ;
    END
  END r_data_o[412]
  PIN r_data_o[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  20.745 190.18 20.885 190.32 ;
    END
  END r_data_o[413]
  PIN r_data_o[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 16.275 0.07 16.345 ;
    END
  END r_data_o[414]
  PIN r_data_o[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 54.635 0.07 54.705 ;
    END
  END r_data_o[415]
  PIN r_data_o[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 92.155 0.07 92.225 ;
    END
  END r_data_o[416]
  PIN r_data_o[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 81.515 0.07 81.585 ;
    END
  END r_data_o[417]
  PIN r_data_o[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  143.945 190.18 144.085 190.32 ;
    END
  END r_data_o[418]
  PIN r_data_o[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 58.555 0.07 58.625 ;
    END
  END r_data_o[419]
  PIN r_data_o[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 162.995 146.865 163.065 ;
    END
  END r_data_o[41]
  PIN r_data_o[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 90.195 146.865 90.265 ;
    END
  END r_data_o[420]
  PIN r_data_o[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 134.155 0.07 134.225 ;
    END
  END r_data_o[421]
  PIN r_data_o[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 178.955 146.865 179.025 ;
    END
  END r_data_o[422]
  PIN r_data_o[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 68.635 146.865 68.705 ;
    END
  END r_data_o[423]
  PIN r_data_o[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 33.355 0.07 33.425 ;
    END
  END r_data_o[424]
  PIN r_data_o[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  44.825 0 44.965 0.14 ;
    END
  END r_data_o[425]
  PIN r_data_o[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 40.635 146.865 40.705 ;
    END
  END r_data_o[426]
  PIN r_data_o[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 166.355 0.07 166.425 ;
    END
  END r_data_o[427]
  PIN r_data_o[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  129.385 190.18 129.525 190.32 ;
    END
  END r_data_o[428]
  PIN r_data_o[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 185.115 0.07 185.185 ;
    END
  END r_data_o[429]
  PIN r_data_o[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 29.435 146.865 29.505 ;
    END
  END r_data_o[42]
  PIN r_data_o[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 70.035 146.865 70.105 ;
    END
  END r_data_o[430]
  PIN r_data_o[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 157.675 146.865 157.745 ;
    END
  END r_data_o[431]
  PIN r_data_o[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 30.555 0.07 30.625 ;
    END
  END r_data_o[432]
  PIN r_data_o[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 32.515 146.865 32.585 ;
    END
  END r_data_o[433]
  PIN r_data_o[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  39.225 190.18 39.365 190.32 ;
    END
  END r_data_o[434]
  PIN r_data_o[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  94.105 190.18 94.245 190.32 ;
    END
  END r_data_o[435]
  PIN r_data_o[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 126.875 146.865 126.945 ;
    END
  END r_data_o[436]
  PIN r_data_o[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 175.035 0.07 175.105 ;
    END
  END r_data_o[437]
  PIN r_data_o[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 98.875 146.865 98.945 ;
    END
  END r_data_o[438]
  PIN r_data_o[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 145.635 146.865 145.705 ;
    END
  END r_data_o[439]
  PIN r_data_o[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 37.275 0.07 37.345 ;
    END
  END r_data_o[43]
  PIN r_data_o[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  58.825 0 58.965 0.14 ;
    END
  END r_data_o[440]
  PIN r_data_o[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 159.635 146.865 159.705 ;
    END
  END r_data_o[441]
  PIN r_data_o[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  19.625 190.18 19.765 190.32 ;
    END
  END r_data_o[442]
  PIN r_data_o[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 47.075 0.07 47.145 ;
    END
  END r_data_o[443]
  PIN r_data_o[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 85.995 146.865 86.065 ;
    END
  END r_data_o[444]
  PIN r_data_o[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 14.595 0.07 14.665 ;
    END
  END r_data_o[445]
  PIN r_data_o[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 165.795 146.865 165.865 ;
    END
  END r_data_o[446]
  PIN r_data_o[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 101.675 146.865 101.745 ;
    END
  END r_data_o[447]
  PIN r_data_o[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 44.555 146.865 44.625 ;
    END
  END r_data_o[448]
  PIN r_data_o[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 49.875 0.07 49.945 ;
    END
  END r_data_o[449]
  PIN r_data_o[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 173.075 146.865 173.145 ;
    END
  END r_data_o[44]
  PIN r_data_o[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  98.585 0 98.725 0.14 ;
    END
  END r_data_o[450]
  PIN r_data_o[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  16.825 0 16.965 0.14 ;
    END
  END r_data_o[451]
  PIN r_data_o[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 74.795 0.07 74.865 ;
    END
  END r_data_o[452]
  PIN r_data_o[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 107.275 0.07 107.345 ;
    END
  END r_data_o[453]
  PIN r_data_o[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 94.115 0.07 94.185 ;
    END
  END r_data_o[454]
  PIN r_data_o[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 189.035 0.07 189.105 ;
    END
  END r_data_o[455]
  PIN r_data_o[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.035 0.07 21.105 ;
    END
  END r_data_o[456]
  PIN r_data_o[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 113.995 0.07 114.065 ;
    END
  END r_data_o[457]
  PIN r_data_o[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 85.155 0.07 85.225 ;
    END
  END r_data_o[458]
  PIN r_data_o[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 42.035 0.07 42.105 ;
    END
  END r_data_o[459]
  PIN r_data_o[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 153.755 0.07 153.825 ;
    END
  END r_data_o[45]
  PIN r_data_o[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 57.435 0.07 57.505 ;
    END
  END r_data_o[460]
  PIN r_data_o[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 121.275 0.07 121.345 ;
    END
  END r_data_o[461]
  PIN r_data_o[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 120.715 0.07 120.785 ;
    END
  END r_data_o[462]
  PIN r_data_o[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 25.795 0.07 25.865 ;
    END
  END r_data_o[463]
  PIN r_data_o[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 129.675 0.07 129.745 ;
    END
  END r_data_o[464]
  PIN r_data_o[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 77.315 146.865 77.385 ;
    END
  END r_data_o[465]
  PIN r_data_o[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 128.275 146.865 128.345 ;
    END
  END r_data_o[466]
  PIN r_data_o[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 17.955 0.07 18.025 ;
    END
  END r_data_o[467]
  PIN r_data_o[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 188.475 0.07 188.545 ;
    END
  END r_data_o[468]
  PIN r_data_o[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  69.465 0 69.605 0.14 ;
    END
  END r_data_o[469]
  PIN r_data_o[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 67.235 146.865 67.305 ;
    END
  END r_data_o[46]
  PIN r_data_o[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 122.395 146.865 122.465 ;
    END
  END r_data_o[470]
  PIN r_data_o[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 114.275 0.07 114.345 ;
    END
  END r_data_o[471]
  PIN r_data_o[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  124.345 0 124.485 0.14 ;
    END
  END r_data_o[472]
  PIN r_data_o[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 36.435 0.07 36.505 ;
    END
  END r_data_o[473]
  PIN r_data_o[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  38.105 0 38.245 0.14 ;
    END
  END r_data_o[474]
  PIN r_data_o[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 154.315 146.865 154.385 ;
    END
  END r_data_o[475]
  PIN r_data_o[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  36.985 0 37.125 0.14 ;
    END
  END r_data_o[476]
  PIN r_data_o[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 106.715 0.07 106.785 ;
    END
  END r_data_o[477]
  PIN r_data_o[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  137.785 0 137.925 0.14 ;
    END
  END r_data_o[478]
  PIN r_data_o[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  18.505 190.18 18.645 190.32 ;
    END
  END r_data_o[479]
  PIN r_data_o[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  48.745 0 48.885 0.14 ;
    END
  END r_data_o[47]
  PIN r_data_o[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 137.515 146.865 137.585 ;
    END
  END r_data_o[480]
  PIN r_data_o[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  64.985 0 65.125 0.14 ;
    END
  END r_data_o[481]
  PIN r_data_o[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 177.835 0.07 177.905 ;
    END
  END r_data_o[482]
  PIN r_data_o[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 161.035 0.07 161.105 ;
    END
  END r_data_o[483]
  PIN r_data_o[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 174.195 0.07 174.265 ;
    END
  END r_data_o[484]
  PIN r_data_o[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  19.625 0 19.765 0.14 ;
    END
  END r_data_o[485]
  PIN r_data_o[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 168.315 146.865 168.385 ;
    END
  END r_data_o[486]
  PIN r_data_o[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 33.075 0.07 33.145 ;
    END
  END r_data_o[487]
  PIN r_data_o[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 55.195 146.865 55.265 ;
    END
  END r_data_o[488]
  PIN r_data_o[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 18.515 146.865 18.585 ;
    END
  END r_data_o[489]
  PIN r_data_o[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 62.475 0.07 62.545 ;
    END
  END r_data_o[48]
  PIN r_data_o[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 152.915 0.07 152.985 ;
    END
  END r_data_o[490]
  PIN r_data_o[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 82.635 146.865 82.705 ;
    END
  END r_data_o[491]
  PIN r_data_o[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 13.755 0.07 13.825 ;
    END
  END r_data_o[492]
  PIN r_data_o[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 129.115 146.865 129.185 ;
    END
  END r_data_o[493]
  PIN r_data_o[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  112.025 190.18 112.165 190.32 ;
    END
  END r_data_o[494]
  PIN r_data_o[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  118.745 0 118.885 0.14 ;
    END
  END r_data_o[495]
  PIN r_data_o[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 144.795 146.865 144.865 ;
    END
  END r_data_o[496]
  PIN r_data_o[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 171.115 0.07 171.185 ;
    END
  END r_data_o[497]
  PIN r_data_o[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  78.425 0 78.565 0.14 ;
    END
  END r_data_o[498]
  PIN r_data_o[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 147.035 146.865 147.105 ;
    END
  END r_data_o[499]
  PIN r_data_o[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 162.435 146.865 162.505 ;
    END
  END r_data_o[49]
  PIN r_data_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 163.835 146.865 163.905 ;
    END
  END r_data_o[4]
  PIN r_data_o[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  84.025 190.18 84.165 190.32 ;
    END
  END r_data_o[500]
  PIN r_data_o[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  108.105 0 108.245 0.14 ;
    END
  END r_data_o[501]
  PIN r_data_o[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  44.825 190.18 44.965 190.32 ;
    END
  END r_data_o[502]
  PIN r_data_o[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 169.435 0.07 169.505 ;
    END
  END r_data_o[503]
  PIN r_data_o[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 86.555 0.07 86.625 ;
    END
  END r_data_o[504]
  PIN r_data_o[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  63.305 190.18 63.445 190.32 ;
    END
  END r_data_o[505]
  PIN r_data_o[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 181.195 146.865 181.265 ;
    END
  END r_data_o[506]
  PIN r_data_o[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 178.395 0.07 178.465 ;
    END
  END r_data_o[507]
  PIN r_data_o[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 29.995 0.07 30.065 ;
    END
  END r_data_o[508]
  PIN r_data_o[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 80.675 146.865 80.745 ;
    END
  END r_data_o[509]
  PIN r_data_o[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 21.875 146.865 21.945 ;
    END
  END r_data_o[50]
  PIN r_data_o[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 161.595 0.07 161.665 ;
    END
  END r_data_o[510]
  PIN r_data_o[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 1.715 0.07 1.785 ;
    END
  END r_data_o[511]
  PIN r_data_o[512]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 92.715 0.07 92.785 ;
    END
  END r_data_o[512]
  PIN r_data_o[513]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  81.225 0 81.365 0.14 ;
    END
  END r_data_o[513]
  PIN r_data_o[514]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  36.985 190.18 37.125 190.32 ;
    END
  END r_data_o[514]
  PIN r_data_o[515]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  40.905 190.18 41.045 190.32 ;
    END
  END r_data_o[515]
  PIN r_data_o[516]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 93.275 0.07 93.345 ;
    END
  END r_data_o[516]
  PIN r_data_o[517]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 138.355 0.07 138.425 ;
    END
  END r_data_o[517]
  PIN r_data_o[518]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 135.555 0.07 135.625 ;
    END
  END r_data_o[518]
  PIN r_data_o[519]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 136.955 0.07 137.025 ;
    END
  END r_data_o[519]
  PIN r_data_o[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 170.555 146.865 170.625 ;
    END
  END r_data_o[51]
  PIN r_data_o[520]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 136.115 0.07 136.185 ;
    END
  END r_data_o[520]
  PIN r_data_o[521]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 69.195 0.07 69.265 ;
    END
  END r_data_o[521]
  PIN r_data_o[522]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 169.715 146.865 169.785 ;
    END
  END r_data_o[522]
  PIN r_data_o[523]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 9.275 0.07 9.345 ;
    END
  END r_data_o[523]
  PIN r_data_o[524]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  100.825 190.18 100.965 190.32 ;
    END
  END r_data_o[524]
  PIN r_data_o[525]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 45.395 146.865 45.465 ;
    END
  END r_data_o[525]
  PIN r_data_o[526]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.675 0.07 31.745 ;
    END
  END r_data_o[526]
  PIN r_data_o[527]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 151.515 146.865 151.585 ;
    END
  END r_data_o[527]
  PIN r_data_o[528]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  66.665 190.18 66.805 190.32 ;
    END
  END r_data_o[528]
  PIN r_data_o[529]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 176.435 146.865 176.505 ;
    END
  END r_data_o[529]
  PIN r_data_o[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 106.155 0.07 106.225 ;
    END
  END r_data_o[52]
  PIN r_data_o[530]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  132.185 190.18 132.325 190.32 ;
    END
  END r_data_o[530]
  PIN r_data_o[531]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 89.635 146.865 89.705 ;
    END
  END r_data_o[531]
  PIN r_data_o[532]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 53.235 146.865 53.305 ;
    END
  END r_data_o[532]
  PIN r_data_o[533]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 88.795 0.07 88.865 ;
    END
  END r_data_o[533]
  PIN r_data_o[534]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 73.955 0.07 74.025 ;
    END
  END r_data_o[534]
  PIN r_data_o[535]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  90.745 0 90.885 0.14 ;
    END
  END r_data_o[535]
  PIN r_data_o[536]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  24.665 0 24.805 0.14 ;
    END
  END r_data_o[536]
  PIN r_data_o[537]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 125.475 146.865 125.545 ;
    END
  END r_data_o[537]
  PIN r_data_o[538]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  39.785 0 39.925 0.14 ;
    END
  END r_data_o[538]
  PIN r_data_o[539]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 35.315 146.865 35.385 ;
    END
  END r_data_o[539]
  PIN r_data_o[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  21.865 190.18 22.005 190.32 ;
    END
  END r_data_o[53]
  PIN r_data_o[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 24.395 0.07 24.465 ;
    END
  END r_data_o[54]
  PIN r_data_o[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  102.505 0 102.645 0.14 ;
    END
  END r_data_o[55]
  PIN r_data_o[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  128.265 0 128.405 0.14 ;
    END
  END r_data_o[56]
  PIN r_data_o[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 110.915 146.865 110.985 ;
    END
  END r_data_o[57]
  PIN r_data_o[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 124.915 146.865 124.985 ;
    END
  END r_data_o[58]
  PIN r_data_o[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 52.675 146.865 52.745 ;
    END
  END r_data_o[59]
  PIN r_data_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  142.825 190.18 142.965 190.32 ;
    END
  END r_data_o[5]
  PIN r_data_o[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  61.065 0 61.205 0.14 ;
    END
  END r_data_o[60]
  PIN r_data_o[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 185.675 146.865 185.745 ;
    END
  END r_data_o[61]
  PIN r_data_o[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 14.595 146.865 14.665 ;
    END
  END r_data_o[62]
  PIN r_data_o[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 176.155 0.07 176.225 ;
    END
  END r_data_o[63]
  PIN r_data_o[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 126.315 146.865 126.385 ;
    END
  END r_data_o[64]
  PIN r_data_o[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  18.505 0 18.645 0.14 ;
    END
  END r_data_o[65]
  PIN r_data_o[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 46.515 0.07 46.585 ;
    END
  END r_data_o[66]
  PIN r_data_o[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  121.545 0 121.685 0.14 ;
    END
  END r_data_o[67]
  PIN r_data_o[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.585 0 14.725 0.14 ;
    END
  END r_data_o[68]
  PIN r_data_o[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 137.795 146.865 137.865 ;
    END
  END r_data_o[69]
  PIN r_data_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 3.675 0.07 3.745 ;
    END
  END r_data_o[6]
  PIN r_data_o[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 133.595 146.865 133.665 ;
    END
  END r_data_o[70]
  PIN r_data_o[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  141.145 0 141.285 0.14 ;
    END
  END r_data_o[71]
  PIN r_data_o[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 130.235 0.07 130.305 ;
    END
  END r_data_o[72]
  PIN r_data_o[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 99.435 0.07 99.505 ;
    END
  END r_data_o[73]
  PIN r_data_o[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  76.185 0 76.325 0.14 ;
    END
  END r_data_o[74]
  PIN r_data_o[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 43.155 146.865 43.225 ;
    END
  END r_data_o[75]
  PIN r_data_o[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  89.065 190.18 89.205 190.32 ;
    END
  END r_data_o[76]
  PIN r_data_o[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.385 0 17.525 0.14 ;
    END
  END r_data_o[77]
  PIN r_data_o[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 87.395 0.07 87.465 ;
    END
  END r_data_o[78]
  PIN r_data_o[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 71.995 146.865 72.065 ;
    END
  END r_data_o[79]
  PIN r_data_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 61.075 0.07 61.145 ;
    END
  END r_data_o[7]
  PIN r_data_o[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.875 0.07 21.945 ;
    END
  END r_data_o[80]
  PIN r_data_o[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 72.835 146.865 72.905 ;
    END
  END r_data_o[81]
  PIN r_data_o[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  96.905 190.18 97.045 190.32 ;
    END
  END r_data_o[82]
  PIN r_data_o[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  15.145 190.18 15.285 190.32 ;
    END
  END r_data_o[83]
  PIN r_data_o[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 13.195 146.865 13.265 ;
    END
  END r_data_o[84]
  PIN r_data_o[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 151.795 146.865 151.865 ;
    END
  END r_data_o[85]
  PIN r_data_o[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  33.065 190.18 33.205 190.32 ;
    END
  END r_data_o[86]
  PIN r_data_o[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  83.465 190.18 83.605 190.32 ;
    END
  END r_data_o[87]
  PIN r_data_o[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 130.235 146.865 130.305 ;
    END
  END r_data_o[88]
  PIN r_data_o[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 28.595 146.865 28.665 ;
    END
  END r_data_o[89]
  PIN r_data_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 106.995 146.865 107.065 ;
    END
  END r_data_o[8]
  PIN r_data_o[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  35.865 0 36.005 0.14 ;
    END
  END r_data_o[90]
  PIN r_data_o[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 94.115 146.865 94.185 ;
    END
  END r_data_o[91]
  PIN r_data_o[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 117.355 0.07 117.425 ;
    END
  END r_data_o[92]
  PIN r_data_o[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 133.035 146.865 133.105 ;
    END
  END r_data_o[93]
  PIN r_data_o[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 89.355 146.865 89.425 ;
    END
  END r_data_o[94]
  PIN r_data_o[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 56.875 146.865 56.945 ;
    END
  END r_data_o[95]
  PIN r_data_o[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  2.265 0 2.405 0.14 ;
    END
  END r_data_o[96]
  PIN r_data_o[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 60.515 146.865 60.585 ;
    END
  END r_data_o[97]
  PIN r_data_o[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 57.155 0.07 57.225 ;
    END
  END r_data_o[98]
  PIN r_data_o[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 165.235 146.865 165.305 ;
    END
  END r_data_o[99]
  PIN r_data_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 86.835 146.865 86.905 ;
    END
  END r_data_o[9]
  PIN r_v_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 173.075 0.07 173.145 ;
    END
  END r_v_i
  PIN w_addr_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 108.115 0.07 108.185 ;
    END
  END w_addr_i
  PIN w_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  8.985 190.18 9.125 190.32 ;
    END
  END w_clk_i
  PIN w_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 120.155 0.07 120.225 ;
    END
  END w_data_i[0]
  PIN w_data_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 164.115 0.07 164.185 ;
    END
  END w_data_i[100]
  PIN w_data_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 5.915 146.865 5.985 ;
    END
  END w_data_i[101]
  PIN w_data_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 5.075 146.865 5.145 ;
    END
  END w_data_i[102]
  PIN w_data_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 157.675 0.07 157.745 ;
    END
  END w_data_i[103]
  PIN w_data_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 22.715 146.865 22.785 ;
    END
  END w_data_i[104]
  PIN w_data_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 74.515 0.07 74.585 ;
    END
  END w_data_i[105]
  PIN w_data_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 51.835 0.07 51.905 ;
    END
  END w_data_i[106]
  PIN w_data_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  72.825 0 72.965 0.14 ;
    END
  END w_data_i[107]
  PIN w_data_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 113.715 146.865 113.785 ;
    END
  END w_data_i[108]
  PIN w_data_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 103.915 0.07 103.985 ;
    END
  END w_data_i[109]
  PIN w_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  16.825 190.18 16.965 190.32 ;
    END
  END w_data_i[10]
  PIN w_data_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 14.035 146.865 14.105 ;
    END
  END w_data_i[110]
  PIN w_data_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 163.555 146.865 163.625 ;
    END
  END w_data_i[111]
  PIN w_data_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 7.315 146.865 7.385 ;
    END
  END w_data_i[112]
  PIN w_data_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 67.515 146.865 67.585 ;
    END
  END w_data_i[113]
  PIN w_data_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  59.385 190.18 59.525 190.32 ;
    END
  END w_data_i[114]
  PIN w_data_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  75.625 0 75.765 0.14 ;
    END
  END w_data_i[115]
  PIN w_data_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 24.675 146.865 24.745 ;
    END
  END w_data_i[116]
  PIN w_data_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  131.625 190.18 131.765 190.32 ;
    END
  END w_data_i[117]
  PIN w_data_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 166.915 0.07 166.985 ;
    END
  END w_data_i[118]
  PIN w_data_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 163.555 0.07 163.625 ;
    END
  END w_data_i[119]
  PIN w_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 139.475 0.07 139.545 ;
    END
  END w_data_i[11]
  PIN w_data_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  53.225 0 53.365 0.14 ;
    END
  END w_data_i[120]
  PIN w_data_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 143.675 0.07 143.745 ;
    END
  END w_data_i[121]
  PIN w_data_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 84.035 146.865 84.105 ;
    END
  END w_data_i[122]
  PIN w_data_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 183.715 146.865 183.785 ;
    END
  END w_data_i[123]
  PIN w_data_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 142.835 0.07 142.905 ;
    END
  END w_data_i[124]
  PIN w_data_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 65.835 0.07 65.905 ;
    END
  END w_data_i[125]
  PIN w_data_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 109.515 0.07 109.585 ;
    END
  END w_data_i[126]
  PIN w_data_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 36.715 146.865 36.785 ;
    END
  END w_data_i[127]
  PIN w_data_i[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 16.555 0.07 16.625 ;
    END
  END w_data_i[128]
  PIN w_data_i[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 31.395 146.865 31.465 ;
    END
  END w_data_i[129]
  PIN w_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  93.545 0 93.685 0.14 ;
    END
  END w_data_i[12]
  PIN w_data_i[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 62.755 146.865 62.825 ;
    END
  END w_data_i[130]
  PIN w_data_i[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 127.435 0.07 127.505 ;
    END
  END w_data_i[131]
  PIN w_data_i[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  57.145 190.18 57.285 190.32 ;
    END
  END w_data_i[132]
  PIN w_data_i[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 166.355 146.865 166.425 ;
    END
  END w_data_i[133]
  PIN w_data_i[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  106.985 0 107.125 0.14 ;
    END
  END w_data_i[134]
  PIN w_data_i[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 35.875 146.865 35.945 ;
    END
  END w_data_i[135]
  PIN w_data_i[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 131.635 0.07 131.705 ;
    END
  END w_data_i[136]
  PIN w_data_i[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 82.635 0.07 82.705 ;
    END
  END w_data_i[137]
  PIN w_data_i[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  42.585 0 42.725 0.14 ;
    END
  END w_data_i[138]
  PIN w_data_i[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 169.155 146.865 169.225 ;
    END
  END w_data_i[139]
  PIN w_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  113.145 190.18 113.285 190.32 ;
    END
  END w_data_i[13]
  PIN w_data_i[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  94.665 190.18 94.805 190.32 ;
    END
  END w_data_i[140]
  PIN w_data_i[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 90.755 146.865 90.825 ;
    END
  END w_data_i[141]
  PIN w_data_i[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 34.475 0.07 34.545 ;
    END
  END w_data_i[142]
  PIN w_data_i[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 133.595 0.07 133.665 ;
    END
  END w_data_i[143]
  PIN w_data_i[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 50.155 146.865 50.225 ;
    END
  END w_data_i[144]
  PIN w_data_i[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 22.435 146.865 22.505 ;
    END
  END w_data_i[145]
  PIN w_data_i[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  136.105 190.18 136.245 190.32 ;
    END
  END w_data_i[146]
  PIN w_data_i[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  121.545 190.18 121.685 190.32 ;
    END
  END w_data_i[147]
  PIN w_data_i[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  8.985 0 9.125 0.14 ;
    END
  END w_data_i[148]
  PIN w_data_i[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 88.515 0.07 88.585 ;
    END
  END w_data_i[149]
  PIN w_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 34.755 146.865 34.825 ;
    END
  END w_data_i[14]
  PIN w_data_i[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 11.795 0.07 11.865 ;
    END
  END w_data_i[150]
  PIN w_data_i[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  45.945 190.18 46.085 190.32 ;
    END
  END w_data_i[151]
  PIN w_data_i[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 5.075 0.07 5.145 ;
    END
  END w_data_i[152]
  PIN w_data_i[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  114.265 190.18 114.405 190.32 ;
    END
  END w_data_i[153]
  PIN w_data_i[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 64.715 146.865 64.785 ;
    END
  END w_data_i[154]
  PIN w_data_i[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  63.865 190.18 64.005 190.32 ;
    END
  END w_data_i[155]
  PIN w_data_i[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  87.945 190.18 88.085 190.32 ;
    END
  END w_data_i[156]
  PIN w_data_i[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 59.395 0.07 59.465 ;
    END
  END w_data_i[157]
  PIN w_data_i[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 144.235 0.07 144.305 ;
    END
  END w_data_i[158]
  PIN w_data_i[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.945 190.18 18.085 190.32 ;
    END
  END w_data_i[159]
  PIN w_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 153.755 146.865 153.825 ;
    END
  END w_data_i[15]
  PIN w_data_i[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 67.235 0.07 67.305 ;
    END
  END w_data_i[160]
  PIN w_data_i[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 96.635 146.865 96.705 ;
    END
  END w_data_i[161]
  PIN w_data_i[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 10.675 146.865 10.745 ;
    END
  END w_data_i[162]
  PIN w_data_i[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  62.185 190.18 62.325 190.32 ;
    END
  END w_data_i[163]
  PIN w_data_i[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  22.425 190.18 22.565 190.32 ;
    END
  END w_data_i[164]
  PIN w_data_i[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  137.225 0 137.365 0.14 ;
    END
  END w_data_i[165]
  PIN w_data_i[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  115.945 0 116.085 0.14 ;
    END
  END w_data_i[166]
  PIN w_data_i[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 183.715 0.07 183.785 ;
    END
  END w_data_i[167]
  PIN w_data_i[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 80.115 0.07 80.185 ;
    END
  END w_data_i[168]
  PIN w_data_i[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 127.715 146.865 127.785 ;
    END
  END w_data_i[169]
  PIN w_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 103.355 0.07 103.425 ;
    END
  END w_data_i[16]
  PIN w_data_i[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 120.995 146.865 121.065 ;
    END
  END w_data_i[170]
  PIN w_data_i[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 78.715 146.865 78.785 ;
    END
  END w_data_i[171]
  PIN w_data_i[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 102.235 0.07 102.305 ;
    END
  END w_data_i[172]
  PIN w_data_i[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 146.195 0.07 146.265 ;
    END
  END w_data_i[173]
  PIN w_data_i[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 58.835 146.865 58.905 ;
    END
  END w_data_i[174]
  PIN w_data_i[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 118.755 146.865 118.825 ;
    END
  END w_data_i[175]
  PIN w_data_i[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 127.995 0.07 128.065 ;
    END
  END w_data_i[176]
  PIN w_data_i[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 47.915 0.07 47.985 ;
    END
  END w_data_i[177]
  PIN w_data_i[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 75.915 146.865 75.985 ;
    END
  END w_data_i[178]
  PIN w_data_i[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 47.355 146.865 47.425 ;
    END
  END w_data_i[179]
  PIN w_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 114.835 0.07 114.905 ;
    END
  END w_data_i[17]
  PIN w_data_i[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 149.555 0.07 149.625 ;
    END
  END w_data_i[180]
  PIN w_data_i[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 108.115 146.865 108.185 ;
    END
  END w_data_i[181]
  PIN w_data_i[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  38.105 190.18 38.245 190.32 ;
    END
  END w_data_i[182]
  PIN w_data_i[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 4.515 146.865 4.585 ;
    END
  END w_data_i[183]
  PIN w_data_i[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 9.275 146.865 9.345 ;
    END
  END w_data_i[184]
  PIN w_data_i[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 1.155 0.07 1.225 ;
    END
  END w_data_i[185]
  PIN w_data_i[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 41.195 146.865 41.265 ;
    END
  END w_data_i[186]
  PIN w_data_i[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 84.875 146.865 84.945 ;
    END
  END w_data_i[187]
  PIN w_data_i[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 11.235 0.07 11.305 ;
    END
  END w_data_i[188]
  PIN w_data_i[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 148.995 0.07 149.065 ;
    END
  END w_data_i[189]
  PIN w_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  28.585 190.18 28.725 190.32 ;
    END
  END w_data_i[18]
  PIN w_data_i[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 136.675 0.07 136.745 ;
    END
  END w_data_i[190]
  PIN w_data_i[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 132.195 146.865 132.265 ;
    END
  END w_data_i[191]
  PIN w_data_i[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 152.355 146.865 152.425 ;
    END
  END w_data_i[192]
  PIN w_data_i[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  138.905 190.18 139.045 190.32 ;
    END
  END w_data_i[193]
  PIN w_data_i[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 157.395 0.07 157.465 ;
    END
  END w_data_i[194]
  PIN w_data_i[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 25.235 0.07 25.305 ;
    END
  END w_data_i[195]
  PIN w_data_i[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 42.595 146.865 42.665 ;
    END
  END w_data_i[196]
  PIN w_data_i[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 110.075 0.07 110.145 ;
    END
  END w_data_i[197]
  PIN w_data_i[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  112.025 0 112.165 0.14 ;
    END
  END w_data_i[198]
  PIN w_data_i[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 141.435 0.07 141.505 ;
    END
  END w_data_i[199]
  PIN w_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 83.475 146.865 83.545 ;
    END
  END w_data_i[19]
  PIN w_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 2.555 146.865 2.625 ;
    END
  END w_data_i[1]
  PIN w_data_i[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.665 0 10.805 0.14 ;
    END
  END w_data_i[200]
  PIN w_data_i[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 153.195 146.865 153.265 ;
    END
  END w_data_i[201]
  PIN w_data_i[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  110.905 0 111.045 0.14 ;
    END
  END w_data_i[202]
  PIN w_data_i[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  142.825 0 142.965 0.14 ;
    END
  END w_data_i[203]
  PIN w_data_i[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  35.865 190.18 36.005 190.32 ;
    END
  END w_data_i[204]
  PIN w_data_i[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 135.555 146.865 135.625 ;
    END
  END w_data_i[205]
  PIN w_data_i[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 83.195 0.07 83.265 ;
    END
  END w_data_i[206]
  PIN w_data_i[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.915 0.07 12.985 ;
    END
  END w_data_i[207]
  PIN w_data_i[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 82.915 146.865 82.985 ;
    END
  END w_data_i[208]
  PIN w_data_i[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 103.635 146.865 103.705 ;
    END
  END w_data_i[209]
  PIN w_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 25.795 146.865 25.865 ;
    END
  END w_data_i[20]
  PIN w_data_i[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 77.315 0.07 77.385 ;
    END
  END w_data_i[210]
  PIN w_data_i[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 19.075 146.865 19.145 ;
    END
  END w_data_i[211]
  PIN w_data_i[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  3.385 0 3.525 0.14 ;
    END
  END w_data_i[212]
  PIN w_data_i[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  39.785 190.18 39.925 190.32 ;
    END
  END w_data_i[213]
  PIN w_data_i[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 142.275 146.865 142.345 ;
    END
  END w_data_i[214]
  PIN w_data_i[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 186.235 0.07 186.305 ;
    END
  END w_data_i[215]
  PIN w_data_i[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 159.075 0.07 159.145 ;
    END
  END w_data_i[216]
  PIN w_data_i[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 48.755 146.865 48.825 ;
    END
  END w_data_i[217]
  PIN w_data_i[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  6.185 0 6.325 0.14 ;
    END
  END w_data_i[218]
  PIN w_data_i[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 117.075 146.865 117.145 ;
    END
  END w_data_i[219]
  PIN w_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 125.755 146.865 125.825 ;
    END
  END w_data_i[21]
  PIN w_data_i[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 146.475 146.865 146.545 ;
    END
  END w_data_i[220]
  PIN w_data_i[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 100.835 0.07 100.905 ;
    END
  END w_data_i[221]
  PIN w_data_i[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 185.115 146.865 185.185 ;
    END
  END w_data_i[222]
  PIN w_data_i[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  106.425 0 106.565 0.14 ;
    END
  END w_data_i[223]
  PIN w_data_i[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 20.475 0.07 20.545 ;
    END
  END w_data_i[224]
  PIN w_data_i[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  55.465 0 55.605 0.14 ;
    END
  END w_data_i[225]
  PIN w_data_i[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  108.105 190.18 108.245 190.32 ;
    END
  END w_data_i[226]
  PIN w_data_i[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 139.755 146.865 139.825 ;
    END
  END w_data_i[227]
  PIN w_data_i[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 83.475 0.07 83.545 ;
    END
  END w_data_i[228]
  PIN w_data_i[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 185.955 146.865 186.025 ;
    END
  END w_data_i[229]
  PIN w_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 61.915 146.865 61.985 ;
    END
  END w_data_i[22]
  PIN w_data_i[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  79.545 190.18 79.685 190.32 ;
    END
  END w_data_i[230]
  PIN w_data_i[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  99.705 190.18 99.845 190.32 ;
    END
  END w_data_i[231]
  PIN w_data_i[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  71.705 190.18 71.845 190.32 ;
    END
  END w_data_i[232]
  PIN w_data_i[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  104.745 190.18 104.885 190.32 ;
    END
  END w_data_i[233]
  PIN w_data_i[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 170.275 146.865 170.345 ;
    END
  END w_data_i[234]
  PIN w_data_i[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 161.875 146.865 161.945 ;
    END
  END w_data_i[235]
  PIN w_data_i[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 164.395 0.07 164.465 ;
    END
  END w_data_i[236]
  PIN w_data_i[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 21.315 146.865 21.385 ;
    END
  END w_data_i[237]
  PIN w_data_i[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 41.475 146.865 41.545 ;
    END
  END w_data_i[238]
  PIN w_data_i[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  126.585 0 126.725 0.14 ;
    END
  END w_data_i[239]
  PIN w_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 38.675 0.07 38.745 ;
    END
  END w_data_i[23]
  PIN w_data_i[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  73.385 190.18 73.525 190.32 ;
    END
  END w_data_i[240]
  PIN w_data_i[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  59.945 190.18 60.085 190.32 ;
    END
  END w_data_i[241]
  PIN w_data_i[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 116.795 146.865 116.865 ;
    END
  END w_data_i[242]
  PIN w_data_i[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 177.555 0.07 177.625 ;
    END
  END w_data_i[243]
  PIN w_data_i[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.025 190.18 14.165 190.32 ;
    END
  END w_data_i[244]
  PIN w_data_i[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  62.745 0 62.885 0.14 ;
    END
  END w_data_i[245]
  PIN w_data_i[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 184.835 0.07 184.905 ;
    END
  END w_data_i[246]
  PIN w_data_i[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 10.395 146.865 10.465 ;
    END
  END w_data_i[247]
  PIN w_data_i[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 16.555 146.865 16.625 ;
    END
  END w_data_i[248]
  PIN w_data_i[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 108.955 146.865 109.025 ;
    END
  END w_data_i[249]
  PIN w_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 104.755 146.865 104.825 ;
    END
  END w_data_i[24]
  PIN w_data_i[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 26.635 0.07 26.705 ;
    END
  END w_data_i[250]
  PIN w_data_i[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 186.515 0.07 186.585 ;
    END
  END w_data_i[251]
  PIN w_data_i[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  107.545 190.18 107.685 190.32 ;
    END
  END w_data_i[252]
  PIN w_data_i[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  120.985 0 121.125 0.14 ;
    END
  END w_data_i[253]
  PIN w_data_i[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 155.155 146.865 155.225 ;
    END
  END w_data_i[254]
  PIN w_data_i[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 6.475 146.865 6.545 ;
    END
  END w_data_i[255]
  PIN w_data_i[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 17.115 146.865 17.185 ;
    END
  END w_data_i[256]
  PIN w_data_i[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 168.875 146.865 168.945 ;
    END
  END w_data_i[257]
  PIN w_data_i[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 160.195 0.07 160.265 ;
    END
  END w_data_i[258]
  PIN w_data_i[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 112.595 0.07 112.665 ;
    END
  END w_data_i[259]
  PIN w_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  26.345 190.18 26.485 190.32 ;
    END
  END w_data_i[25]
  PIN w_data_i[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  145.625 0 145.765 0.14 ;
    END
  END w_data_i[260]
  PIN w_data_i[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  79.545 0 79.685 0.14 ;
    END
  END w_data_i[261]
  PIN w_data_i[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 184.555 146.865 184.625 ;
    END
  END w_data_i[262]
  PIN w_data_i[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 46.795 146.865 46.865 ;
    END
  END w_data_i[263]
  PIN w_data_i[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 164.395 146.865 164.465 ;
    END
  END w_data_i[264]
  PIN w_data_i[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  96.905 0 97.045 0.14 ;
    END
  END w_data_i[265]
  PIN w_data_i[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 28.315 0.07 28.385 ;
    END
  END w_data_i[266]
  PIN w_data_i[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 116.795 0.07 116.865 ;
    END
  END w_data_i[267]
  PIN w_data_i[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 110.075 146.865 110.145 ;
    END
  END w_data_i[268]
  PIN w_data_i[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 64.155 146.865 64.225 ;
    END
  END w_data_i[269]
  PIN w_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 68.075 146.865 68.145 ;
    END
  END w_data_i[26]
  PIN w_data_i[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 172.235 146.865 172.305 ;
    END
  END w_data_i[270]
  PIN w_data_i[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 37.835 0.07 37.905 ;
    END
  END w_data_i[271]
  PIN w_data_i[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  123.785 0 123.925 0.14 ;
    END
  END w_data_i[272]
  PIN w_data_i[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 66.675 0.07 66.745 ;
    END
  END w_data_i[273]
  PIN w_data_i[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 157.115 146.865 157.185 ;
    END
  END w_data_i[274]
  PIN w_data_i[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 51.835 146.865 51.905 ;
    END
  END w_data_i[275]
  PIN w_data_i[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 5.915 0.07 5.985 ;
    END
  END w_data_i[276]
  PIN w_data_i[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  91.865 190.18 92.005 190.32 ;
    END
  END w_data_i[277]
  PIN w_data_i[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 110.355 146.865 110.425 ;
    END
  END w_data_i[278]
  PIN w_data_i[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 102.795 0.07 102.865 ;
    END
  END w_data_i[279]
  PIN w_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  11.785 0 11.925 0.14 ;
    END
  END w_data_i[27]
  PIN w_data_i[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 7.035 146.865 7.105 ;
    END
  END w_data_i[280]
  PIN w_data_i[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 54.075 0.07 54.145 ;
    END
  END w_data_i[281]
  PIN w_data_i[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 38.395 0.07 38.465 ;
    END
  END w_data_i[282]
  PIN w_data_i[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 126.035 0.07 126.105 ;
    END
  END w_data_i[283]
  PIN w_data_i[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  50.425 190.18 50.565 190.32 ;
    END
  END w_data_i[284]
  PIN w_data_i[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 49.035 0.07 49.105 ;
    END
  END w_data_i[285]
  PIN w_data_i[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 179.235 146.865 179.305 ;
    END
  END w_data_i[286]
  PIN w_data_i[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  134.985 0 135.125 0.14 ;
    END
  END w_data_i[287]
  PIN w_data_i[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 112.035 146.865 112.105 ;
    END
  END w_data_i[288]
  PIN w_data_i[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 23.835 0.07 23.905 ;
    END
  END w_data_i[289]
  PIN w_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 147.595 0.07 147.665 ;
    END
  END w_data_i[28]
  PIN w_data_i[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  61.065 190.18 61.205 190.32 ;
    END
  END w_data_i[290]
  PIN w_data_i[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.875 0.07 7.945 ;
    END
  END w_data_i[291]
  PIN w_data_i[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  65.545 0 65.685 0.14 ;
    END
  END w_data_i[292]
  PIN w_data_i[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  72.825 190.18 72.965 190.32 ;
    END
  END w_data_i[293]
  PIN w_data_i[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 124.075 146.865 124.145 ;
    END
  END w_data_i[294]
  PIN w_data_i[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 73.955 146.865 74.025 ;
    END
  END w_data_i[295]
  PIN w_data_i[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 160.195 146.865 160.265 ;
    END
  END w_data_i[296]
  PIN w_data_i[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 162.435 0.07 162.505 ;
    END
  END w_data_i[297]
  PIN w_data_i[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 141.715 0.07 141.785 ;
    END
  END w_data_i[298]
  PIN w_data_i[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 100.835 146.865 100.905 ;
    END
  END w_data_i[299]
  PIN w_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 63.315 146.865 63.385 ;
    END
  END w_data_i[29]
  PIN w_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  75.625 190.18 75.765 190.32 ;
    END
  END w_data_i[2]
  PIN w_data_i[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 137.515 0.07 137.585 ;
    END
  END w_data_i[300]
  PIN w_data_i[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 113.435 0.07 113.505 ;
    END
  END w_data_i[301]
  PIN w_data_i[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 48.475 0.07 48.545 ;
    END
  END w_data_i[302]
  PIN w_data_i[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 82.075 0.07 82.145 ;
    END
  END w_data_i[303]
  PIN w_data_i[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  103.625 190.18 103.765 190.32 ;
    END
  END w_data_i[304]
  PIN w_data_i[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.035 0.07 7.105 ;
    END
  END w_data_i[305]
  PIN w_data_i[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 178.395 146.865 178.465 ;
    END
  END w_data_i[306]
  PIN w_data_i[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 148.995 146.865 149.065 ;
    END
  END w_data_i[307]
  PIN w_data_i[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 146.755 0.07 146.825 ;
    END
  END w_data_i[308]
  PIN w_data_i[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 134.435 146.865 134.505 ;
    END
  END w_data_i[309]
  PIN w_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 89.355 0.07 89.425 ;
    END
  END w_data_i[30]
  PIN w_data_i[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 95.515 146.865 95.585 ;
    END
  END w_data_i[310]
  PIN w_data_i[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 94.675 0.07 94.745 ;
    END
  END w_data_i[311]
  PIN w_data_i[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 51.275 0.07 51.345 ;
    END
  END w_data_i[312]
  PIN w_data_i[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  109.225 0 109.365 0.14 ;
    END
  END w_data_i[313]
  PIN w_data_i[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 184.275 146.865 184.345 ;
    END
  END w_data_i[314]
  PIN w_data_i[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 69.475 0.07 69.545 ;
    END
  END w_data_i[315]
  PIN w_data_i[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 40.635 0.07 40.705 ;
    END
  END w_data_i[316]
  PIN w_data_i[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 180.355 0.07 180.425 ;
    END
  END w_data_i[317]
  PIN w_data_i[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 58.555 146.865 58.625 ;
    END
  END w_data_i[318]
  PIN w_data_i[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 33.355 146.865 33.425 ;
    END
  END w_data_i[319]
  PIN w_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  25.225 0 25.365 0.14 ;
    END
  END w_data_i[31]
  PIN w_data_i[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  38.665 0 38.805 0.14 ;
    END
  END w_data_i[320]
  PIN w_data_i[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 84.595 146.865 84.665 ;
    END
  END w_data_i[321]
  PIN w_data_i[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 109.235 0.07 109.305 ;
    END
  END w_data_i[322]
  PIN w_data_i[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 150.955 0.07 151.025 ;
    END
  END w_data_i[323]
  PIN w_data_i[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 160.475 146.865 160.545 ;
    END
  END w_data_i[324]
  PIN w_data_i[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 91.315 0.07 91.385 ;
    END
  END w_data_i[325]
  PIN w_data_i[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  28.025 0 28.165 0.14 ;
    END
  END w_data_i[326]
  PIN w_data_i[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 140.875 0.07 140.945 ;
    END
  END w_data_i[327]
  PIN w_data_i[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 37.275 146.865 37.345 ;
    END
  END w_data_i[328]
  PIN w_data_i[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  113.705 0 113.845 0.14 ;
    END
  END w_data_i[329]
  PIN w_data_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 43.435 146.865 43.505 ;
    END
  END w_data_i[32]
  PIN w_data_i[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 133.315 0.07 133.385 ;
    END
  END w_data_i[330]
  PIN w_data_i[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 119.595 146.865 119.665 ;
    END
  END w_data_i[331]
  PIN w_data_i[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  130.505 190.18 130.645 190.32 ;
    END
  END w_data_i[332]
  PIN w_data_i[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 25.235 146.865 25.305 ;
    END
  END w_data_i[333]
  PIN w_data_i[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 2.555 0.07 2.625 ;
    END
  END w_data_i[334]
  PIN w_data_i[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 150.395 0.07 150.465 ;
    END
  END w_data_i[335]
  PIN w_data_i[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 26.075 146.865 26.145 ;
    END
  END w_data_i[336]
  PIN w_data_i[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 145.635 0.07 145.705 ;
    END
  END w_data_i[337]
  PIN w_data_i[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  50.425 0 50.565 0.14 ;
    END
  END w_data_i[338]
  PIN w_data_i[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 69.475 146.865 69.545 ;
    END
  END w_data_i[339]
  PIN w_data_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 85.435 146.865 85.505 ;
    END
  END w_data_i[33]
  PIN w_data_i[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  119.865 190.18 120.005 190.32 ;
    END
  END w_data_i[340]
  PIN w_data_i[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 18.515 0.07 18.585 ;
    END
  END w_data_i[341]
  PIN w_data_i[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 125.475 0.07 125.545 ;
    END
  END w_data_i[342]
  PIN w_data_i[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 97.195 0.07 97.265 ;
    END
  END w_data_i[343]
  PIN w_data_i[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 64.435 0.07 64.505 ;
    END
  END w_data_i[344]
  PIN w_data_i[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  132.185 0 132.325 0.14 ;
    END
  END w_data_i[345]
  PIN w_data_i[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 152.355 0.07 152.425 ;
    END
  END w_data_i[346]
  PIN w_data_i[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 105.315 0.07 105.385 ;
    END
  END w_data_i[347]
  PIN w_data_i[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 70.035 0.07 70.105 ;
    END
  END w_data_i[348]
  PIN w_data_i[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 34.475 146.865 34.545 ;
    END
  END w_data_i[349]
  PIN w_data_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 95.235 0.07 95.305 ;
    END
  END w_data_i[34]
  PIN w_data_i[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  120.985 190.18 121.125 190.32 ;
    END
  END w_data_i[350]
  PIN w_data_i[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 15.995 146.865 16.065 ;
    END
  END w_data_i[351]
  PIN w_data_i[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 120.155 146.865 120.225 ;
    END
  END w_data_i[352]
  PIN w_data_i[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 93.555 146.865 93.625 ;
    END
  END w_data_i[353]
  PIN w_data_i[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 140.315 146.865 140.385 ;
    END
  END w_data_i[354]
  PIN w_data_i[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 45.955 0.07 46.025 ;
    END
  END w_data_i[355]
  PIN w_data_i[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  131.065 0 131.205 0.14 ;
    END
  END w_data_i[356]
  PIN w_data_i[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 70.595 0.07 70.665 ;
    END
  END w_data_i[357]
  PIN w_data_i[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 110.635 0.07 110.705 ;
    END
  END w_data_i[358]
  PIN w_data_i[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 178.955 0.07 179.025 ;
    END
  END w_data_i[359]
  PIN w_data_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 68.915 146.865 68.985 ;
    END
  END w_data_i[35]
  PIN w_data_i[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 67.795 0.07 67.865 ;
    END
  END w_data_i[360]
  PIN w_data_i[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 14.315 0.07 14.385 ;
    END
  END w_data_i[361]
  PIN w_data_i[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 8.435 0.07 8.505 ;
    END
  END w_data_i[362]
  PIN w_data_i[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 189.035 146.865 189.105 ;
    END
  END w_data_i[363]
  PIN w_data_i[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 19.915 146.865 19.985 ;
    END
  END w_data_i[364]
  PIN w_data_i[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 37.835 146.865 37.905 ;
    END
  END w_data_i[365]
  PIN w_data_i[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  89.065 0 89.205 0.14 ;
    END
  END w_data_i[366]
  PIN w_data_i[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 33.915 0.07 33.985 ;
    END
  END w_data_i[367]
  PIN w_data_i[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 56.595 146.865 56.665 ;
    END
  END w_data_i[368]
  PIN w_data_i[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 72.555 146.865 72.625 ;
    END
  END w_data_i[369]
  PIN w_data_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 9.835 0.07 9.905 ;
    END
  END w_data_i[36]
  PIN w_data_i[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  99.705 0 99.845 0.14 ;
    END
  END w_data_i[370]
  PIN w_data_i[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  11.225 190.18 11.365 190.32 ;
    END
  END w_data_i[371]
  PIN w_data_i[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 59.955 146.865 60.025 ;
    END
  END w_data_i[372]
  PIN w_data_i[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 148.155 146.865 148.225 ;
    END
  END w_data_i[373]
  PIN w_data_i[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 162.995 0.07 163.065 ;
    END
  END w_data_i[374]
  PIN w_data_i[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 158.795 0.07 158.865 ;
    END
  END w_data_i[375]
  PIN w_data_i[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 98.315 146.865 98.385 ;
    END
  END w_data_i[376]
  PIN w_data_i[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 3.955 146.865 4.025 ;
    END
  END w_data_i[377]
  PIN w_data_i[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 71.995 0.07 72.065 ;
    END
  END w_data_i[378]
  PIN w_data_i[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 89.915 0.07 89.985 ;
    END
  END w_data_i[379]
  PIN w_data_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 96.075 0.07 96.145 ;
    END
  END w_data_i[37]
  PIN w_data_i[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 164.955 0.07 165.025 ;
    END
  END w_data_i[380]
  PIN w_data_i[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  86.825 0 86.965 0.14 ;
    END
  END w_data_i[381]
  PIN w_data_i[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  145.625 190.18 145.765 190.32 ;
    END
  END w_data_i[382]
  PIN w_data_i[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 49.875 146.865 49.945 ;
    END
  END w_data_i[383]
  PIN w_data_i[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 10.395 0.07 10.465 ;
    END
  END w_data_i[384]
  PIN w_data_i[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 186.515 146.865 186.585 ;
    END
  END w_data_i[385]
  PIN w_data_i[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 138.075 0.07 138.145 ;
    END
  END w_data_i[386]
  PIN w_data_i[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 158.235 0.07 158.305 ;
    END
  END w_data_i[387]
  PIN w_data_i[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  134.425 0 134.565 0.14 ;
    END
  END w_data_i[388]
  PIN w_data_i[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  90.745 190.18 90.885 190.32 ;
    END
  END w_data_i[389]
  PIN w_data_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 85.435 0.07 85.505 ;
    END
  END w_data_i[38]
  PIN w_data_i[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 60.515 0.07 60.585 ;
    END
  END w_data_i[390]
  PIN w_data_i[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.955 0.07 32.025 ;
    END
  END w_data_i[391]
  PIN w_data_i[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 129.395 0.07 129.465 ;
    END
  END w_data_i[392]
  PIN w_data_i[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 23.835 146.865 23.905 ;
    END
  END w_data_i[393]
  PIN w_data_i[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 12.635 146.865 12.705 ;
    END
  END w_data_i[394]
  PIN w_data_i[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  35.305 190.18 35.445 190.32 ;
    END
  END w_data_i[395]
  PIN w_data_i[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 154.875 146.865 154.945 ;
    END
  END w_data_i[396]
  PIN w_data_i[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 100.275 146.865 100.345 ;
    END
  END w_data_i[397]
  PIN w_data_i[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 182.315 146.865 182.385 ;
    END
  END w_data_i[398]
  PIN w_data_i[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 32.795 146.865 32.865 ;
    END
  END w_data_i[399]
  PIN w_data_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 39.795 0.07 39.865 ;
    END
  END w_data_i[39]
  PIN w_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 140.315 0.07 140.385 ;
    END
  END w_data_i[3]
  PIN w_data_i[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  80.665 190.18 80.805 190.32 ;
    END
  END w_data_i[400]
  PIN w_data_i[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 143.115 146.865 143.185 ;
    END
  END w_data_i[401]
  PIN w_data_i[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 166.915 146.865 166.985 ;
    END
  END w_data_i[402]
  PIN w_data_i[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 61.355 146.865 61.425 ;
    END
  END w_data_i[403]
  PIN w_data_i[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 129.675 146.865 129.745 ;
    END
  END w_data_i[404]
  PIN w_data_i[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  127.705 190.18 127.845 190.32 ;
    END
  END w_data_i[405]
  PIN w_data_i[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 3.115 0.07 3.185 ;
    END
  END w_data_i[406]
  PIN w_data_i[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  26.345 0 26.485 0.14 ;
    END
  END w_data_i[407]
  PIN w_data_i[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 13.755 146.865 13.825 ;
    END
  END w_data_i[408]
  PIN w_data_i[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  91.865 0 92.005 0.14 ;
    END
  END w_data_i[409]
  PIN w_data_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 43.155 0.07 43.225 ;
    END
  END w_data_i[40]
  PIN w_data_i[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  21.305 0 21.445 0.14 ;
    END
  END w_data_i[410]
  PIN w_data_i[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 36.995 0.07 37.065 ;
    END
  END w_data_i[411]
  PIN w_data_i[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 23.275 0.07 23.345 ;
    END
  END w_data_i[412]
  PIN w_data_i[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  58.265 190.18 58.405 190.32 ;
    END
  END w_data_i[413]
  PIN w_data_i[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 152.915 146.865 152.985 ;
    END
  END w_data_i[414]
  PIN w_data_i[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.745 0 34.885 0.14 ;
    END
  END w_data_i[415]
  PIN w_data_i[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 50.715 0.07 50.785 ;
    END
  END w_data_i[416]
  PIN w_data_i[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 38.115 146.865 38.185 ;
    END
  END w_data_i[417]
  PIN w_data_i[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  2.265 190.18 2.405 190.32 ;
    END
  END w_data_i[418]
  PIN w_data_i[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 29.995 146.865 30.065 ;
    END
  END w_data_i[419]
  PIN w_data_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 56.595 0.07 56.665 ;
    END
  END w_data_i[41]
  PIN w_data_i[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  42.585 190.18 42.725 190.32 ;
    END
  END w_data_i[420]
  PIN w_data_i[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  8.425 190.18 8.565 190.32 ;
    END
  END w_data_i[421]
  PIN w_data_i[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 71.435 0.07 71.505 ;
    END
  END w_data_i[422]
  PIN w_data_i[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 17.115 0.07 17.185 ;
    END
  END w_data_i[423]
  PIN w_data_i[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 100.555 0.07 100.625 ;
    END
  END w_data_i[424]
  PIN w_data_i[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  104.185 0 104.325 0.14 ;
    END
  END w_data_i[425]
  PIN w_data_i[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 94.955 146.865 95.025 ;
    END
  END w_data_i[426]
  PIN w_data_i[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 134.155 146.865 134.225 ;
    END
  END w_data_i[427]
  PIN w_data_i[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 173.635 146.865 173.705 ;
    END
  END w_data_i[428]
  PIN w_data_i[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 134.995 0.07 135.065 ;
    END
  END w_data_i[429]
  PIN w_data_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 48.475 146.865 48.545 ;
    END
  END w_data_i[42]
  PIN w_data_i[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  109.225 190.18 109.365 190.32 ;
    END
  END w_data_i[430]
  PIN w_data_i[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 187.635 146.865 187.705 ;
    END
  END w_data_i[431]
  PIN w_data_i[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 73.115 0.07 73.185 ;
    END
  END w_data_i[432]
  PIN w_data_i[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  82.345 190.18 82.485 190.32 ;
    END
  END w_data_i[433]
  PIN w_data_i[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 70.875 146.865 70.945 ;
    END
  END w_data_i[434]
  PIN w_data_i[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 40.355 0.07 40.425 ;
    END
  END w_data_i[435]
  PIN w_data_i[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 65.275 146.865 65.345 ;
    END
  END w_data_i[436]
  PIN w_data_i[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 91.595 146.865 91.665 ;
    END
  END w_data_i[437]
  PIN w_data_i[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  56.025 0 56.165 0.14 ;
    END
  END w_data_i[438]
  PIN w_data_i[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  84.025 0 84.165 0.14 ;
    END
  END w_data_i[439]
  PIN w_data_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 19.635 0.07 19.705 ;
    END
  END w_data_i[43]
  PIN w_data_i[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 127.435 146.865 127.505 ;
    END
  END w_data_i[440]
  PIN w_data_i[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  114.825 190.18 114.965 190.32 ;
    END
  END w_data_i[441]
  PIN w_data_i[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 145.355 0.07 145.425 ;
    END
  END w_data_i[442]
  PIN w_data_i[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 138.915 0.07 138.985 ;
    END
  END w_data_i[443]
  PIN w_data_i[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 115.395 0.07 115.465 ;
    END
  END w_data_i[444]
  PIN w_data_i[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 6.475 0.07 6.545 ;
    END
  END w_data_i[445]
  PIN w_data_i[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  87.385 190.18 87.525 190.32 ;
    END
  END w_data_i[446]
  PIN w_data_i[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 88.235 146.865 88.305 ;
    END
  END w_data_i[447]
  PIN w_data_i[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 108.675 0.07 108.745 ;
    END
  END w_data_i[448]
  PIN w_data_i[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  66.665 0 66.805 0.14 ;
    END
  END w_data_i[449]
  PIN w_data_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  124.905 190.18 125.045 190.32 ;
    END
  END w_data_i[44]
  PIN w_data_i[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 176.995 0.07 177.065 ;
    END
  END w_data_i[450]
  PIN w_data_i[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 168.315 0.07 168.385 ;
    END
  END w_data_i[451]
  PIN w_data_i[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  11.785 190.18 11.925 190.32 ;
    END
  END w_data_i[452]
  PIN w_data_i[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  27.465 190.18 27.605 190.32 ;
    END
  END w_data_i[453]
  PIN w_data_i[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  30.265 190.18 30.405 190.32 ;
    END
  END w_data_i[454]
  PIN w_data_i[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 17.395 146.865 17.465 ;
    END
  END w_data_i[455]
  PIN w_data_i[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 154.875 0.07 154.945 ;
    END
  END w_data_i[456]
  PIN w_data_i[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 32.515 0.07 32.585 ;
    END
  END w_data_i[457]
  PIN w_data_i[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  5.065 0 5.205 0.14 ;
    END
  END w_data_i[458]
  PIN w_data_i[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 60.795 146.865 60.865 ;
    END
  END w_data_i[459]
  PIN w_data_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 17.955 146.865 18.025 ;
    END
  END w_data_i[45]
  PIN w_data_i[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 107.555 146.865 107.625 ;
    END
  END w_data_i[460]
  PIN w_data_i[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 172.235 0.07 172.305 ;
    END
  END w_data_i[461]
  PIN w_data_i[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 120.715 146.865 120.785 ;
    END
  END w_data_i[462]
  PIN w_data_i[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 73.395 0.07 73.465 ;
    END
  END w_data_i[463]
  PIN w_data_i[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.025 0 14.165 0.14 ;
    END
  END w_data_i[464]
  PIN w_data_i[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  67.785 0 67.925 0.14 ;
    END
  END w_data_i[465]
  PIN w_data_i[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 3.675 146.865 3.745 ;
    END
  END w_data_i[466]
  PIN w_data_i[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 156.275 0.07 156.345 ;
    END
  END w_data_i[467]
  PIN w_data_i[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 63.875 146.865 63.945 ;
    END
  END w_data_i[468]
  PIN w_data_i[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  129.385 0 129.525 0.14 ;
    END
  END w_data_i[469]
  PIN w_data_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 54.635 146.865 54.705 ;
    END
  END w_data_i[46]
  PIN w_data_i[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 177.275 146.865 177.345 ;
    END
  END w_data_i[470]
  PIN w_data_i[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  110.345 190.18 110.485 190.32 ;
    END
  END w_data_i[471]
  PIN w_data_i[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 57.435 146.865 57.505 ;
    END
  END w_data_i[472]
  PIN w_data_i[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 78.155 0.07 78.225 ;
    END
  END w_data_i[473]
  PIN w_data_i[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 92.715 146.865 92.785 ;
    END
  END w_data_i[474]
  PIN w_data_i[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  126.585 190.18 126.725 190.32 ;
    END
  END w_data_i[475]
  PIN w_data_i[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 140.035 0.07 140.105 ;
    END
  END w_data_i[476]
  PIN w_data_i[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 177.835 146.865 177.905 ;
    END
  END w_data_i[477]
  PIN w_data_i[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 53.515 146.865 53.585 ;
    END
  END w_data_i[478]
  PIN w_data_i[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 176.435 0.07 176.505 ;
    END
  END w_data_i[479]
  PIN w_data_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 108.675 146.865 108.745 ;
    END
  END w_data_i[47]
  PIN w_data_i[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 130.795 0.07 130.865 ;
    END
  END w_data_i[480]
  PIN w_data_i[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 79.275 146.865 79.345 ;
    END
  END w_data_i[481]
  PIN w_data_i[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 75.355 0.07 75.425 ;
    END
  END w_data_i[482]
  PIN w_data_i[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  41.465 0 41.605 0.14 ;
    END
  END w_data_i[483]
  PIN w_data_i[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 171.115 146.865 171.185 ;
    END
  END w_data_i[484]
  PIN w_data_i[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 19.355 146.865 19.425 ;
    END
  END w_data_i[485]
  PIN w_data_i[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  134.425 190.18 134.565 190.32 ;
    END
  END w_data_i[486]
  PIN w_data_i[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  82.905 0 83.045 0.14 ;
    END
  END w_data_i[487]
  PIN w_data_i[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 80.955 146.865 81.025 ;
    END
  END w_data_i[488]
  PIN w_data_i[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 90.755 0.07 90.825 ;
    END
  END w_data_i[489]
  PIN w_data_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 181.755 0.07 181.825 ;
    END
  END w_data_i[48]
  PIN w_data_i[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  106.425 190.18 106.565 190.32 ;
    END
  END w_data_i[490]
  PIN w_data_i[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 86.835 0.07 86.905 ;
    END
  END w_data_i[491]
  PIN w_data_i[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 101.955 0.07 102.025 ;
    END
  END w_data_i[492]
  PIN w_data_i[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 114.275 146.865 114.345 ;
    END
  END w_data_i[493]
  PIN w_data_i[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 79.835 0.07 79.905 ;
    END
  END w_data_i[494]
  PIN w_data_i[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 140.875 146.865 140.945 ;
    END
  END w_data_i[495]
  PIN w_data_i[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 156.835 0.07 156.905 ;
    END
  END w_data_i[496]
  PIN w_data_i[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 124.635 0.07 124.705 ;
    END
  END w_data_i[497]
  PIN w_data_i[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 63.315 0.07 63.385 ;
    END
  END w_data_i[498]
  PIN w_data_i[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  29.145 0 29.285 0.14 ;
    END
  END w_data_i[499]
  PIN w_data_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 15.715 146.865 15.785 ;
    END
  END w_data_i[49]
  PIN w_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  128.825 190.18 128.965 190.32 ;
    END
  END w_data_i[4]
  PIN w_data_i[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 188.475 146.865 188.545 ;
    END
  END w_data_i[500]
  PIN w_data_i[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 26.355 0.07 26.425 ;
    END
  END w_data_i[501]
  PIN w_data_i[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 175.875 146.865 175.945 ;
    END
  END w_data_i[502]
  PIN w_data_i[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 131.075 146.865 131.145 ;
    END
  END w_data_i[503]
  PIN w_data_i[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 76.755 146.865 76.825 ;
    END
  END w_data_i[504]
  PIN w_data_i[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 162.155 0.07 162.225 ;
    END
  END w_data_i[505]
  PIN w_data_i[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.185 190.18 34.325 190.32 ;
    END
  END w_data_i[506]
  PIN w_data_i[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 15.155 146.865 15.225 ;
    END
  END w_data_i[507]
  PIN w_data_i[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 52.115 146.865 52.185 ;
    END
  END w_data_i[508]
  PIN w_data_i[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 115.675 146.865 115.745 ;
    END
  END w_data_i[509]
  PIN w_data_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 85.995 0.07 86.065 ;
    END
  END w_data_i[50]
  PIN w_data_i[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 11.235 146.865 11.305 ;
    END
  END w_data_i[510]
  PIN w_data_i[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  33.065 0 33.205 0.14 ;
    END
  END w_data_i[511]
  PIN w_data_i[512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 121.555 0.07 121.625 ;
    END
  END w_data_i[512]
  PIN w_data_i[513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 167.195 146.865 167.265 ;
    END
  END w_data_i[513]
  PIN w_data_i[514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  78.425 190.18 78.565 190.32 ;
    END
  END w_data_i[514]
  PIN w_data_i[515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  117.625 0 117.765 0.14 ;
    END
  END w_data_i[515]
  PIN w_data_i[516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  6.185 190.18 6.325 190.32 ;
    END
  END w_data_i[516]
  PIN w_data_i[517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 141.155 146.865 141.225 ;
    END
  END w_data_i[517]
  PIN w_data_i[518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 44.835 146.865 44.905 ;
    END
  END w_data_i[518]
  PIN w_data_i[519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  3.385 190.18 3.525 190.32 ;
    END
  END w_data_i[519]
  PIN w_data_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 40.075 146.865 40.145 ;
    END
  END w_data_i[51]
  PIN w_data_i[520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  94.665 0 94.805 0.14 ;
    END
  END w_data_i[520]
  PIN w_data_i[521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  15.705 0 15.845 0.14 ;
    END
  END w_data_i[521]
  PIN w_data_i[522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 76.195 146.865 76.265 ;
    END
  END w_data_i[522]
  PIN w_data_i[523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 116.235 146.865 116.305 ;
    END
  END w_data_i[523]
  PIN w_data_i[524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 128.275 0.07 128.345 ;
    END
  END w_data_i[524]
  PIN w_data_i[525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  118.185 190.18 118.325 190.32 ;
    END
  END w_data_i[525]
  PIN w_data_i[526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 50.435 0.07 50.505 ;
    END
  END w_data_i[526]
  PIN w_data_i[527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 61.355 0.07 61.425 ;
    END
  END w_data_i[527]
  PIN w_data_i[528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 57.995 0.07 58.065 ;
    END
  END w_data_i[528]
  PIN w_data_i[529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.905 0 13.045 0.14 ;
    END
  END w_data_i[529]
  PIN w_data_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  63.865 0 64.005 0.14 ;
    END
  END w_data_i[52]
  PIN w_data_i[530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 149.555 146.865 149.625 ;
    END
  END w_data_i[530]
  PIN w_data_i[531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 11.795 146.865 11.865 ;
    END
  END w_data_i[531]
  PIN w_data_i[532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 188.195 0.07 188.265 ;
    END
  END w_data_i[532]
  PIN w_data_i[533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  68.905 190.18 69.045 190.32 ;
    END
  END w_data_i[533]
  PIN w_data_i[534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 98.595 0.07 98.665 ;
    END
  END w_data_i[534]
  PIN w_data_i[535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  45.385 0 45.525 0.14 ;
    END
  END w_data_i[535]
  PIN w_data_i[536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 5.635 0.07 5.705 ;
    END
  END w_data_i[536]
  PIN w_data_i[537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  81.225 190.18 81.365 190.32 ;
    END
  END w_data_i[537]
  PIN w_data_i[538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 22.995 0.07 23.065 ;
    END
  END w_data_i[538]
  PIN w_data_i[539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 183.155 146.865 183.225 ;
    END
  END w_data_i[539]
  PIN w_data_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 118.195 146.865 118.265 ;
    END
  END w_data_i[53]
  PIN w_data_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 27.195 146.865 27.265 ;
    END
  END w_data_i[54]
  PIN w_data_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  52.665 190.18 52.805 190.32 ;
    END
  END w_data_i[55]
  PIN w_data_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 132.195 0.07 132.265 ;
    END
  END w_data_i[56]
  PIN w_data_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  89.625 0 89.765 0.14 ;
    END
  END w_data_i[57]
  PIN w_data_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 155.715 146.865 155.785 ;
    END
  END w_data_i[58]
  PIN w_data_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 43.995 146.865 44.065 ;
    END
  END w_data_i[59]
  PIN w_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 111.475 146.865 111.545 ;
    END
  END w_data_i[5]
  PIN w_data_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 35.875 0.07 35.945 ;
    END
  END w_data_i[60]
  PIN w_data_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 74.235 146.865 74.305 ;
    END
  END w_data_i[61]
  PIN w_data_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  46.505 0 46.645 0.14 ;
    END
  END w_data_i[62]
  PIN w_data_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  140.025 0 140.165 0.14 ;
    END
  END w_data_i[63]
  PIN w_data_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 128.835 146.865 128.905 ;
    END
  END w_data_i[64]
  PIN w_data_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  53.225 190.18 53.365 190.32 ;
    END
  END w_data_i[65]
  PIN w_data_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  140.025 190.18 140.165 190.32 ;
    END
  END w_data_i[66]
  PIN w_data_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 74.795 146.865 74.865 ;
    END
  END w_data_i[67]
  PIN w_data_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  23.545 0 23.685 0.14 ;
    END
  END w_data_i[68]
  PIN w_data_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 146.195 146.865 146.265 ;
    END
  END w_data_i[69]
  PIN w_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.305 0 7.445 0.14 ;
    END
  END w_data_i[6]
  PIN w_data_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  137.225 190.18 137.365 190.32 ;
    END
  END w_data_i[70]
  PIN w_data_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 4.515 0.07 4.585 ;
    END
  END w_data_i[71]
  PIN w_data_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 82.075 146.865 82.145 ;
    END
  END w_data_i[72]
  PIN w_data_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  42.025 190.18 42.165 190.32 ;
    END
  END w_data_i[73]
  PIN w_data_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 20.755 146.865 20.825 ;
    END
  END w_data_i[74]
  PIN w_data_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 19.075 0.07 19.145 ;
    END
  END w_data_i[75]
  PIN w_data_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 20.475 146.865 20.545 ;
    END
  END w_data_i[76]
  PIN w_data_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END w_data_i[77]
  PIN w_data_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 36.435 146.865 36.505 ;
    END
  END w_data_i[78]
  PIN w_data_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 44.555 0.07 44.625 ;
    END
  END w_data_i[79]
  PIN w_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 98.035 0.07 98.105 ;
    END
  END w_data_i[7]
  PIN w_data_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 154.315 0.07 154.385 ;
    END
  END w_data_i[80]
  PIN w_data_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 27.195 0.07 27.265 ;
    END
  END w_data_i[81]
  PIN w_data_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  58.265 0 58.405 0.14 ;
    END
  END w_data_i[82]
  PIN w_data_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  20.745 0 20.885 0.14 ;
    END
  END w_data_i[83]
  PIN w_data_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 190.18 0.725 190.32 ;
    END
  END w_data_i[84]
  PIN w_data_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 159.635 0.07 159.705 ;
    END
  END w_data_i[85]
  PIN w_data_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 1.155 146.865 1.225 ;
    END
  END w_data_i[86]
  PIN w_data_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  49.305 190.18 49.445 190.32 ;
    END
  END w_data_i[87]
  PIN w_data_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 99.995 146.865 100.065 ;
    END
  END w_data_i[88]
  PIN w_data_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 76.755 0.07 76.825 ;
    END
  END w_data_i[89]
  PIN w_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 164.955 146.865 165.025 ;
    END
  END w_data_i[8]
  PIN w_data_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  59.945 0 60.085 0.14 ;
    END
  END w_data_i[90]
  PIN w_data_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  103.625 0 103.765 0.14 ;
    END
  END w_data_i[91]
  PIN w_data_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 8.435 146.865 8.505 ;
    END
  END w_data_i[92]
  PIN w_data_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 159.075 146.865 159.145 ;
    END
  END w_data_i[93]
  PIN w_data_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 8.715 146.865 8.785 ;
    END
  END w_data_i[94]
  PIN w_data_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  48.745 190.18 48.885 190.32 ;
    END
  END w_data_i[95]
  PIN w_data_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  46.505 190.18 46.645 190.32 ;
    END
  END w_data_i[96]
  PIN w_data_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 118.195 0.07 118.265 ;
    END
  END w_data_i[97]
  PIN w_data_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 142.275 0.07 142.345 ;
    END
  END w_data_i[98]
  PIN w_data_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 23.275 146.865 23.345 ;
    END
  END w_data_i[99]
  PIN w_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 27.755 0.07 27.825 ;
    END
  END w_data_i[9]
  PIN w_reset_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 107.555 0.07 107.625 ;
    END
  END w_reset_i
  PIN w_v_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  146.795 123.515 146.865 123.585 ;
    END
  END w_v_i
  OBS
    LAYER metal1 ;
     RECT  0 -0.085 3.23 190.32 ;
     RECT  3.23 0 146.865 190.32 ;
    LAYER metal2 ;
     RECT  0 0 146.865 190.32 ;
    LAYER metal3 ;
     RECT  0 0 146.865 190.32 ;
    LAYER metal4 ;
     RECT  0 0 146.865 190.32 ;
  END
END bsg_mem_p540
END LIBRARY
