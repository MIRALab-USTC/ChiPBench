VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MACRO bsg_mem_p28
  FOREIGN bsg_mem_p28 0 0 ;
  CLASS BLOCK ;
  SIZE 33.37 BY 23.96 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 20.915 32.3 21.085 ;
        RECT  1.14 18.115 32.3 18.285 ;
        RECT  1.14 15.315 32.3 15.485 ;
        RECT  1.14 12.515 32.3 12.685 ;
        RECT  1.14 9.715 32.3 9.885 ;
        RECT  1.14 6.915 32.3 7.085 ;
        RECT  1.14 4.115 32.3 4.285 ;
        RECT  1.14 1.315 32.3 1.485 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 22.315 32.3 22.485 ;
        RECT  1.14 19.515 32.3 19.685 ;
        RECT  1.14 16.715 32.3 16.885 ;
        RECT  1.14 13.915 32.3 14.085 ;
        RECT  1.14 11.115 32.3 11.285 ;
        RECT  1.14 8.315 32.3 8.485 ;
        RECT  1.14 5.515 32.3 5.685 ;
        RECT  1.14 2.715 32.3 2.885 ;
    END
  END VDD
  PIN r_addr_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 20.755 0.07 20.825 ;
    END
  END r_addr_i
  PIN r_data_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  33.3 15.715 33.37 15.785 ;
    END
  END r_data_o[0]
  PIN r_data_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  22.985 23.82 23.125 23.96 ;
    END
  END r_data_o[10]
  PIN r_data_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  33.3 7.035 33.37 7.105 ;
    END
  END r_data_o[11]
  PIN r_data_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  33.3 21.875 33.37 21.945 ;
    END
  END r_data_o[12]
  PIN r_data_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  33.3 9.555 33.37 9.625 ;
    END
  END r_data_o[13]
  PIN r_data_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 5.635 0.07 5.705 ;
    END
  END r_data_o[14]
  PIN r_data_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.105 0 10.245 0.14 ;
    END
  END r_data_o[15]
  PIN r_data_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 4.515 0.07 4.585 ;
    END
  END r_data_o[16]
  PIN r_data_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 3.115 0.07 3.185 ;
    END
  END r_data_o[17]
  PIN r_data_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  33.3 10.675 33.37 10.745 ;
    END
  END r_data_o[18]
  PIN r_data_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  33.3 20.755 33.37 20.825 ;
    END
  END r_data_o[19]
  PIN r_data_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  2.825 0 2.965 0.14 ;
    END
  END r_data_o[1]
  PIN r_data_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 13.195 0.07 13.265 ;
    END
  END r_data_o[20]
  PIN r_data_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.865 0 8.005 0.14 ;
    END
  END r_data_o[21]
  PIN r_data_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.905 23.82 13.045 23.96 ;
    END
  END r_data_o[22]
  PIN r_data_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  33.3 4.515 33.37 4.585 ;
    END
  END r_data_o[23]
  PIN r_data_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.945 23.82 18.085 23.96 ;
    END
  END r_data_o[24]
  PIN r_data_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  33.3 14.315 33.37 14.385 ;
    END
  END r_data_o[25]
  PIN r_data_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.105 23.82 10.245 23.96 ;
    END
  END r_data_o[26]
  PIN r_data_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 14.315 0.07 14.385 ;
    END
  END r_data_o[27]
  PIN r_data_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  32.505 0 32.645 0.14 ;
    END
  END r_data_o[2]
  PIN r_data_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  30.265 0 30.405 0.14 ;
    END
  END r_data_o[3]
  PIN r_data_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 9.555 0.07 9.625 ;
    END
  END r_data_o[4]
  PIN r_data_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  33.3 16.835 33.37 16.905 ;
    END
  END r_data_o[5]
  PIN r_data_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  27.465 0 27.605 0.14 ;
    END
  END r_data_o[6]
  PIN r_data_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  20.185 23.82 20.325 23.96 ;
    END
  END r_data_o[7]
  PIN r_data_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  33.3 1.995 33.37 2.065 ;
    END
  END r_data_o[8]
  PIN r_data_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  33.3 5.635 33.37 5.705 ;
    END
  END r_data_o[9]
  PIN r_v_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  22.985 0 23.125 0.14 ;
    END
  END r_v_i
  PIN w_addr_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  33.3 8.155 33.37 8.225 ;
    END
  END w_addr_i
  PIN w_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 15.715 0.07 15.785 ;
    END
  END w_clk_i
  PIN w_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 10.675 0.07 10.745 ;
    END
  END w_data_i[0]
  PIN w_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 8.155 0.07 8.225 ;
    END
  END w_data_i[10]
  PIN w_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 19.355 0.07 19.425 ;
    END
  END w_data_i[11]
  PIN w_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.945 0 18.085 0.14 ;
    END
  END w_data_i[12]
  PIN w_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  25.225 23.82 25.365 23.96 ;
    END
  END w_data_i[13]
  PIN w_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  2.825 23.82 2.965 23.96 ;
    END
  END w_data_i[14]
  PIN w_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  33.3 19.355 33.37 19.425 ;
    END
  END w_data_i[15]
  PIN w_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  15.145 23.82 15.285 23.96 ;
    END
  END w_data_i[16]
  PIN w_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 16.835 0.07 16.905 ;
    END
  END w_data_i[17]
  PIN w_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END w_data_i[18]
  PIN w_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.875 0.07 21.945 ;
    END
  END w_data_i[19]
  PIN w_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  32.505 23.82 32.645 23.96 ;
    END
  END w_data_i[1]
  PIN w_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  15.145 0 15.285 0.14 ;
    END
  END w_data_i[20]
  PIN w_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  33.3 18.235 33.37 18.305 ;
    END
  END w_data_i[21]
  PIN w_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  33.3 3.115 33.37 3.185 ;
    END
  END w_data_i[22]
  PIN w_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.865 23.82 8.005 23.96 ;
    END
  END w_data_i[23]
  PIN w_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  33.3 11.795 33.37 11.865 ;
    END
  END w_data_i[24]
  PIN w_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  5.065 0 5.205 0.14 ;
    END
  END w_data_i[25]
  PIN w_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.905 0 13.045 0.14 ;
    END
  END w_data_i[26]
  PIN w_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.075 0.07 12.145 ;
    END
  END w_data_i[27]
  PIN w_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 1.995 0.07 2.065 ;
    END
  END w_data_i[2]
  PIN w_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  20.185 0 20.325 0.14 ;
    END
  END w_data_i[3]
  PIN w_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  30.265 23.82 30.405 23.96 ;
    END
  END w_data_i[4]
  PIN w_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  28.025 23.82 28.165 23.96 ;
    END
  END w_data_i[5]
  PIN w_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 23.82 0.725 23.96 ;
    END
  END w_data_i[6]
  PIN w_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  5.625 23.82 5.765 23.96 ;
    END
  END w_data_i[7]
  PIN w_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  25.225 0 25.365 0.14 ;
    END
  END w_data_i[8]
  PIN w_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.035 0.07 7.105 ;
    END
  END w_data_i[9]
  PIN w_reset_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 18.235 0.07 18.305 ;
    END
  END w_reset_i
  PIN w_v_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  33.3 13.195 33.37 13.265 ;
    END
  END w_v_i
  OBS
    LAYER metal1 ;
     RECT  0 -0.085 3.23 23.96 ;
     RECT  3.23 0 33.37 23.96 ;
    LAYER metal2 ;
     RECT  0 0 33.37 23.96 ;
    LAYER metal3 ;
     RECT  0 0 33.37 23.96 ;
    LAYER metal4 ;
     RECT  0 0 33.37 23.96 ;
  END
END bsg_mem_p28
END LIBRARY
