VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MACRO bsg_mem_p99
  FOREIGN bsg_mem_p99 0 0 ;
  CLASS BLOCK ;
  SIZE 69.605 BY 35.805 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 32.115 68.59 32.285 ;
        RECT  1.14 29.315 68.59 29.485 ;
        RECT  1.14 26.515 68.59 26.685 ;
        RECT  1.14 23.715 68.59 23.885 ;
        RECT  1.14 20.915 68.59 21.085 ;
        RECT  1.14 18.115 68.59 18.285 ;
        RECT  1.14 15.315 68.59 15.485 ;
        RECT  1.14 12.515 68.59 12.685 ;
        RECT  1.14 9.715 68.59 9.885 ;
        RECT  1.14 6.915 68.59 7.085 ;
        RECT  1.14 4.115 68.59 4.285 ;
        RECT  1.14 1.315 68.59 1.485 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 33.515 68.59 33.685 ;
        RECT  1.14 30.715 68.59 30.885 ;
        RECT  1.14 27.915 68.59 28.085 ;
        RECT  1.14 25.115 68.59 25.285 ;
        RECT  1.14 22.315 68.59 22.485 ;
        RECT  1.14 19.515 68.59 19.685 ;
        RECT  1.14 16.715 68.59 16.885 ;
        RECT  1.14 13.915 68.59 14.085 ;
        RECT  1.14 11.115 68.59 11.285 ;
        RECT  1.14 8.315 68.59 8.485 ;
        RECT  1.14 5.515 68.59 5.685 ;
        RECT  1.14 2.715 68.59 2.885 ;
    END
  END VDD
  PIN r_addr_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  44.825 0 44.965 0.14 ;
    END
  END r_addr_i
  PIN r_data_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 9.275 69.605 9.345 ;
    END
  END r_data_o[0]
  PIN r_data_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.035 0.07 21.105 ;
    END
  END r_data_o[10]
  PIN r_data_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 26.915 0.07 26.985 ;
    END
  END r_data_o[11]
  PIN r_data_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 34.195 69.605 34.265 ;
    END
  END r_data_o[12]
  PIN r_data_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 25.515 0.07 25.585 ;
    END
  END r_data_o[13]
  PIN r_data_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.675 0.07 31.745 ;
    END
  END r_data_o[14]
  PIN r_data_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 27.475 69.605 27.545 ;
    END
  END r_data_o[15]
  PIN r_data_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.185 35.665 34.325 35.805 ;
    END
  END r_data_o[16]
  PIN r_data_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  21.865 0 22.005 0.14 ;
    END
  END r_data_o[17]
  PIN r_data_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  38.105 0 38.245 0.14 ;
    END
  END r_data_o[18]
  PIN r_data_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 18.795 69.605 18.865 ;
    END
  END r_data_o[19]
  PIN r_data_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 5.355 69.605 5.425 ;
    END
  END r_data_o[1]
  PIN r_data_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  11.225 35.665 11.365 35.805 ;
    END
  END r_data_o[20]
  PIN r_data_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  51.545 0 51.685 0.14 ;
    END
  END r_data_o[21]
  PIN r_data_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.185 0 34.325 0.14 ;
    END
  END r_data_o[22]
  PIN r_data_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  46.505 35.665 46.645 35.805 ;
    END
  END r_data_o[23]
  PIN r_data_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 22.715 69.605 22.785 ;
    END
  END r_data_o[24]
  PIN r_data_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  56.585 0 56.725 0.14 ;
    END
  END r_data_o[25]
  PIN r_data_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 32.795 69.605 32.865 ;
    END
  END r_data_o[26]
  PIN r_data_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 30.275 69.605 30.345 ;
    END
  END r_data_o[27]
  PIN r_data_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  59.385 0 59.525 0.14 ;
    END
  END r_data_o[28]
  PIN r_data_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 20.755 69.605 20.825 ;
    END
  END r_data_o[29]
  PIN r_data_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 20.195 69.605 20.265 ;
    END
  END r_data_o[2]
  PIN r_data_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  19.625 35.665 19.765 35.805 ;
    END
  END r_data_o[30]
  PIN r_data_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 7.315 69.605 7.385 ;
    END
  END r_data_o[31]
  PIN r_data_o[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  40.905 35.665 41.045 35.805 ;
    END
  END r_data_o[32]
  PIN r_data_o[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 21.315 69.605 21.385 ;
    END
  END r_data_o[33]
  PIN r_data_o[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 30.275 0.07 30.345 ;
    END
  END r_data_o[34]
  PIN r_data_o[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  64.985 35.665 65.125 35.805 ;
    END
  END r_data_o[35]
  PIN r_data_o[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 26.915 69.605 26.985 ;
    END
  END r_data_o[36]
  PIN r_data_o[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  57.145 35.665 57.285 35.805 ;
    END
  END r_data_o[37]
  PIN r_data_o[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 13.475 69.605 13.545 ;
    END
  END r_data_o[38]
  PIN r_data_o[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  47.625 0 47.765 0.14 ;
    END
  END r_data_o[39]
  PIN r_data_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.385 0 31.525 0.14 ;
    END
  END r_data_o[3]
  PIN r_data_o[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  1.705 35.665 1.845 35.805 ;
    END
  END r_data_o[40]
  PIN r_data_o[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 1.995 69.605 2.065 ;
    END
  END r_data_o[41]
  PIN r_data_o[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  21.865 35.665 22.005 35.805 ;
    END
  END r_data_o[42]
  PIN r_data_o[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.945 35.665 18.085 35.805 ;
    END
  END r_data_o[43]
  PIN r_data_o[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.945 0 18.085 0.14 ;
    END
  END r_data_o[44]
  PIN r_data_o[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  24.665 0 24.805 0.14 ;
    END
  END r_data_o[45]
  PIN r_data_o[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.915 0.07 12.985 ;
    END
  END r_data_o[46]
  PIN r_data_o[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 33.075 0.07 33.145 ;
    END
  END r_data_o[47]
  PIN r_data_o[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 18.795 0.07 18.865 ;
    END
  END r_data_o[48]
  PIN r_data_o[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 22.995 0.07 23.065 ;
    END
  END r_data_o[49]
  PIN r_data_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 11.235 69.605 11.305 ;
    END
  END r_data_o[4]
  PIN r_data_o[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  67.785 0 67.925 0.14 ;
    END
  END r_data_o[50]
  PIN r_data_o[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 22.155 0.07 22.225 ;
    END
  END r_data_o[51]
  PIN r_data_o[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  26.345 35.665 26.485 35.805 ;
    END
  END r_data_o[52]
  PIN r_data_o[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  15.145 35.665 15.285 35.805 ;
    END
  END r_data_o[53]
  PIN r_data_o[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 28.035 69.605 28.105 ;
    END
  END r_data_o[54]
  PIN r_data_o[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 15.435 69.605 15.505 ;
    END
  END r_data_o[55]
  PIN r_data_o[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  55.465 0 55.605 0.14 ;
    END
  END r_data_o[56]
  PIN r_data_o[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 2.555 69.605 2.625 ;
    END
  END r_data_o[57]
  PIN r_data_o[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  38.105 35.665 38.245 35.805 ;
    END
  END r_data_o[58]
  PIN r_data_o[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 32.235 69.605 32.305 ;
    END
  END r_data_o[59]
  PIN r_data_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.305 35.665 7.445 35.805 ;
    END
  END r_data_o[5]
  PIN r_data_o[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  58.265 35.665 58.405 35.805 ;
    END
  END r_data_o[60]
  PIN r_data_o[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 6.195 0.07 6.265 ;
    END
  END r_data_o[61]
  PIN r_data_o[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 16.275 0.07 16.345 ;
    END
  END r_data_o[62]
  PIN r_data_o[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 30.835 69.605 30.905 ;
    END
  END r_data_o[63]
  PIN r_data_o[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  23.545 35.665 23.685 35.805 ;
    END
  END r_data_o[64]
  PIN r_data_o[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  16.825 35.665 16.965 35.805 ;
    END
  END r_data_o[65]
  PIN r_data_o[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  66.105 0 66.245 0.14 ;
    END
  END r_data_o[66]
  PIN r_data_o[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 17.675 0.07 17.745 ;
    END
  END r_data_o[67]
  PIN r_data_o[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 28.875 0.07 28.945 ;
    END
  END r_data_o[68]
  PIN r_data_o[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  20.745 35.665 20.885 35.805 ;
    END
  END r_data_o[69]
  PIN r_data_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.305 0 7.445 0.14 ;
    END
  END r_data_o[6]
  PIN r_data_o[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 9.555 0.07 9.625 ;
    END
  END r_data_o[70]
  PIN r_data_o[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 3.955 69.605 4.025 ;
    END
  END r_data_o[71]
  PIN r_data_o[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.075 0.07 12.145 ;
    END
  END r_data_o[72]
  PIN r_data_o[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 15.435 0.07 15.505 ;
    END
  END r_data_o[73]
  PIN r_data_o[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  53.225 35.665 53.365 35.805 ;
    END
  END r_data_o[74]
  PIN r_data_o[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  24.665 35.665 24.805 35.805 ;
    END
  END r_data_o[75]
  PIN r_data_o[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  67.785 35.665 67.925 35.805 ;
    END
  END r_data_o[76]
  PIN r_data_o[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  28.585 0 28.725 0.14 ;
    END
  END r_data_o[77]
  PIN r_data_o[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 15.995 69.605 16.065 ;
    END
  END r_data_o[78]
  PIN r_data_o[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  55.465 35.665 55.605 35.805 ;
    END
  END r_data_o[79]
  PIN r_data_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 25.515 69.605 25.585 ;
    END
  END r_data_o[7]
  PIN r_data_o[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 10.675 69.605 10.745 ;
    END
  END r_data_o[80]
  PIN r_data_o[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  58.265 0 58.405 0.14 ;
    END
  END r_data_o[81]
  PIN r_data_o[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  27.465 35.665 27.605 35.805 ;
    END
  END r_data_o[82]
  PIN r_data_o[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 7.875 69.605 7.945 ;
    END
  END r_data_o[83]
  PIN r_data_o[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 20.195 0.07 20.265 ;
    END
  END r_data_o[84]
  PIN r_data_o[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 4.795 0.07 4.865 ;
    END
  END r_data_o[85]
  PIN r_data_o[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  36.425 0 36.565 0.14 ;
    END
  END r_data_o[86]
  PIN r_data_o[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 22.155 69.605 22.225 ;
    END
  END r_data_o[87]
  PIN r_data_o[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 23.555 0.07 23.625 ;
    END
  END r_data_o[88]
  PIN r_data_o[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.115 0.07 31.185 ;
    END
  END r_data_o[89]
  PIN r_data_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  22.985 0 23.125 0.14 ;
    END
  END r_data_o[8]
  PIN r_data_o[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  28.585 35.665 28.725 35.805 ;
    END
  END r_data_o[90]
  PIN r_data_o[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  11.225 0 11.365 0.14 ;
    END
  END r_data_o[91]
  PIN r_data_o[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  51.545 35.665 51.685 35.805 ;
    END
  END r_data_o[92]
  PIN r_data_o[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  68.905 35.665 69.045 35.805 ;
    END
  END r_data_o[93]
  PIN r_data_o[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 12.635 69.605 12.705 ;
    END
  END r_data_o[94]
  PIN r_data_o[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  59.945 35.665 60.085 35.805 ;
    END
  END r_data_o[95]
  PIN r_data_o[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 24.395 0.07 24.465 ;
    END
  END r_data_o[96]
  PIN r_data_o[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  35.305 35.665 35.445 35.805 ;
    END
  END r_data_o[97]
  PIN r_data_o[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  52.665 0 52.805 0.14 ;
    END
  END r_data_o[98]
  PIN r_data_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 28.875 69.605 28.945 ;
    END
  END r_data_o[9]
  PIN r_v_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  50.425 35.665 50.565 35.805 ;
    END
  END r_v_i
  PIN w_addr_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 19.355 69.605 19.425 ;
    END
  END w_addr_i
  PIN w_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 10.955 0.07 11.025 ;
    END
  END w_clk_i
  PIN w_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 35.665 0.725 35.805 ;
    END
  END w_data_i[0]
  PIN w_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 26.355 0.07 26.425 ;
    END
  END w_data_i[10]
  PIN w_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 2.835 0.07 2.905 ;
    END
  END w_data_i[11]
  PIN w_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  43.705 35.665 43.845 35.805 ;
    END
  END w_data_i[12]
  PIN w_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 5.915 69.605 5.985 ;
    END
  END w_data_i[13]
  PIN w_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 1.995 0.07 2.065 ;
    END
  END w_data_i[14]
  PIN w_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  4.505 35.665 4.645 35.805 ;
    END
  END w_data_i[15]
  PIN w_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  63.305 0 63.445 0.14 ;
    END
  END w_data_i[16]
  PIN w_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  45.945 0 46.085 0.14 ;
    END
  END w_data_i[17]
  PIN w_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.905 35.665 13.045 35.805 ;
    END
  END w_data_i[18]
  PIN w_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  42.025 35.665 42.165 35.805 ;
    END
  END w_data_i[19]
  PIN w_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 5.355 0.07 5.425 ;
    END
  END w_data_i[1]
  PIN w_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  36.985 35.665 37.125 35.805 ;
    END
  END w_data_i[20]
  PIN w_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  61.065 0 61.205 0.14 ;
    END
  END w_data_i[21]
  PIN w_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  62.185 35.665 62.325 35.805 ;
    END
  END w_data_i[22]
  PIN w_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  27.465 0 27.605 0.14 ;
    END
  END w_data_i[23]
  PIN w_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  5.625 0 5.765 0.14 ;
    END
  END w_data_i[24]
  PIN w_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 28.315 0.07 28.385 ;
    END
  END w_data_i[25]
  PIN w_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 6.755 69.605 6.825 ;
    END
  END w_data_i[26]
  PIN w_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 16.835 69.605 16.905 ;
    END
  END w_data_i[27]
  PIN w_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  20.745 0 20.885 0.14 ;
    END
  END w_data_i[28]
  PIN w_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 23.555 69.605 23.625 ;
    END
  END w_data_i[29]
  PIN w_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 3.395 69.605 3.465 ;
    END
  END w_data_i[2]
  PIN w_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  3.385 35.665 3.525 35.805 ;
    END
  END w_data_i[30]
  PIN w_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.025 35.665 14.165 35.805 ;
    END
  END w_data_i[31]
  PIN w_data_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  39.225 0 39.365 0.14 ;
    END
  END w_data_i[32]
  PIN w_data_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  16.265 0 16.405 0.14 ;
    END
  END w_data_i[33]
  PIN w_data_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  2.825 0 2.965 0.14 ;
    END
  END w_data_i[34]
  PIN w_data_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  54.345 0 54.485 0.14 ;
    END
  END w_data_i[35]
  PIN w_data_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  68.905 0 69.045 0.14 ;
    END
  END w_data_i[36]
  PIN w_data_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  61.065 35.665 61.205 35.805 ;
    END
  END w_data_i[37]
  PIN w_data_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 1.435 0.07 1.505 ;
    END
  END w_data_i[38]
  PIN w_data_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 13.475 0.07 13.545 ;
    END
  END w_data_i[39]
  PIN w_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  33.065 35.665 33.205 35.805 ;
    END
  END w_data_i[3]
  PIN w_data_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 16.835 0.07 16.905 ;
    END
  END w_data_i[40]
  PIN w_data_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 18.235 0.07 18.305 ;
    END
  END w_data_i[41]
  PIN w_data_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.345 0 12.485 0.14 ;
    END
  END w_data_i[42]
  PIN w_data_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 11.515 0.07 11.585 ;
    END
  END w_data_i[43]
  PIN w_data_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  32.505 0 32.645 0.14 ;
    END
  END w_data_i[44]
  PIN w_data_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 31.395 69.605 31.465 ;
    END
  END w_data_i[45]
  PIN w_data_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  8.425 35.665 8.565 35.805 ;
    END
  END w_data_i[46]
  PIN w_data_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  39.785 35.665 39.925 35.805 ;
    END
  END w_data_i[47]
  PIN w_data_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  8.425 0 8.565 0.14 ;
    END
  END w_data_i[48]
  PIN w_data_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 12.075 69.605 12.145 ;
    END
  END w_data_i[49]
  PIN w_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 10.115 0.07 10.185 ;
    END
  END w_data_i[4]
  PIN w_data_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 4.235 0.07 4.305 ;
    END
  END w_data_i[50]
  PIN w_data_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 17.955 69.605 18.025 ;
    END
  END w_data_i[51]
  PIN w_data_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 32.235 0.07 32.305 ;
    END
  END w_data_i[52]
  PIN w_data_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 8.155 0.07 8.225 ;
    END
  END w_data_i[53]
  PIN w_data_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 29.435 69.605 29.505 ;
    END
  END w_data_i[54]
  PIN w_data_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 14.315 0.07 14.385 ;
    END
  END w_data_i[55]
  PIN w_data_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  19.065 0 19.205 0.14 ;
    END
  END w_data_i[56]
  PIN w_data_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 14.035 69.605 14.105 ;
    END
  END w_data_i[57]
  PIN w_data_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 3.395 0.07 3.465 ;
    END
  END w_data_i[58]
  PIN w_data_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 4.515 69.605 4.585 ;
    END
  END w_data_i[59]
  PIN w_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 34.475 0.07 34.545 ;
    END
  END w_data_i[5]
  PIN w_data_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  62.185 0 62.325 0.14 ;
    END
  END w_data_i[60]
  PIN w_data_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  9.545 0 9.685 0.14 ;
    END
  END w_data_i[61]
  PIN w_data_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  29.705 0 29.845 0.14 ;
    END
  END w_data_i[62]
  PIN w_data_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 10.115 69.605 10.185 ;
    END
  END w_data_i[63]
  PIN w_data_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 33.635 69.605 33.705 ;
    END
  END w_data_i[64]
  PIN w_data_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.595 0.07 7.665 ;
    END
  END w_data_i[65]
  PIN w_data_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  64.985 0 65.125 0.14 ;
    END
  END w_data_i[66]
  PIN w_data_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 14.875 0.07 14.945 ;
    END
  END w_data_i[67]
  PIN w_data_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 14.595 69.605 14.665 ;
    END
  END w_data_i[68]
  PIN w_data_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  1.705 0 1.845 0.14 ;
    END
  END w_data_i[69]
  PIN w_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 26.075 69.605 26.145 ;
    END
  END w_data_i[6]
  PIN w_data_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  66.665 35.665 66.805 35.805 ;
    END
  END w_data_i[70]
  PIN w_data_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 1.155 69.605 1.225 ;
    END
  END w_data_i[71]
  PIN w_data_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  63.865 35.665 64.005 35.805 ;
    END
  END w_data_i[72]
  PIN w_data_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  42.025 0 42.165 0.14 ;
    END
  END w_data_i[73]
  PIN w_data_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.595 0.07 21.665 ;
    END
  END w_data_i[74]
  PIN w_data_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  43.145 0 43.285 0.14 ;
    END
  END w_data_i[75]
  PIN w_data_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END w_data_i[76]
  PIN w_data_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  49.865 0 50.005 0.14 ;
    END
  END w_data_i[77]
  PIN w_data_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 24.955 0.07 25.025 ;
    END
  END w_data_i[78]
  PIN w_data_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  6.185 35.665 6.325 35.805 ;
    END
  END w_data_i[79]
  PIN w_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.385 35.665 31.525 35.805 ;
    END
  END w_data_i[7]
  PIN w_data_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 19.635 0.07 19.705 ;
    END
  END w_data_i[80]
  PIN w_data_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.025 0 14.165 0.14 ;
    END
  END w_data_i[81]
  PIN w_data_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  4.505 0 4.645 0.14 ;
    END
  END w_data_i[82]
  PIN w_data_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  44.825 35.665 44.965 35.805 ;
    END
  END w_data_i[83]
  PIN w_data_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  30.265 35.665 30.405 35.805 ;
    END
  END w_data_i[84]
  PIN w_data_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  35.305 0 35.445 0.14 ;
    END
  END w_data_i[85]
  PIN w_data_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  54.345 35.665 54.485 35.805 ;
    END
  END w_data_i[86]
  PIN w_data_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 8.715 69.605 8.785 ;
    END
  END w_data_i[87]
  PIN w_data_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 27.755 0.07 27.825 ;
    END
  END w_data_i[88]
  PIN w_data_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 24.675 69.605 24.745 ;
    END
  END w_data_i[89]
  PIN w_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  15.145 0 15.285 0.14 ;
    END
  END w_data_i[8]
  PIN w_data_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  25.785 0 25.925 0.14 ;
    END
  END w_data_i[90]
  PIN w_data_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 6.755 0.07 6.825 ;
    END
  END w_data_i[91]
  PIN w_data_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 24.115 69.605 24.185 ;
    END
  END w_data_i[92]
  PIN w_data_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  40.905 0 41.045 0.14 ;
    END
  END w_data_i[93]
  PIN w_data_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  48.745 35.665 48.885 35.805 ;
    END
  END w_data_i[94]
  PIN w_data_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  47.625 35.665 47.765 35.805 ;
    END
  END w_data_i[95]
  PIN w_data_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 33.635 0.07 33.705 ;
    END
  END w_data_i[96]
  PIN w_data_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.105 35.665 10.245 35.805 ;
    END
  END w_data_i[97]
  PIN w_data_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  48.745 0 48.885 0.14 ;
    END
  END w_data_i[98]
  PIN w_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 8.715 0.07 8.785 ;
    END
  END w_data_i[9]
  PIN w_reset_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 29.715 0.07 29.785 ;
    END
  END w_reset_i
  PIN w_v_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  69.535 17.395 69.605 17.465 ;
    END
  END w_v_i
  OBS
    LAYER metal1 ;
     RECT  0 -0.085 3.23 35.805 ;
     RECT  3.23 0 69.605 35.805 ;
    LAYER metal2 ;
     RECT  0 0 69.605 35.805 ;
    LAYER metal3 ;
     RECT  0 0 69.605 35.805 ;
    LAYER metal4 ;
     RECT  0 0 69.605 35.805 ;
  END
END bsg_mem_p99
END LIBRARY
