VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MACRO bsg_mem_p567
  FOREIGN bsg_mem_p567 0 0 ;
  CLASS BLOCK ;
  SIZE 94.11 BY 140.16 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 138.515 93.1 138.685 ;
        RECT  1.14 135.715 93.1 135.885 ;
        RECT  1.14 132.915 93.1 133.085 ;
        RECT  1.14 130.115 93.1 130.285 ;
        RECT  1.14 127.315 93.1 127.485 ;
        RECT  1.14 124.515 93.1 124.685 ;
        RECT  1.14 121.715 93.1 121.885 ;
        RECT  1.14 118.915 93.1 119.085 ;
        RECT  1.14 116.115 93.1 116.285 ;
        RECT  1.14 113.315 93.1 113.485 ;
        RECT  1.14 110.515 93.1 110.685 ;
        RECT  1.14 107.715 93.1 107.885 ;
        RECT  1.14 104.915 93.1 105.085 ;
        RECT  1.14 102.115 93.1 102.285 ;
        RECT  1.14 99.315 93.1 99.485 ;
        RECT  1.14 96.515 93.1 96.685 ;
        RECT  1.14 93.715 93.1 93.885 ;
        RECT  1.14 90.915 93.1 91.085 ;
        RECT  1.14 88.115 93.1 88.285 ;
        RECT  1.14 85.315 93.1 85.485 ;
        RECT  1.14 82.515 93.1 82.685 ;
        RECT  1.14 79.715 93.1 79.885 ;
        RECT  1.14 76.915 93.1 77.085 ;
        RECT  1.14 74.115 93.1 74.285 ;
        RECT  1.14 71.315 93.1 71.485 ;
        RECT  1.14 68.515 93.1 68.685 ;
        RECT  1.14 65.715 93.1 65.885 ;
        RECT  1.14 62.915 93.1 63.085 ;
        RECT  1.14 60.115 93.1 60.285 ;
        RECT  1.14 57.315 93.1 57.485 ;
        RECT  1.14 54.515 93.1 54.685 ;
        RECT  1.14 51.715 93.1 51.885 ;
        RECT  1.14 48.915 93.1 49.085 ;
        RECT  1.14 46.115 93.1 46.285 ;
        RECT  1.14 43.315 93.1 43.485 ;
        RECT  1.14 40.515 93.1 40.685 ;
        RECT  1.14 37.715 93.1 37.885 ;
        RECT  1.14 34.915 93.1 35.085 ;
        RECT  1.14 32.115 93.1 32.285 ;
        RECT  1.14 29.315 93.1 29.485 ;
        RECT  1.14 26.515 93.1 26.685 ;
        RECT  1.14 23.715 93.1 23.885 ;
        RECT  1.14 20.915 93.1 21.085 ;
        RECT  1.14 18.115 93.1 18.285 ;
        RECT  1.14 15.315 93.1 15.485 ;
        RECT  1.14 12.515 93.1 12.685 ;
        RECT  1.14 9.715 93.1 9.885 ;
        RECT  1.14 6.915 93.1 7.085 ;
        RECT  1.14 4.115 93.1 4.285 ;
        RECT  1.14 1.315 93.1 1.485 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 137.115 93.1 137.285 ;
        RECT  1.14 134.315 93.1 134.485 ;
        RECT  1.14 131.515 93.1 131.685 ;
        RECT  1.14 128.715 93.1 128.885 ;
        RECT  1.14 125.915 93.1 126.085 ;
        RECT  1.14 123.115 93.1 123.285 ;
        RECT  1.14 120.315 93.1 120.485 ;
        RECT  1.14 117.515 93.1 117.685 ;
        RECT  1.14 114.715 93.1 114.885 ;
        RECT  1.14 111.915 93.1 112.085 ;
        RECT  1.14 109.115 93.1 109.285 ;
        RECT  1.14 106.315 93.1 106.485 ;
        RECT  1.14 103.515 93.1 103.685 ;
        RECT  1.14 100.715 93.1 100.885 ;
        RECT  1.14 97.915 93.1 98.085 ;
        RECT  1.14 95.115 93.1 95.285 ;
        RECT  1.14 92.315 93.1 92.485 ;
        RECT  1.14 89.515 93.1 89.685 ;
        RECT  1.14 86.715 93.1 86.885 ;
        RECT  1.14 83.915 93.1 84.085 ;
        RECT  1.14 81.115 93.1 81.285 ;
        RECT  1.14 78.315 93.1 78.485 ;
        RECT  1.14 75.515 93.1 75.685 ;
        RECT  1.14 72.715 93.1 72.885 ;
        RECT  1.14 69.915 93.1 70.085 ;
        RECT  1.14 67.115 93.1 67.285 ;
        RECT  1.14 64.315 93.1 64.485 ;
        RECT  1.14 61.515 93.1 61.685 ;
        RECT  1.14 58.715 93.1 58.885 ;
        RECT  1.14 55.915 93.1 56.085 ;
        RECT  1.14 53.115 93.1 53.285 ;
        RECT  1.14 50.315 93.1 50.485 ;
        RECT  1.14 47.515 93.1 47.685 ;
        RECT  1.14 44.715 93.1 44.885 ;
        RECT  1.14 41.915 93.1 42.085 ;
        RECT  1.14 39.115 93.1 39.285 ;
        RECT  1.14 36.315 93.1 36.485 ;
        RECT  1.14 33.515 93.1 33.685 ;
        RECT  1.14 30.715 93.1 30.885 ;
        RECT  1.14 27.915 93.1 28.085 ;
        RECT  1.14 25.115 93.1 25.285 ;
        RECT  1.14 22.315 93.1 22.485 ;
        RECT  1.14 19.515 93.1 19.685 ;
        RECT  1.14 16.715 93.1 16.885 ;
        RECT  1.14 13.915 93.1 14.085 ;
        RECT  1.14 11.115 93.1 11.285 ;
        RECT  1.14 8.315 93.1 8.485 ;
        RECT  1.14 5.515 93.1 5.685 ;
        RECT  1.14 2.715 93.1 2.885 ;
    END
  END VDD
  PIN r_addr_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 36.155 94.11 36.225 ;
    END
  END r_addr_i
  PIN r_data_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 51.275 94.11 51.345 ;
    END
  END r_data_o[0]
  PIN r_data_o[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 23.275 0.07 23.345 ;
    END
  END r_data_o[100]
  PIN r_data_o[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 80.955 94.11 81.025 ;
    END
  END r_data_o[101]
  PIN r_data_o[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 56.875 94.11 56.945 ;
    END
  END r_data_o[102]
  PIN r_data_o[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 86.555 0.07 86.625 ;
    END
  END r_data_o[103]
  PIN r_data_o[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  70.585 140.02 70.725 140.16 ;
    END
  END r_data_o[104]
  PIN r_data_o[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 94.955 0.07 95.025 ;
    END
  END r_data_o[105]
  PIN r_data_o[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 132.755 94.11 132.825 ;
    END
  END r_data_o[106]
  PIN r_data_o[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 31.955 94.11 32.025 ;
    END
  END r_data_o[107]
  PIN r_data_o[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 66.675 94.11 66.745 ;
    END
  END r_data_o[108]
  PIN r_data_o[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 17.675 0.07 17.745 ;
    END
  END r_data_o[109]
  PIN r_data_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 32.235 0.07 32.305 ;
    END
  END r_data_o[10]
  PIN r_data_o[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.875 0.07 21.945 ;
    END
  END r_data_o[110]
  PIN r_data_o[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  57.705 140.02 57.845 140.16 ;
    END
  END r_data_o[111]
  PIN r_data_o[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  35.865 140.02 36.005 140.16 ;
    END
  END r_data_o[112]
  PIN r_data_o[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 119.595 0.07 119.665 ;
    END
  END r_data_o[113]
  PIN r_data_o[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 5.635 0.07 5.705 ;
    END
  END r_data_o[114]
  PIN r_data_o[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 64.995 94.11 65.065 ;
    END
  END r_data_o[115]
  PIN r_data_o[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 75.075 94.11 75.145 ;
    END
  END r_data_o[116]
  PIN r_data_o[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 69.475 0.07 69.545 ;
    END
  END r_data_o[117]
  PIN r_data_o[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  35.305 0 35.445 0.14 ;
    END
  END r_data_o[118]
  PIN r_data_o[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 88.235 94.11 88.305 ;
    END
  END r_data_o[119]
  PIN r_data_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 84.875 94.11 84.945 ;
    END
  END r_data_o[11]
  PIN r_data_o[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  40.905 140.02 41.045 140.16 ;
    END
  END r_data_o[120]
  PIN r_data_o[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 82.635 0.07 82.705 ;
    END
  END r_data_o[121]
  PIN r_data_o[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  39.785 140.02 39.925 140.16 ;
    END
  END r_data_o[122]
  PIN r_data_o[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  50.425 140.02 50.565 140.16 ;
    END
  END r_data_o[123]
  PIN r_data_o[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 11.795 94.11 11.865 ;
    END
  END r_data_o[124]
  PIN r_data_o[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 75.355 0.07 75.425 ;
    END
  END r_data_o[125]
  PIN r_data_o[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  15.705 0 15.845 0.14 ;
    END
  END r_data_o[126]
  PIN r_data_o[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 56.035 0.07 56.105 ;
    END
  END r_data_o[127]
  PIN r_data_o[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 128.835 94.11 128.905 ;
    END
  END r_data_o[128]
  PIN r_data_o[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 123.795 94.11 123.865 ;
    END
  END r_data_o[129]
  PIN r_data_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 88.795 0.07 88.865 ;
    END
  END r_data_o[12]
  PIN r_data_o[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 40.915 94.11 40.985 ;
    END
  END r_data_o[130]
  PIN r_data_o[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 99.995 94.11 100.065 ;
    END
  END r_data_o[131]
  PIN r_data_o[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 127.715 94.11 127.785 ;
    END
  END r_data_o[132]
  PIN r_data_o[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  46.505 0 46.645 0.14 ;
    END
  END r_data_o[133]
  PIN r_data_o[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 98.035 0.07 98.105 ;
    END
  END r_data_o[134]
  PIN r_data_o[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 66.395 94.11 66.465 ;
    END
  END r_data_o[135]
  PIN r_data_o[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 38.395 0.07 38.465 ;
    END
  END r_data_o[136]
  PIN r_data_o[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 32.515 94.11 32.585 ;
    END
  END r_data_o[137]
  PIN r_data_o[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 133.875 0.07 133.945 ;
    END
  END r_data_o[138]
  PIN r_data_o[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 73.395 0.07 73.465 ;
    END
  END r_data_o[139]
  PIN r_data_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  21.305 140.02 21.445 140.16 ;
    END
  END r_data_o[13]
  PIN r_data_o[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 22.435 94.11 22.505 ;
    END
  END r_data_o[140]
  PIN r_data_o[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 115.395 0.07 115.465 ;
    END
  END r_data_o[141]
  PIN r_data_o[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 28.595 0.07 28.665 ;
    END
  END r_data_o[142]
  PIN r_data_o[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 53.515 94.11 53.585 ;
    END
  END r_data_o[143]
  PIN r_data_o[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 132.195 0.07 132.265 ;
    END
  END r_data_o[144]
  PIN r_data_o[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 53.235 0.07 53.305 ;
    END
  END r_data_o[145]
  PIN r_data_o[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  61.625 140.02 61.765 140.16 ;
    END
  END r_data_o[146]
  PIN r_data_o[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  8.985 140.02 9.125 140.16 ;
    END
  END r_data_o[147]
  PIN r_data_o[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 32.515 0.07 32.585 ;
    END
  END r_data_o[148]
  PIN r_data_o[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 4.515 0.07 4.585 ;
    END
  END r_data_o[149]
  PIN r_data_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 73.675 94.11 73.745 ;
    END
  END r_data_o[14]
  PIN r_data_o[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  84.585 0 84.725 0.14 ;
    END
  END r_data_o[150]
  PIN r_data_o[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  66.105 140.02 66.245 140.16 ;
    END
  END r_data_o[151]
  PIN r_data_o[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  43.705 0 43.845 0.14 ;
    END
  END r_data_o[152]
  PIN r_data_o[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 57.155 94.11 57.225 ;
    END
  END r_data_o[153]
  PIN r_data_o[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 59.395 94.11 59.465 ;
    END
  END r_data_o[154]
  PIN r_data_o[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 26.635 94.11 26.705 ;
    END
  END r_data_o[155]
  PIN r_data_o[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 77.595 0.07 77.665 ;
    END
  END r_data_o[156]
  PIN r_data_o[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 116.795 94.11 116.865 ;
    END
  END r_data_o[157]
  PIN r_data_o[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 7.595 94.11 7.665 ;
    END
  END r_data_o[158]
  PIN r_data_o[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 96.355 94.11 96.425 ;
    END
  END r_data_o[159]
  PIN r_data_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 29.715 94.11 29.785 ;
    END
  END r_data_o[15]
  PIN r_data_o[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  59.945 0 60.085 0.14 ;
    END
  END r_data_o[160]
  PIN r_data_o[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 102.795 0.07 102.865 ;
    END
  END r_data_o[161]
  PIN r_data_o[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  79.545 0 79.685 0.14 ;
    END
  END r_data_o[162]
  PIN r_data_o[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 121.555 0.07 121.625 ;
    END
  END r_data_o[163]
  PIN r_data_o[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 113.155 94.11 113.225 ;
    END
  END r_data_o[164]
  PIN r_data_o[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 125.755 94.11 125.825 ;
    END
  END r_data_o[165]
  PIN r_data_o[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  44.265 0 44.405 0.14 ;
    END
  END r_data_o[166]
  PIN r_data_o[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 109.515 94.11 109.585 ;
    END
  END r_data_o[167]
  PIN r_data_o[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.635 0.07 12.705 ;
    END
  END r_data_o[168]
  PIN r_data_o[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  78.425 140.02 78.565 140.16 ;
    END
  END r_data_o[169]
  PIN r_data_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  58.265 0 58.405 0.14 ;
    END
  END r_data_o[16]
  PIN r_data_o[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 43.435 94.11 43.505 ;
    END
  END r_data_o[170]
  PIN r_data_o[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 39.795 0.07 39.865 ;
    END
  END r_data_o[171]
  PIN r_data_o[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 16.835 94.11 16.905 ;
    END
  END r_data_o[172]
  PIN r_data_o[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 97.755 94.11 97.825 ;
    END
  END r_data_o[173]
  PIN r_data_o[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 114.275 94.11 114.345 ;
    END
  END r_data_o[174]
  PIN r_data_o[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  1.145 0 1.285 0.14 ;
    END
  END r_data_o[175]
  PIN r_data_o[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 52.675 0.07 52.745 ;
    END
  END r_data_o[176]
  PIN r_data_o[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 59.115 94.11 59.185 ;
    END
  END r_data_o[177]
  PIN r_data_o[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 28.315 0.07 28.385 ;
    END
  END r_data_o[178]
  PIN r_data_o[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 137.795 0.07 137.865 ;
    END
  END r_data_o[179]
  PIN r_data_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  87.945 0 88.085 0.14 ;
    END
  END r_data_o[17]
  PIN r_data_o[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  72.265 0 72.405 0.14 ;
    END
  END r_data_o[180]
  PIN r_data_o[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  50.425 0 50.565 0.14 ;
    END
  END r_data_o[181]
  PIN r_data_o[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  52.105 140.02 52.245 140.16 ;
    END
  END r_data_o[182]
  PIN r_data_o[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 111.755 0.07 111.825 ;
    END
  END r_data_o[183]
  PIN r_data_o[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 127.435 0.07 127.505 ;
    END
  END r_data_o[184]
  PIN r_data_o[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 54.635 0.07 54.705 ;
    END
  END r_data_o[185]
  PIN r_data_o[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  82.905 140.02 83.045 140.16 ;
    END
  END r_data_o[186]
  PIN r_data_o[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 126.595 0.07 126.665 ;
    END
  END r_data_o[187]
  PIN r_data_o[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 45.115 0.07 45.185 ;
    END
  END r_data_o[188]
  PIN r_data_o[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 55.195 0.07 55.265 ;
    END
  END r_data_o[189]
  PIN r_data_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  88.505 0 88.645 0.14 ;
    END
  END r_data_o[18]
  PIN r_data_o[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 99.155 94.11 99.225 ;
    END
  END r_data_o[190]
  PIN r_data_o[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 33.635 0.07 33.705 ;
    END
  END r_data_o[191]
  PIN r_data_o[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 79.835 0.07 79.905 ;
    END
  END r_data_o[192]
  PIN r_data_o[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 96.915 0.07 96.985 ;
    END
  END r_data_o[193]
  PIN r_data_o[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 34.475 94.11 34.545 ;
    END
  END r_data_o[194]
  PIN r_data_o[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 123.235 0.07 123.305 ;
    END
  END r_data_o[195]
  PIN r_data_o[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 44.835 94.11 44.905 ;
    END
  END r_data_o[196]
  PIN r_data_o[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 77.315 94.11 77.385 ;
    END
  END r_data_o[197]
  PIN r_data_o[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 45.955 94.11 46.025 ;
    END
  END r_data_o[198]
  PIN r_data_o[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  11.785 0 11.925 0.14 ;
    END
  END r_data_o[199]
  PIN r_data_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 47.915 0.07 47.985 ;
    END
  END r_data_o[19]
  PIN r_data_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 76.755 0.07 76.825 ;
    END
  END r_data_o[1]
  PIN r_data_o[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 62.755 94.11 62.825 ;
    END
  END r_data_o[200]
  PIN r_data_o[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 9.835 94.11 9.905 ;
    END
  END r_data_o[201]
  PIN r_data_o[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 118.195 0.07 118.265 ;
    END
  END r_data_o[202]
  PIN r_data_o[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 56.875 0.07 56.945 ;
    END
  END r_data_o[203]
  PIN r_data_o[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.945 0 32.085 0.14 ;
    END
  END r_data_o[204]
  PIN r_data_o[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 38.675 94.11 38.745 ;
    END
  END r_data_o[205]
  PIN r_data_o[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 114.835 0.07 114.905 ;
    END
  END r_data_o[206]
  PIN r_data_o[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 113.995 94.11 114.065 ;
    END
  END r_data_o[207]
  PIN r_data_o[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 10.115 0.07 10.185 ;
    END
  END r_data_o[208]
  PIN r_data_o[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 15.155 0.07 15.225 ;
    END
  END r_data_o[209]
  PIN r_data_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 121.275 0.07 121.345 ;
    END
  END r_data_o[20]
  PIN r_data_o[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 131.355 94.11 131.425 ;
    END
  END r_data_o[210]
  PIN r_data_o[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 129.395 0.07 129.465 ;
    END
  END r_data_o[211]
  PIN r_data_o[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 108.115 94.11 108.185 ;
    END
  END r_data_o[212]
  PIN r_data_o[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 89.915 94.11 89.985 ;
    END
  END r_data_o[213]
  PIN r_data_o[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 122.115 0.07 122.185 ;
    END
  END r_data_o[214]
  PIN r_data_o[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 36.435 0.07 36.505 ;
    END
  END r_data_o[215]
  PIN r_data_o[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 64.435 94.11 64.505 ;
    END
  END r_data_o[216]
  PIN r_data_o[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 101.115 94.11 101.185 ;
    END
  END r_data_o[217]
  PIN r_data_o[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  52.105 0 52.245 0.14 ;
    END
  END r_data_o[218]
  PIN r_data_o[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 81.795 94.11 81.865 ;
    END
  END r_data_o[219]
  PIN r_data_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 110.915 0.07 110.985 ;
    END
  END r_data_o[21]
  PIN r_data_o[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  27.465 0 27.605 0.14 ;
    END
  END r_data_o[220]
  PIN r_data_o[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 20.475 0.07 20.545 ;
    END
  END r_data_o[221]
  PIN r_data_o[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 98.875 0.07 98.945 ;
    END
  END r_data_o[222]
  PIN r_data_o[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  2.825 0 2.965 0.14 ;
    END
  END r_data_o[223]
  PIN r_data_o[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 5.355 94.11 5.425 ;
    END
  END r_data_o[224]
  PIN r_data_o[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 140.02 0.725 140.16 ;
    END
  END r_data_o[225]
  PIN r_data_o[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  92.985 0 93.125 0.14 ;
    END
  END r_data_o[226]
  PIN r_data_o[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 137.515 0.07 137.585 ;
    END
  END r_data_o[227]
  PIN r_data_o[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  91.305 0 91.445 0.14 ;
    END
  END r_data_o[228]
  PIN r_data_o[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  64.425 140.02 64.565 140.16 ;
    END
  END r_data_o[229]
  PIN r_data_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 92.995 94.11 93.065 ;
    END
  END r_data_o[22]
  PIN r_data_o[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  25.785 0 25.925 0.14 ;
    END
  END r_data_o[230]
  PIN r_data_o[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 26.355 0.07 26.425 ;
    END
  END r_data_o[231]
  PIN r_data_o[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  22.425 0 22.565 0.14 ;
    END
  END r_data_o[232]
  PIN r_data_o[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.305 140.02 7.445 140.16 ;
    END
  END r_data_o[233]
  PIN r_data_o[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 45.115 94.11 45.185 ;
    END
  END r_data_o[234]
  PIN r_data_o[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 94.955 94.11 95.025 ;
    END
  END r_data_o[235]
  PIN r_data_o[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 74.235 0.07 74.305 ;
    END
  END r_data_o[236]
  PIN r_data_o[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 54.355 94.11 54.425 ;
    END
  END r_data_o[237]
  PIN r_data_o[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 54.075 0.07 54.145 ;
    END
  END r_data_o[238]
  PIN r_data_o[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 136.675 94.11 136.745 ;
    END
  END r_data_o[239]
  PIN r_data_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  20.745 140.02 20.885 140.16 ;
    END
  END r_data_o[23]
  PIN r_data_o[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  63.305 0 63.445 0.14 ;
    END
  END r_data_o[240]
  PIN r_data_o[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 47.635 94.11 47.705 ;
    END
  END r_data_o[241]
  PIN r_data_o[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  47.065 0 47.205 0.14 ;
    END
  END r_data_o[242]
  PIN r_data_o[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.875 0.07 7.945 ;
    END
  END r_data_o[243]
  PIN r_data_o[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 0.875 94.11 0.945 ;
    END
  END r_data_o[244]
  PIN r_data_o[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  6.185 0 6.325 0.14 ;
    END
  END r_data_o[245]
  PIN r_data_o[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 56.315 0.07 56.385 ;
    END
  END r_data_o[246]
  PIN r_data_o[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  84.585 140.02 84.725 140.16 ;
    END
  END r_data_o[247]
  PIN r_data_o[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 16.555 0.07 16.625 ;
    END
  END r_data_o[248]
  PIN r_data_o[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 49.035 0.07 49.105 ;
    END
  END r_data_o[249]
  PIN r_data_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 83.195 94.11 83.265 ;
    END
  END r_data_o[24]
  PIN r_data_o[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 87.675 0.07 87.745 ;
    END
  END r_data_o[250]
  PIN r_data_o[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 14.595 0.07 14.665 ;
    END
  END r_data_o[251]
  PIN r_data_o[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 30.275 0.07 30.345 ;
    END
  END r_data_o[252]
  PIN r_data_o[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  4.505 140.02 4.645 140.16 ;
    END
  END r_data_o[253]
  PIN r_data_o[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 70.315 0.07 70.385 ;
    END
  END r_data_o[254]
  PIN r_data_o[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 67.235 94.11 67.305 ;
    END
  END r_data_o[255]
  PIN r_data_o[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 10.675 94.11 10.745 ;
    END
  END r_data_o[256]
  PIN r_data_o[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 85.155 94.11 85.225 ;
    END
  END r_data_o[257]
  PIN r_data_o[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.185 0 34.325 0.14 ;
    END
  END r_data_o[258]
  PIN r_data_o[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  80.105 0 80.245 0.14 ;
    END
  END r_data_o[259]
  PIN r_data_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 70.595 94.11 70.665 ;
    END
  END r_data_o[25]
  PIN r_data_o[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 28.595 94.11 28.665 ;
    END
  END r_data_o[260]
  PIN r_data_o[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 94.115 94.11 94.185 ;
    END
  END r_data_o[261]
  PIN r_data_o[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  13.465 140.02 13.605 140.16 ;
    END
  END r_data_o[262]
  PIN r_data_o[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  30.265 140.02 30.405 140.16 ;
    END
  END r_data_o[263]
  PIN r_data_o[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 136.395 0.07 136.465 ;
    END
  END r_data_o[264]
  PIN r_data_o[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 61.915 0.07 61.985 ;
    END
  END r_data_o[265]
  PIN r_data_o[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.945 140.02 32.085 140.16 ;
    END
  END r_data_o[266]
  PIN r_data_o[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  30.825 0 30.965 0.14 ;
    END
  END r_data_o[267]
  PIN r_data_o[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 121.555 94.11 121.625 ;
    END
  END r_data_o[268]
  PIN r_data_o[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  15.145 140.02 15.285 140.16 ;
    END
  END r_data_o[269]
  PIN r_data_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 37.835 0.07 37.905 ;
    END
  END r_data_o[26]
  PIN r_data_o[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  73.385 140.02 73.525 140.16 ;
    END
  END r_data_o[270]
  PIN r_data_o[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 65.275 0.07 65.345 ;
    END
  END r_data_o[271]
  PIN r_data_o[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 116.515 0.07 116.585 ;
    END
  END r_data_o[272]
  PIN r_data_o[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  47.065 140.02 47.205 140.16 ;
    END
  END r_data_o[273]
  PIN r_data_o[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 131.635 0.07 131.705 ;
    END
  END r_data_o[274]
  PIN r_data_o[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 105.315 0.07 105.385 ;
    END
  END r_data_o[275]
  PIN r_data_o[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 79.275 0.07 79.345 ;
    END
  END r_data_o[276]
  PIN r_data_o[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 32.795 0.07 32.865 ;
    END
  END r_data_o[277]
  PIN r_data_o[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 73.115 94.11 73.185 ;
    END
  END r_data_o[278]
  PIN r_data_o[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 105.035 0.07 105.105 ;
    END
  END r_data_o[279]
  PIN r_data_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.105 140.02 10.245 140.16 ;
    END
  END r_data_o[27]
  PIN r_data_o[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 17.115 94.11 17.185 ;
    END
  END r_data_o[280]
  PIN r_data_o[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  75.625 140.02 75.765 140.16 ;
    END
  END r_data_o[281]
  PIN r_data_o[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 70.875 94.11 70.945 ;
    END
  END r_data_o[282]
  PIN r_data_o[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  70.585 0 70.725 0.14 ;
    END
  END r_data_o[283]
  PIN r_data_o[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 117.075 0.07 117.145 ;
    END
  END r_data_o[284]
  PIN r_data_o[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 30.835 0.07 30.905 ;
    END
  END r_data_o[285]
  PIN r_data_o[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 35.315 94.11 35.385 ;
    END
  END r_data_o[286]
  PIN r_data_o[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 46.235 94.11 46.305 ;
    END
  END r_data_o[287]
  PIN r_data_o[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 119.875 0.07 119.945 ;
    END
  END r_data_o[288]
  PIN r_data_o[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  54.905 0 55.045 0.14 ;
    END
  END r_data_o[289]
  PIN r_data_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 89.635 0.07 89.705 ;
    END
  END r_data_o[28]
  PIN r_data_o[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 1.715 0.07 1.785 ;
    END
  END r_data_o[290]
  PIN r_data_o[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 6.195 0.07 6.265 ;
    END
  END r_data_o[291]
  PIN r_data_o[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 34.195 94.11 34.265 ;
    END
  END r_data_o[292]
  PIN r_data_o[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 138.635 0.07 138.705 ;
    END
  END r_data_o[293]
  PIN r_data_o[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 136.955 94.11 137.025 ;
    END
  END r_data_o[294]
  PIN r_data_o[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 123.515 94.11 123.585 ;
    END
  END r_data_o[295]
  PIN r_data_o[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 55.755 94.11 55.825 ;
    END
  END r_data_o[296]
  PIN r_data_o[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  72.265 140.02 72.405 140.16 ;
    END
  END r_data_o[297]
  PIN r_data_o[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 100.555 0.07 100.625 ;
    END
  END r_data_o[298]
  PIN r_data_o[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 61.075 94.11 61.145 ;
    END
  END r_data_o[299]
  PIN r_data_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 7.875 94.11 7.945 ;
    END
  END r_data_o[29]
  PIN r_data_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  2.265 140.02 2.405 140.16 ;
    END
  END r_data_o[2]
  PIN r_data_o[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 24.115 0.07 24.185 ;
    END
  END r_data_o[300]
  PIN r_data_o[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 94.395 94.11 94.465 ;
    END
  END r_data_o[301]
  PIN r_data_o[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 81.235 0.07 81.305 ;
    END
  END r_data_o[302]
  PIN r_data_o[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  1.705 0 1.845 0.14 ;
    END
  END r_data_o[303]
  PIN r_data_o[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 65.835 94.11 65.905 ;
    END
  END r_data_o[304]
  PIN r_data_o[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 15.435 0.07 15.505 ;
    END
  END r_data_o[305]
  PIN r_data_o[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  81.785 140.02 81.925 140.16 ;
    END
  END r_data_o[306]
  PIN r_data_o[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 54.915 94.11 54.985 ;
    END
  END r_data_o[307]
  PIN r_data_o[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 114.275 0.07 114.345 ;
    END
  END r_data_o[308]
  PIN r_data_o[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 78.435 0.07 78.505 ;
    END
  END r_data_o[309]
  PIN r_data_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  38.105 0 38.245 0.14 ;
    END
  END r_data_o[30]
  PIN r_data_o[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 22.715 0.07 22.785 ;
    END
  END r_data_o[310]
  PIN r_data_o[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 8.435 94.11 8.505 ;
    END
  END r_data_o[311]
  PIN r_data_o[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 115.675 94.11 115.745 ;
    END
  END r_data_o[312]
  PIN r_data_o[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 137.795 94.11 137.865 ;
    END
  END r_data_o[313]
  PIN r_data_o[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 76.755 94.11 76.825 ;
    END
  END r_data_o[314]
  PIN r_data_o[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 98.315 94.11 98.385 ;
    END
  END r_data_o[315]
  PIN r_data_o[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 66.955 0.07 67.025 ;
    END
  END r_data_o[316]
  PIN r_data_o[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 10.115 94.11 10.185 ;
    END
  END r_data_o[317]
  PIN r_data_o[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  59.385 0 59.525 0.14 ;
    END
  END r_data_o[318]
  PIN r_data_o[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  55.465 0 55.605 0.14 ;
    END
  END r_data_o[319]
  PIN r_data_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 14.315 94.11 14.385 ;
    END
  END r_data_o[31]
  PIN r_data_o[320]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 106.155 94.11 106.225 ;
    END
  END r_data_o[320]
  PIN r_data_o[321]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 46.795 0.07 46.865 ;
    END
  END r_data_o[321]
  PIN r_data_o[322]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 101.395 0.07 101.465 ;
    END
  END r_data_o[322]
  PIN r_data_o[323]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 138.355 94.11 138.425 ;
    END
  END r_data_o[323]
  PIN r_data_o[324]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 89.635 94.11 89.705 ;
    END
  END r_data_o[324]
  PIN r_data_o[325]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 115.955 0.07 116.025 ;
    END
  END r_data_o[325]
  PIN r_data_o[326]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 117.355 94.11 117.425 ;
    END
  END r_data_o[326]
  PIN r_data_o[327]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 121.275 94.11 121.345 ;
    END
  END r_data_o[327]
  PIN r_data_o[328]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 56.595 0.07 56.665 ;
    END
  END r_data_o[328]
  PIN r_data_o[329]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  62.185 0 62.325 0.14 ;
    END
  END r_data_o[329]
  PIN r_data_o[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 80.115 94.11 80.185 ;
    END
  END r_data_o[32]
  PIN r_data_o[330]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 127.155 0.07 127.225 ;
    END
  END r_data_o[330]
  PIN r_data_o[331]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  59.945 140.02 60.085 140.16 ;
    END
  END r_data_o[331]
  PIN r_data_o[332]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 25.795 0.07 25.865 ;
    END
  END r_data_o[332]
  PIN r_data_o[333]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  86.825 0 86.965 0.14 ;
    END
  END r_data_o[333]
  PIN r_data_o[334]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 89.355 0.07 89.425 ;
    END
  END r_data_o[334]
  PIN r_data_o[335]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 63.035 0.07 63.105 ;
    END
  END r_data_o[335]
  PIN r_data_o[336]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 138.635 94.11 138.705 ;
    END
  END r_data_o[336]
  PIN r_data_o[337]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 96.075 94.11 96.145 ;
    END
  END r_data_o[337]
  PIN r_data_o[338]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 113.995 0.07 114.065 ;
    END
  END r_data_o[338]
  PIN r_data_o[339]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 33.915 0.07 33.985 ;
    END
  END r_data_o[339]
  PIN r_data_o[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 101.955 0.07 102.025 ;
    END
  END r_data_o[33]
  PIN r_data_o[340]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  38.665 0 38.805 0.14 ;
    END
  END r_data_o[340]
  PIN r_data_o[341]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 65.555 0.07 65.625 ;
    END
  END r_data_o[341]
  PIN r_data_o[342]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  75.065 0 75.205 0.14 ;
    END
  END r_data_o[342]
  PIN r_data_o[343]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.585 0 14.725 0.14 ;
    END
  END r_data_o[343]
  PIN r_data_o[344]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 122.675 94.11 122.745 ;
    END
  END r_data_o[344]
  PIN r_data_o[345]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 81.235 94.11 81.305 ;
    END
  END r_data_o[345]
  PIN r_data_o[346]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 31.395 94.11 31.465 ;
    END
  END r_data_o[346]
  PIN r_data_o[347]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 109.795 94.11 109.865 ;
    END
  END r_data_o[347]
  PIN r_data_o[348]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  85.705 140.02 85.845 140.16 ;
    END
  END r_data_o[348]
  PIN r_data_o[349]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 47.075 94.11 47.145 ;
    END
  END r_data_o[349]
  PIN r_data_o[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 29.995 0.07 30.065 ;
    END
  END r_data_o[34]
  PIN r_data_o[350]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 83.755 94.11 83.825 ;
    END
  END r_data_o[350]
  PIN r_data_o[351]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 110.075 94.11 110.145 ;
    END
  END r_data_o[351]
  PIN r_data_o[352]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 50.435 94.11 50.505 ;
    END
  END r_data_o[352]
  PIN r_data_o[353]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 133.875 94.11 133.945 ;
    END
  END r_data_o[353]
  PIN r_data_o[354]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 78.155 94.11 78.225 ;
    END
  END r_data_o[354]
  PIN r_data_o[355]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 99.715 94.11 99.785 ;
    END
  END r_data_o[355]
  PIN r_data_o[356]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 65.275 94.11 65.345 ;
    END
  END r_data_o[356]
  PIN r_data_o[357]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 43.155 0.07 43.225 ;
    END
  END r_data_o[357]
  PIN r_data_o[358]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.025 140.02 14.165 140.16 ;
    END
  END r_data_o[358]
  PIN r_data_o[359]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 48.755 94.11 48.825 ;
    END
  END r_data_o[359]
  PIN r_data_o[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 5.915 94.11 5.985 ;
    END
  END r_data_o[35]
  PIN r_data_o[360]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 61.355 0.07 61.425 ;
    END
  END r_data_o[360]
  PIN r_data_o[361]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.385 140.02 31.525 140.16 ;
    END
  END r_data_o[361]
  PIN r_data_o[362]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 90.755 94.11 90.825 ;
    END
  END r_data_o[362]
  PIN r_data_o[363]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 84.595 0.07 84.665 ;
    END
  END r_data_o[363]
  PIN r_data_o[364]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.905 140.02 13.045 140.16 ;
    END
  END r_data_o[364]
  PIN r_data_o[365]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.385 0 17.525 0.14 ;
    END
  END r_data_o[365]
  PIN r_data_o[366]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  21.865 0 22.005 0.14 ;
    END
  END r_data_o[366]
  PIN r_data_o[367]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 108.115 0.07 108.185 ;
    END
  END r_data_o[367]
  PIN r_data_o[368]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 29.995 94.11 30.065 ;
    END
  END r_data_o[368]
  PIN r_data_o[369]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 3.115 0.07 3.185 ;
    END
  END r_data_o[369]
  PIN r_data_o[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 99.435 94.11 99.505 ;
    END
  END r_data_o[36]
  PIN r_data_o[370]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 28.035 94.11 28.105 ;
    END
  END r_data_o[370]
  PIN r_data_o[371]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 72.835 94.11 72.905 ;
    END
  END r_data_o[371]
  PIN r_data_o[372]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 38.955 0.07 39.025 ;
    END
  END r_data_o[372]
  PIN r_data_o[373]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 137.515 94.11 137.585 ;
    END
  END r_data_o[373]
  PIN r_data_o[374]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  64.985 0 65.125 0.14 ;
    END
  END r_data_o[374]
  PIN r_data_o[375]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 40.355 0.07 40.425 ;
    END
  END r_data_o[375]
  PIN r_data_o[376]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 119.315 0.07 119.385 ;
    END
  END r_data_o[376]
  PIN r_data_o[377]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  33.625 140.02 33.765 140.16 ;
    END
  END r_data_o[377]
  PIN r_data_o[378]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 18.515 0.07 18.585 ;
    END
  END r_data_o[378]
  PIN r_data_o[379]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 10.395 0.07 10.465 ;
    END
  END r_data_o[379]
  PIN r_data_o[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 82.915 0.07 82.985 ;
    END
  END r_data_o[37]
  PIN r_data_o[380]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 72.555 94.11 72.625 ;
    END
  END r_data_o[380]
  PIN r_data_o[381]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 76.195 0.07 76.265 ;
    END
  END r_data_o[381]
  PIN r_data_o[382]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 3.395 94.11 3.465 ;
    END
  END r_data_o[382]
  PIN r_data_o[383]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 115.115 0.07 115.185 ;
    END
  END r_data_o[383]
  PIN r_data_o[384]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 68.355 0.07 68.425 ;
    END
  END r_data_o[384]
  PIN r_data_o[385]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  79.545 140.02 79.685 140.16 ;
    END
  END r_data_o[385]
  PIN r_data_o[386]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 11.515 0.07 11.585 ;
    END
  END r_data_o[386]
  PIN r_data_o[387]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  66.665 0 66.805 0.14 ;
    END
  END r_data_o[387]
  PIN r_data_o[388]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 52.395 0.07 52.465 ;
    END
  END r_data_o[388]
  PIN r_data_o[389]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 118.475 94.11 118.545 ;
    END
  END r_data_o[389]
  PIN r_data_o[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  77.865 140.02 78.005 140.16 ;
    END
  END r_data_o[38]
  PIN r_data_o[390]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 49.315 94.11 49.385 ;
    END
  END r_data_o[390]
  PIN r_data_o[391]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 55.195 94.11 55.265 ;
    END
  END r_data_o[391]
  PIN r_data_o[392]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  80.105 140.02 80.245 140.16 ;
    END
  END r_data_o[392]
  PIN r_data_o[393]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 135.835 94.11 135.905 ;
    END
  END r_data_o[393]
  PIN r_data_o[394]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  82.905 0 83.045 0.14 ;
    END
  END r_data_o[394]
  PIN r_data_o[395]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 105.875 0.07 105.945 ;
    END
  END r_data_o[395]
  PIN r_data_o[396]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  80.665 140.02 80.805 140.16 ;
    END
  END r_data_o[396]
  PIN r_data_o[397]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 80.955 0.07 81.025 ;
    END
  END r_data_o[397]
  PIN r_data_o[398]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  68.905 0 69.045 0.14 ;
    END
  END r_data_o[398]
  PIN r_data_o[399]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  87.385 140.02 87.525 140.16 ;
    END
  END r_data_o[399]
  PIN r_data_o[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 93.555 94.11 93.625 ;
    END
  END r_data_o[39]
  PIN r_data_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 133.595 0.07 133.665 ;
    END
  END r_data_o[3]
  PIN r_data_o[400]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 124.635 94.11 124.705 ;
    END
  END r_data_o[400]
  PIN r_data_o[401]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 42.315 0.07 42.385 ;
    END
  END r_data_o[401]
  PIN r_data_o[402]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 53.235 94.11 53.305 ;
    END
  END r_data_o[402]
  PIN r_data_o[403]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  83.465 0 83.605 0.14 ;
    END
  END r_data_o[403]
  PIN r_data_o[404]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  22.985 0 23.125 0.14 ;
    END
  END r_data_o[404]
  PIN r_data_o[405]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 105.035 94.11 105.105 ;
    END
  END r_data_o[405]
  PIN r_data_o[406]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 65.555 94.11 65.625 ;
    END
  END r_data_o[406]
  PIN r_data_o[407]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 124.075 0.07 124.145 ;
    END
  END r_data_o[407]
  PIN r_data_o[408]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 49.315 0.07 49.385 ;
    END
  END r_data_o[408]
  PIN r_data_o[409]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 66.395 0.07 66.465 ;
    END
  END r_data_o[409]
  PIN r_data_o[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 131.635 94.11 131.705 ;
    END
  END r_data_o[40]
  PIN r_data_o[410]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  70.025 140.02 70.165 140.16 ;
    END
  END r_data_o[410]
  PIN r_data_o[411]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 44.275 0.07 44.345 ;
    END
  END r_data_o[411]
  PIN r_data_o[412]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 101.395 94.11 101.465 ;
    END
  END r_data_o[412]
  PIN r_data_o[413]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 106.715 0.07 106.785 ;
    END
  END r_data_o[413]
  PIN r_data_o[414]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 103.355 0.07 103.425 ;
    END
  END r_data_o[414]
  PIN r_data_o[415]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 135.555 0.07 135.625 ;
    END
  END r_data_o[415]
  PIN r_data_o[416]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 20.475 94.11 20.545 ;
    END
  END r_data_o[416]
  PIN r_data_o[417]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 116.235 94.11 116.305 ;
    END
  END r_data_o[417]
  PIN r_data_o[418]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 118.475 0.07 118.545 ;
    END
  END r_data_o[418]
  PIN r_data_o[419]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 112.875 0.07 112.945 ;
    END
  END r_data_o[419]
  PIN r_data_o[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 103.915 94.11 103.985 ;
    END
  END r_data_o[41]
  PIN r_data_o[420]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 1.995 94.11 2.065 ;
    END
  END r_data_o[420]
  PIN r_data_o[421]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  11.225 140.02 11.365 140.16 ;
    END
  END r_data_o[421]
  PIN r_data_o[422]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 69.755 94.11 69.825 ;
    END
  END r_data_o[422]
  PIN r_data_o[423]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 139.195 0.07 139.265 ;
    END
  END r_data_o[423]
  PIN r_data_o[424]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 78.715 0.07 78.785 ;
    END
  END r_data_o[424]
  PIN r_data_o[425]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 21.035 94.11 21.105 ;
    END
  END r_data_o[425]
  PIN r_data_o[426]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 74.795 94.11 74.865 ;
    END
  END r_data_o[426]
  PIN r_data_o[427]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  28.585 140.02 28.725 140.16 ;
    END
  END r_data_o[427]
  PIN r_data_o[428]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  42.025 0 42.165 0.14 ;
    END
  END r_data_o[428]
  PIN r_data_o[429]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 38.115 0.07 38.185 ;
    END
  END r_data_o[429]
  PIN r_data_o[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  67.225 0 67.365 0.14 ;
    END
  END r_data_o[42]
  PIN r_data_o[430]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  43.705 140.02 43.845 140.16 ;
    END
  END r_data_o[430]
  PIN r_data_o[431]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 95.235 94.11 95.305 ;
    END
  END r_data_o[431]
  PIN r_data_o[432]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 4.515 94.11 4.585 ;
    END
  END r_data_o[432]
  PIN r_data_o[433]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 42.875 94.11 42.945 ;
    END
  END r_data_o[433]
  PIN r_data_o[434]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 48.195 0.07 48.265 ;
    END
  END r_data_o[434]
  PIN r_data_o[435]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 60.795 94.11 60.865 ;
    END
  END r_data_o[435]
  PIN r_data_o[436]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 35.595 0.07 35.665 ;
    END
  END r_data_o[436]
  PIN r_data_o[437]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 9.555 0.07 9.625 ;
    END
  END r_data_o[437]
  PIN r_data_o[438]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 78.995 94.11 79.065 ;
    END
  END r_data_o[438]
  PIN r_data_o[439]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 122.395 94.11 122.465 ;
    END
  END r_data_o[439]
  PIN r_data_o[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 39.235 94.11 39.305 ;
    END
  END r_data_o[43]
  PIN r_data_o[440]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 28.035 0.07 28.105 ;
    END
  END r_data_o[440]
  PIN r_data_o[441]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  48.185 140.02 48.325 140.16 ;
    END
  END r_data_o[441]
  PIN r_data_o[442]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  53.785 140.02 53.925 140.16 ;
    END
  END r_data_o[442]
  PIN r_data_o[443]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  64.425 0 64.565 0.14 ;
    END
  END r_data_o[443]
  PIN r_data_o[444]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 115.675 0.07 115.745 ;
    END
  END r_data_o[444]
  PIN r_data_o[445]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  27.465 140.02 27.605 140.16 ;
    END
  END r_data_o[445]
  PIN r_data_o[446]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  5.625 0 5.765 0.14 ;
    END
  END r_data_o[446]
  PIN r_data_o[447]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 39.515 94.11 39.585 ;
    END
  END r_data_o[447]
  PIN r_data_o[448]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 105.315 94.11 105.385 ;
    END
  END r_data_o[448]
  PIN r_data_o[449]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 2.555 94.11 2.625 ;
    END
  END r_data_o[449]
  PIN r_data_o[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  80.665 0 80.805 0.14 ;
    END
  END r_data_o[44]
  PIN r_data_o[450]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 93.835 0.07 93.905 ;
    END
  END r_data_o[450]
  PIN r_data_o[451]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 84.595 94.11 84.665 ;
    END
  END r_data_o[451]
  PIN r_data_o[452]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  86.265 0 86.405 0.14 ;
    END
  END r_data_o[452]
  PIN r_data_o[453]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  18.505 140.02 18.645 140.16 ;
    END
  END r_data_o[453]
  PIN r_data_o[454]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 33.355 94.11 33.425 ;
    END
  END r_data_o[454]
  PIN r_data_o[455]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  24.105 0 24.245 0.14 ;
    END
  END r_data_o[455]
  PIN r_data_o[456]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  89.625 140.02 89.765 140.16 ;
    END
  END r_data_o[456]
  PIN r_data_o[457]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  38.665 140.02 38.805 140.16 ;
    END
  END r_data_o[457]
  PIN r_data_o[458]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 109.515 0.07 109.585 ;
    END
  END r_data_o[458]
  PIN r_data_o[459]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  57.145 140.02 57.285 140.16 ;
    END
  END r_data_o[459]
  PIN r_data_o[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 57.435 0.07 57.505 ;
    END
  END r_data_o[45]
  PIN r_data_o[460]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 129.395 94.11 129.465 ;
    END
  END r_data_o[460]
  PIN r_data_o[461]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  71.705 0 71.845 0.14 ;
    END
  END r_data_o[461]
  PIN r_data_o[462]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  51.545 0 51.685 0.14 ;
    END
  END r_data_o[462]
  PIN r_data_o[463]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  54.345 0 54.485 0.14 ;
    END
  END r_data_o[463]
  PIN r_data_o[464]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 85.435 0.07 85.505 ;
    END
  END r_data_o[464]
  PIN r_data_o[465]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 57.995 0.07 58.065 ;
    END
  END r_data_o[465]
  PIN r_data_o[466]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 81.515 94.11 81.585 ;
    END
  END r_data_o[466]
  PIN r_data_o[467]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 63.035 94.11 63.105 ;
    END
  END r_data_o[467]
  PIN r_data_o[468]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 102.235 94.11 102.305 ;
    END
  END r_data_o[468]
  PIN r_data_o[469]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 37.835 94.11 37.905 ;
    END
  END r_data_o[469]
  PIN r_data_o[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 79.835 94.11 79.905 ;
    END
  END r_data_o[46]
  PIN r_data_o[470]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 125.475 0.07 125.545 ;
    END
  END r_data_o[470]
  PIN r_data_o[471]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 123.235 94.11 123.305 ;
    END
  END r_data_o[471]
  PIN r_data_o[472]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 36.995 0.07 37.065 ;
    END
  END r_data_o[472]
  PIN r_data_o[473]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 89.075 0.07 89.145 ;
    END
  END r_data_o[473]
  PIN r_data_o[474]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  91.305 140.02 91.445 140.16 ;
    END
  END r_data_o[474]
  PIN r_data_o[475]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 41.195 94.11 41.265 ;
    END
  END r_data_o[475]
  PIN r_data_o[476]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 32.235 94.11 32.305 ;
    END
  END r_data_o[476]
  PIN r_data_o[477]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 7.315 94.11 7.385 ;
    END
  END r_data_o[477]
  PIN r_data_o[478]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 46.515 0.07 46.585 ;
    END
  END r_data_o[478]
  PIN r_data_o[479]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  39.225 140.02 39.365 140.16 ;
    END
  END r_data_o[479]
  PIN r_data_o[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 128.275 0.07 128.345 ;
    END
  END r_data_o[47]
  PIN r_data_o[480]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 83.475 94.11 83.545 ;
    END
  END r_data_o[480]
  PIN r_data_o[481]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 112.315 94.11 112.385 ;
    END
  END r_data_o[481]
  PIN r_data_o[482]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 35.035 94.11 35.105 ;
    END
  END r_data_o[482]
  PIN r_data_o[483]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 103.075 94.11 103.145 ;
    END
  END r_data_o[483]
  PIN r_data_o[484]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.305 0 7.445 0.14 ;
    END
  END r_data_o[484]
  PIN r_data_o[485]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 85.715 94.11 85.785 ;
    END
  END r_data_o[485]
  PIN r_data_o[486]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 97.475 94.11 97.545 ;
    END
  END r_data_o[486]
  PIN r_data_o[487]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  16.825 140.02 16.965 140.16 ;
    END
  END r_data_o[487]
  PIN r_data_o[488]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  19.625 0 19.765 0.14 ;
    END
  END r_data_o[488]
  PIN r_data_o[489]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 117.915 0.07 117.985 ;
    END
  END r_data_o[489]
  PIN r_data_o[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 126.315 94.11 126.385 ;
    END
  END r_data_o[48]
  PIN r_data_o[490]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  74.505 140.02 74.645 140.16 ;
    END
  END r_data_o[490]
  PIN r_data_o[491]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 132.475 94.11 132.545 ;
    END
  END r_data_o[491]
  PIN r_data_o[492]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 19.355 0.07 19.425 ;
    END
  END r_data_o[492]
  PIN r_data_o[493]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 5.915 0.07 5.985 ;
    END
  END r_data_o[493]
  PIN r_data_o[494]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 25.235 94.11 25.305 ;
    END
  END r_data_o[494]
  PIN r_data_o[495]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  63.305 140.02 63.445 140.16 ;
    END
  END r_data_o[495]
  PIN r_data_o[496]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 29.435 0.07 29.505 ;
    END
  END r_data_o[496]
  PIN r_data_o[497]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 30.555 0.07 30.625 ;
    END
  END r_data_o[497]
  PIN r_data_o[498]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 131.075 0.07 131.145 ;
    END
  END r_data_o[498]
  PIN r_data_o[499]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 44.835 0.07 44.905 ;
    END
  END r_data_o[499]
  PIN r_data_o[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 49.875 0.07 49.945 ;
    END
  END r_data_o[49]
  PIN r_data_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 134.995 94.11 135.065 ;
    END
  END r_data_o[4]
  PIN r_data_o[500]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.665 140.02 10.805 140.16 ;
    END
  END r_data_o[500]
  PIN r_data_o[501]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 80.395 0.07 80.465 ;
    END
  END r_data_o[501]
  PIN r_data_o[502]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 85.715 0.07 85.785 ;
    END
  END r_data_o[502]
  PIN r_data_o[503]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 48.475 0.07 48.545 ;
    END
  END r_data_o[503]
  PIN r_data_o[504]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 107.275 94.11 107.345 ;
    END
  END r_data_o[504]
  PIN r_data_o[505]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 12.635 94.11 12.705 ;
    END
  END r_data_o[505]
  PIN r_data_o[506]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 67.235 0.07 67.305 ;
    END
  END r_data_o[506]
  PIN r_data_o[507]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 17.955 94.11 18.025 ;
    END
  END r_data_o[507]
  PIN r_data_o[508]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 71.155 0.07 71.225 ;
    END
  END r_data_o[508]
  PIN r_data_o[509]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 117.635 94.11 117.705 ;
    END
  END r_data_o[509]
  PIN r_data_o[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 5.635 94.11 5.705 ;
    END
  END r_data_o[50]
  PIN r_data_o[510]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  90.185 140.02 90.325 140.16 ;
    END
  END r_data_o[510]
  PIN r_data_o[511]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 74.515 94.11 74.585 ;
    END
  END r_data_o[511]
  PIN r_data_o[512]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 95.515 0.07 95.585 ;
    END
  END r_data_o[512]
  PIN r_data_o[513]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 68.355 94.11 68.425 ;
    END
  END r_data_o[513]
  PIN r_data_o[514]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  29.705 0 29.845 0.14 ;
    END
  END r_data_o[514]
  PIN r_data_o[515]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.355 0.07 12.425 ;
    END
  END r_data_o[515]
  PIN r_data_o[516]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 36.155 0.07 36.225 ;
    END
  END r_data_o[516]
  PIN r_data_o[517]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  52.665 0 52.805 0.14 ;
    END
  END r_data_o[517]
  PIN r_data_o[518]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 63.315 0.07 63.385 ;
    END
  END r_data_o[518]
  PIN r_data_o[519]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 134.435 94.11 134.505 ;
    END
  END r_data_o[519]
  PIN r_data_o[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 15.995 0.07 16.065 ;
    END
  END r_data_o[51]
  PIN r_data_o[520]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 71.435 0.07 71.505 ;
    END
  END r_data_o[520]
  PIN r_data_o[521]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.905 0 13.045 0.14 ;
    END
  END r_data_o[521]
  PIN r_data_o[522]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  29.145 0 29.285 0.14 ;
    END
  END r_data_o[522]
  PIN r_data_o[523]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 127.995 0.07 128.065 ;
    END
  END r_data_o[523]
  PIN r_data_o[524]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  59.385 140.02 59.525 140.16 ;
    END
  END r_data_o[524]
  PIN r_data_o[525]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  35.865 0 36.005 0.14 ;
    END
  END r_data_o[525]
  PIN r_data_o[526]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 119.035 0.07 119.105 ;
    END
  END r_data_o[526]
  PIN r_data_o[527]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 1.435 0.07 1.505 ;
    END
  END r_data_o[527]
  PIN r_data_o[528]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  37.545 0 37.685 0.14 ;
    END
  END r_data_o[528]
  PIN r_data_o[529]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 71.715 94.11 71.785 ;
    END
  END r_data_o[529]
  PIN r_data_o[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  48.745 0 48.885 0.14 ;
    END
  END r_data_o[52]
  PIN r_data_o[530]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  51.545 140.02 51.685 140.16 ;
    END
  END r_data_o[530]
  PIN r_data_o[531]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 26.635 0.07 26.705 ;
    END
  END r_data_o[531]
  PIN r_data_o[532]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  77.305 0 77.445 0.14 ;
    END
  END r_data_o[532]
  PIN r_data_o[533]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 64.715 0.07 64.785 ;
    END
  END r_data_o[533]
  PIN r_data_o[534]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 81.515 0.07 81.585 ;
    END
  END r_data_o[534]
  PIN r_data_o[535]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 119.595 94.11 119.665 ;
    END
  END r_data_o[535]
  PIN r_data_o[536]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 133.595 94.11 133.665 ;
    END
  END r_data_o[536]
  PIN r_data_o[537]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 92.435 0.07 92.505 ;
    END
  END r_data_o[537]
  PIN r_data_o[538]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 42.035 94.11 42.105 ;
    END
  END r_data_o[538]
  PIN r_data_o[539]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 138.355 0.07 138.425 ;
    END
  END r_data_o[539]
  PIN r_data_o[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 42.035 0.07 42.105 ;
    END
  END r_data_o[53]
  PIN r_data_o[540]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 36.435 94.11 36.505 ;
    END
  END r_data_o[540]
  PIN r_data_o[541]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.745 140.02 34.885 140.16 ;
    END
  END r_data_o[541]
  PIN r_data_o[542]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 90.755 0.07 90.825 ;
    END
  END r_data_o[542]
  PIN r_data_o[543]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  90.185 0 90.325 0.14 ;
    END
  END r_data_o[543]
  PIN r_data_o[544]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 3.955 0.07 4.025 ;
    END
  END r_data_o[544]
  PIN r_data_o[545]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 60.515 94.11 60.585 ;
    END
  END r_data_o[545]
  PIN r_data_o[546]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 37.555 0.07 37.625 ;
    END
  END r_data_o[546]
  PIN r_data_o[547]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  58.825 140.02 58.965 140.16 ;
    END
  END r_data_o[547]
  PIN r_data_o[548]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  50.985 140.02 51.125 140.16 ;
    END
  END r_data_o[548]
  PIN r_data_o[549]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 43.155 94.11 43.225 ;
    END
  END r_data_o[549]
  PIN r_data_o[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  78.425 0 78.565 0.14 ;
    END
  END r_data_o[54]
  PIN r_data_o[550]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  1.145 140.02 1.285 140.16 ;
    END
  END r_data_o[550]
  PIN r_data_o[551]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 26.355 94.11 26.425 ;
    END
  END r_data_o[551]
  PIN r_data_o[552]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  50.985 0 51.125 0.14 ;
    END
  END r_data_o[552]
  PIN r_data_o[553]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 104.195 94.11 104.265 ;
    END
  END r_data_o[553]
  PIN r_data_o[554]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 112.315 0.07 112.385 ;
    END
  END r_data_o[554]
  PIN r_data_o[555]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.075 0.07 12.145 ;
    END
  END r_data_o[555]
  PIN r_data_o[556]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 21.595 94.11 21.665 ;
    END
  END r_data_o[556]
  PIN r_data_o[557]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 103.075 0.07 103.145 ;
    END
  END r_data_o[557]
  PIN r_data_o[558]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 69.195 94.11 69.265 ;
    END
  END r_data_o[558]
  PIN r_data_o[559]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 91.595 0.07 91.665 ;
    END
  END r_data_o[559]
  PIN r_data_o[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  71.145 140.02 71.285 140.16 ;
    END
  END r_data_o[55]
  PIN r_data_o[560]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  84.025 140.02 84.165 140.16 ;
    END
  END r_data_o[560]
  PIN r_data_o[561]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 114.555 94.11 114.625 ;
    END
  END r_data_o[561]
  PIN r_data_o[562]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  61.625 0 61.765 0.14 ;
    END
  END r_data_o[562]
  PIN r_data_o[563]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 77.875 0.07 77.945 ;
    END
  END r_data_o[563]
  PIN r_data_o[564]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.035 0.07 7.105 ;
    END
  END r_data_o[564]
  PIN r_data_o[565]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  26.345 0 26.485 0.14 ;
    END
  END r_data_o[565]
  PIN r_data_o[566]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 126.595 94.11 126.665 ;
    END
  END r_data_o[566]
  PIN r_data_o[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 28.315 94.11 28.385 ;
    END
  END r_data_o[56]
  PIN r_data_o[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 27.195 94.11 27.265 ;
    END
  END r_data_o[57]
  PIN r_data_o[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  91.865 0 92.005 0.14 ;
    END
  END r_data_o[58]
  PIN r_data_o[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 1.995 0.07 2.065 ;
    END
  END r_data_o[59]
  PIN r_data_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 89.355 94.11 89.425 ;
    END
  END r_data_o[5]
  PIN r_data_o[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 96.075 0.07 96.145 ;
    END
  END r_data_o[60]
  PIN r_data_o[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 77.035 0.07 77.105 ;
    END
  END r_data_o[61]
  PIN r_data_o[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 77.315 0.07 77.385 ;
    END
  END r_data_o[62]
  PIN r_data_o[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 29.715 0.07 29.785 ;
    END
  END r_data_o[63]
  PIN r_data_o[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 120.435 94.11 120.505 ;
    END
  END r_data_o[64]
  PIN r_data_o[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 105.595 0.07 105.665 ;
    END
  END r_data_o[65]
  PIN r_data_o[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 72.275 0.07 72.345 ;
    END
  END r_data_o[66]
  PIN r_data_o[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 79.555 94.11 79.625 ;
    END
  END r_data_o[67]
  PIN r_data_o[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 60.795 0.07 60.865 ;
    END
  END r_data_o[68]
  PIN r_data_o[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 11.795 0.07 11.865 ;
    END
  END r_data_o[69]
  PIN r_data_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 75.635 94.11 75.705 ;
    END
  END r_data_o[6]
  PIN r_data_o[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 48.195 94.11 48.265 ;
    END
  END r_data_o[70]
  PIN r_data_o[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 137.235 0.07 137.305 ;
    END
  END r_data_o[71]
  PIN r_data_o[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 46.795 94.11 46.865 ;
    END
  END r_data_o[72]
  PIN r_data_o[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 64.435 0.07 64.505 ;
    END
  END r_data_o[73]
  PIN r_data_o[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 97.475 0.07 97.545 ;
    END
  END r_data_o[74]
  PIN r_data_o[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 101.955 94.11 102.025 ;
    END
  END r_data_o[75]
  PIN r_data_o[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 38.675 0.07 38.745 ;
    END
  END r_data_o[76]
  PIN r_data_o[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 74.515 0.07 74.585 ;
    END
  END r_data_o[77]
  PIN r_data_o[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 63.875 94.11 63.945 ;
    END
  END r_data_o[78]
  PIN r_data_o[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 67.515 0.07 67.585 ;
    END
  END r_data_o[79]
  PIN r_data_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.185 140.02 34.325 140.16 ;
    END
  END r_data_o[7]
  PIN r_data_o[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 73.115 0.07 73.185 ;
    END
  END r_data_o[80]
  PIN r_data_o[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 91.035 94.11 91.105 ;
    END
  END r_data_o[81]
  PIN r_data_o[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 58.835 0.07 58.905 ;
    END
  END r_data_o[82]
  PIN r_data_o[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 47.355 94.11 47.425 ;
    END
  END r_data_o[83]
  PIN r_data_o[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 75.635 0.07 75.705 ;
    END
  END r_data_o[84]
  PIN r_data_o[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 124.355 0.07 124.425 ;
    END
  END r_data_o[85]
  PIN r_data_o[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 50.715 94.11 50.785 ;
    END
  END r_data_o[86]
  PIN r_data_o[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 98.595 0.07 98.665 ;
    END
  END r_data_o[87]
  PIN r_data_o[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 131.915 0.07 131.985 ;
    END
  END r_data_o[88]
  PIN r_data_o[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  6.745 140.02 6.885 140.16 ;
    END
  END r_data_o[89]
  PIN r_data_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.025 0 14.165 0.14 ;
    END
  END r_data_o[8]
  PIN r_data_o[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 99.435 0.07 99.505 ;
    END
  END r_data_o[90]
  PIN r_data_o[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  90.745 0 90.885 0.14 ;
    END
  END r_data_o[91]
  PIN r_data_o[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 8.155 0.07 8.225 ;
    END
  END r_data_o[92]
  PIN r_data_o[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 110.635 94.11 110.705 ;
    END
  END r_data_o[93]
  PIN r_data_o[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  90.745 140.02 90.885 140.16 ;
    END
  END r_data_o[94]
  PIN r_data_o[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 107.555 94.11 107.625 ;
    END
  END r_data_o[95]
  PIN r_data_o[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 6.475 94.11 6.545 ;
    END
  END r_data_o[96]
  PIN r_data_o[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 134.155 94.11 134.225 ;
    END
  END r_data_o[97]
  PIN r_data_o[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 128.555 0.07 128.625 ;
    END
  END r_data_o[98]
  PIN r_data_o[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  56.585 0 56.725 0.14 ;
    END
  END r_data_o[99]
  PIN r_data_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 40.075 94.11 40.145 ;
    END
  END r_data_o[9]
  PIN r_v_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 14.595 94.11 14.665 ;
    END
  END r_v_i
  PIN w_addr_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  13.465 0 13.605 0.14 ;
    END
  END w_addr_i
  PIN w_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 78.715 94.11 78.785 ;
    END
  END w_clk_i
  PIN w_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 61.355 94.11 61.425 ;
    END
  END w_data_i[0]
  PIN w_data_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 104.195 0.07 104.265 ;
    END
  END w_data_i[100]
  PIN w_data_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.745 0 34.885 0.14 ;
    END
  END w_data_i[101]
  PIN w_data_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 39.235 0.07 39.305 ;
    END
  END w_data_i[102]
  PIN w_data_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 92.715 0.07 92.785 ;
    END
  END w_data_i[103]
  PIN w_data_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 45.675 0.07 45.745 ;
    END
  END w_data_i[104]
  PIN w_data_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 72.835 0.07 72.905 ;
    END
  END w_data_i[105]
  PIN w_data_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 120.715 94.11 120.785 ;
    END
  END w_data_i[106]
  PIN w_data_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 41.755 0.07 41.825 ;
    END
  END w_data_i[107]
  PIN w_data_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 66.115 0.07 66.185 ;
    END
  END w_data_i[108]
  PIN w_data_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 104.475 94.11 104.545 ;
    END
  END w_data_i[109]
  PIN w_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 20.195 0.07 20.265 ;
    END
  END w_data_i[10]
  PIN w_data_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 87.115 94.11 87.185 ;
    END
  END w_data_i[110]
  PIN w_data_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  26.905 0 27.045 0.14 ;
    END
  END w_data_i[111]
  PIN w_data_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 82.355 0.07 82.425 ;
    END
  END w_data_i[112]
  PIN w_data_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 59.395 0.07 59.465 ;
    END
  END w_data_i[113]
  PIN w_data_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 36.715 0.07 36.785 ;
    END
  END w_data_i[114]
  PIN w_data_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  45.385 140.02 45.525 140.16 ;
    END
  END w_data_i[115]
  PIN w_data_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 125.755 0.07 125.825 ;
    END
  END w_data_i[116]
  PIN w_data_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 136.115 0.07 136.185 ;
    END
  END w_data_i[117]
  PIN w_data_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 55.475 0.07 55.545 ;
    END
  END w_data_i[118]
  PIN w_data_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 52.115 0.07 52.185 ;
    END
  END w_data_i[119]
  PIN w_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 111.475 0.07 111.545 ;
    END
  END w_data_i[11]
  PIN w_data_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 71.995 94.11 72.065 ;
    END
  END w_data_i[120]
  PIN w_data_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 93.555 0.07 93.625 ;
    END
  END w_data_i[121]
  PIN w_data_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 3.675 94.11 3.745 ;
    END
  END w_data_i[122]
  PIN w_data_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.385 140.02 17.525 140.16 ;
    END
  END w_data_i[123]
  PIN w_data_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 35.875 94.11 35.945 ;
    END
  END w_data_i[124]
  PIN w_data_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.595 0.07 21.665 ;
    END
  END w_data_i[125]
  PIN w_data_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 12.075 94.11 12.145 ;
    END
  END w_data_i[126]
  PIN w_data_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 120.995 0.07 121.065 ;
    END
  END w_data_i[127]
  PIN w_data_i[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  29.705 140.02 29.845 140.16 ;
    END
  END w_data_i[128]
  PIN w_data_i[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.955 0.07 32.025 ;
    END
  END w_data_i[129]
  PIN w_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 60.515 0.07 60.585 ;
    END
  END w_data_i[12]
  PIN w_data_i[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 122.395 0.07 122.465 ;
    END
  END w_data_i[130]
  PIN w_data_i[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  53.785 0 53.925 0.14 ;
    END
  END w_data_i[131]
  PIN w_data_i[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 46.235 0.07 46.305 ;
    END
  END w_data_i[132]
  PIN w_data_i[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 106.155 0.07 106.225 ;
    END
  END w_data_i[133]
  PIN w_data_i[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  25.785 140.02 25.925 140.16 ;
    END
  END w_data_i[134]
  PIN w_data_i[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 48.755 0.07 48.825 ;
    END
  END w_data_i[135]
  PIN w_data_i[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 128.275 94.11 128.345 ;
    END
  END w_data_i[136]
  PIN w_data_i[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 12.915 94.11 12.985 ;
    END
  END w_data_i[137]
  PIN w_data_i[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 57.435 94.11 57.505 ;
    END
  END w_data_i[138]
  PIN w_data_i[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 4.795 94.11 4.865 ;
    END
  END w_data_i[139]
  PIN w_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  56.025 0 56.165 0.14 ;
    END
  END w_data_i[13]
  PIN w_data_i[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 26.075 94.11 26.145 ;
    END
  END w_data_i[140]
  PIN w_data_i[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  66.665 140.02 66.805 140.16 ;
    END
  END w_data_i[141]
  PIN w_data_i[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 18.235 0.07 18.305 ;
    END
  END w_data_i[142]
  PIN w_data_i[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 126.035 0.07 126.105 ;
    END
  END w_data_i[143]
  PIN w_data_i[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 68.915 0.07 68.985 ;
    END
  END w_data_i[144]
  PIN w_data_i[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  39.225 0 39.365 0.14 ;
    END
  END w_data_i[145]
  PIN w_data_i[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 97.195 0.07 97.265 ;
    END
  END w_data_i[146]
  PIN w_data_i[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 69.475 94.11 69.545 ;
    END
  END w_data_i[147]
  PIN w_data_i[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.945 140.02 18.085 140.16 ;
    END
  END w_data_i[148]
  PIN w_data_i[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 95.515 94.11 95.585 ;
    END
  END w_data_i[149]
  PIN w_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 126.035 94.11 126.105 ;
    END
  END w_data_i[14]
  PIN w_data_i[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  82.345 140.02 82.485 140.16 ;
    END
  END w_data_i[150]
  PIN w_data_i[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 34.755 94.11 34.825 ;
    END
  END w_data_i[151]
  PIN w_data_i[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  3.385 140.02 3.525 140.16 ;
    END
  END w_data_i[152]
  PIN w_data_i[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 87.115 0.07 87.185 ;
    END
  END w_data_i[153]
  PIN w_data_i[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 45.955 0.07 46.025 ;
    END
  END w_data_i[154]
  PIN w_data_i[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 54.075 94.11 54.145 ;
    END
  END w_data_i[155]
  PIN w_data_i[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 101.675 0.07 101.745 ;
    END
  END w_data_i[156]
  PIN w_data_i[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 9.555 94.11 9.625 ;
    END
  END w_data_i[157]
  PIN w_data_i[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 129.955 94.11 130.025 ;
    END
  END w_data_i[158]
  PIN w_data_i[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 108.675 0.07 108.745 ;
    END
  END w_data_i[159]
  PIN w_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 25.515 0.07 25.585 ;
    END
  END w_data_i[15]
  PIN w_data_i[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 103.635 0.07 103.705 ;
    END
  END w_data_i[160]
  PIN w_data_i[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 15.435 94.11 15.505 ;
    END
  END w_data_i[161]
  PIN w_data_i[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.385 0 31.525 0.14 ;
    END
  END w_data_i[162]
  PIN w_data_i[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 131.915 94.11 131.985 ;
    END
  END w_data_i[163]
  PIN w_data_i[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  54.345 140.02 54.485 140.16 ;
    END
  END w_data_i[164]
  PIN w_data_i[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  41.465 140.02 41.605 140.16 ;
    END
  END w_data_i[165]
  PIN w_data_i[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 73.955 94.11 74.025 ;
    END
  END w_data_i[166]
  PIN w_data_i[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  58.265 140.02 58.405 140.16 ;
    END
  END w_data_i[167]
  PIN w_data_i[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 70.035 94.11 70.105 ;
    END
  END w_data_i[168]
  PIN w_data_i[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 44.275 94.11 44.345 ;
    END
  END w_data_i[169]
  PIN w_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 23.835 94.11 23.905 ;
    END
  END w_data_i[16]
  PIN w_data_i[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 23.555 0.07 23.625 ;
    END
  END w_data_i[170]
  PIN w_data_i[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 62.195 0.07 62.265 ;
    END
  END w_data_i[171]
  PIN w_data_i[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  6.745 0 6.885 0.14 ;
    END
  END w_data_i[172]
  PIN w_data_i[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 112.595 94.11 112.665 ;
    END
  END w_data_i[173]
  PIN w_data_i[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 73.675 0.07 73.745 ;
    END
  END w_data_i[174]
  PIN w_data_i[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 130.235 0.07 130.305 ;
    END
  END w_data_i[175]
  PIN w_data_i[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  73.945 140.02 74.085 140.16 ;
    END
  END w_data_i[176]
  PIN w_data_i[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.585 140.02 14.725 140.16 ;
    END
  END w_data_i[177]
  PIN w_data_i[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 121.835 0.07 121.905 ;
    END
  END w_data_i[178]
  PIN w_data_i[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 54.635 94.11 54.705 ;
    END
  END w_data_i[179]
  PIN w_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  61.065 140.02 61.205 140.16 ;
    END
  END w_data_i[17]
  PIN w_data_i[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 130.515 0.07 130.585 ;
    END
  END w_data_i[180]
  PIN w_data_i[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  76.185 0 76.325 0.14 ;
    END
  END w_data_i[181]
  PIN w_data_i[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  18.505 0 18.645 0.14 ;
    END
  END w_data_i[182]
  PIN w_data_i[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 93.275 94.11 93.345 ;
    END
  END w_data_i[183]
  PIN w_data_i[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 120.155 94.11 120.225 ;
    END
  END w_data_i[184]
  PIN w_data_i[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.665 0 10.805 0.14 ;
    END
  END w_data_i[185]
  PIN w_data_i[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 77.875 94.11 77.945 ;
    END
  END w_data_i[186]
  PIN w_data_i[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 70.875 0.07 70.945 ;
    END
  END w_data_i[187]
  PIN w_data_i[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 11.235 0.07 11.305 ;
    END
  END w_data_i[188]
  PIN w_data_i[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 111.475 94.11 111.545 ;
    END
  END w_data_i[189]
  PIN w_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 4.235 94.11 4.305 ;
    END
  END w_data_i[18]
  PIN w_data_i[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  85.145 0 85.285 0.14 ;
    END
  END w_data_i[190]
  PIN w_data_i[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  86.265 140.02 86.405 140.16 ;
    END
  END w_data_i[191]
  PIN w_data_i[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 61.635 94.11 61.705 ;
    END
  END w_data_i[192]
  PIN w_data_i[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 100.835 94.11 100.905 ;
    END
  END w_data_i[193]
  PIN w_data_i[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 80.675 94.11 80.745 ;
    END
  END w_data_i[194]
  PIN w_data_i[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 106.995 0.07 107.065 ;
    END
  END w_data_i[195]
  PIN w_data_i[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 64.715 94.11 64.785 ;
    END
  END w_data_i[196]
  PIN w_data_i[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 31.115 94.11 31.185 ;
    END
  END w_data_i[197]
  PIN w_data_i[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 58.555 0.07 58.625 ;
    END
  END w_data_i[198]
  PIN w_data_i[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 87.395 0.07 87.465 ;
    END
  END w_data_i[199]
  PIN w_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 93.835 94.11 93.905 ;
    END
  END w_data_i[19]
  PIN w_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  62.185 140.02 62.325 140.16 ;
    END
  END w_data_i[1]
  PIN w_data_i[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  67.225 140.02 67.365 140.16 ;
    END
  END w_data_i[200]
  PIN w_data_i[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 62.475 94.11 62.545 ;
    END
  END w_data_i[201]
  PIN w_data_i[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 2.555 0.07 2.625 ;
    END
  END w_data_i[202]
  PIN w_data_i[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 63.595 0.07 63.665 ;
    END
  END w_data_i[203]
  PIN w_data_i[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 129.115 0.07 129.185 ;
    END
  END w_data_i[204]
  PIN w_data_i[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 116.235 0.07 116.305 ;
    END
  END w_data_i[205]
  PIN w_data_i[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  2.825 140.02 2.965 140.16 ;
    END
  END w_data_i[206]
  PIN w_data_i[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 10.395 94.11 10.465 ;
    END
  END w_data_i[207]
  PIN w_data_i[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.315 0.07 21.385 ;
    END
  END w_data_i[208]
  PIN w_data_i[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 97.195 94.11 97.265 ;
    END
  END w_data_i[209]
  PIN w_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 36.995 94.11 37.065 ;
    END
  END w_data_i[20]
  PIN w_data_i[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 68.915 94.11 68.985 ;
    END
  END w_data_i[210]
  PIN w_data_i[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 5.075 0.07 5.145 ;
    END
  END w_data_i[211]
  PIN w_data_i[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 77.035 94.11 77.105 ;
    END
  END w_data_i[212]
  PIN w_data_i[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 22.435 0.07 22.505 ;
    END
  END w_data_i[213]
  PIN w_data_i[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 24.115 94.11 24.185 ;
    END
  END w_data_i[214]
  PIN w_data_i[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 103.635 94.11 103.705 ;
    END
  END w_data_i[215]
  PIN w_data_i[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 19.635 0.07 19.705 ;
    END
  END w_data_i[216]
  PIN w_data_i[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 92.995 0.07 93.065 ;
    END
  END w_data_i[217]
  PIN w_data_i[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 27.755 0.07 27.825 ;
    END
  END w_data_i[218]
  PIN w_data_i[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 102.515 94.11 102.585 ;
    END
  END w_data_i[219]
  PIN w_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 38.115 94.11 38.185 ;
    END
  END w_data_i[21]
  PIN w_data_i[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 117.635 0.07 117.705 ;
    END
  END w_data_i[220]
  PIN w_data_i[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 94.115 0.07 94.185 ;
    END
  END w_data_i[221]
  PIN w_data_i[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 28.875 94.11 28.945 ;
    END
  END w_data_i[222]
  PIN w_data_i[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 67.795 94.11 67.865 ;
    END
  END w_data_i[223]
  PIN w_data_i[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 8.715 94.11 8.785 ;
    END
  END w_data_i[224]
  PIN w_data_i[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.865 0 8.005 0.14 ;
    END
  END w_data_i[225]
  PIN w_data_i[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 118.755 94.11 118.825 ;
    END
  END w_data_i[226]
  PIN w_data_i[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  81.225 0 81.365 0.14 ;
    END
  END w_data_i[227]
  PIN w_data_i[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 6.475 0.07 6.545 ;
    END
  END w_data_i[228]
  PIN w_data_i[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  1.705 140.02 1.845 140.16 ;
    END
  END w_data_i[229]
  PIN w_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 34.475 0.07 34.545 ;
    END
  END w_data_i[22]
  PIN w_data_i[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 58.555 94.11 58.625 ;
    END
  END w_data_i[230]
  PIN w_data_i[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 115.395 94.11 115.465 ;
    END
  END w_data_i[231]
  PIN w_data_i[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 23.835 0.07 23.905 ;
    END
  END w_data_i[232]
  PIN w_data_i[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 122.955 0.07 123.025 ;
    END
  END w_data_i[233]
  PIN w_data_i[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 25.795 94.11 25.865 ;
    END
  END w_data_i[234]
  PIN w_data_i[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  75.625 0 75.765 0.14 ;
    END
  END w_data_i[235]
  PIN w_data_i[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 20.755 94.11 20.825 ;
    END
  END w_data_i[236]
  PIN w_data_i[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  2.265 0 2.405 0.14 ;
    END
  END w_data_i[237]
  PIN w_data_i[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  5.625 140.02 5.765 140.16 ;
    END
  END w_data_i[238]
  PIN w_data_i[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 110.355 94.11 110.425 ;
    END
  END w_data_i[239]
  PIN w_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 35.875 0.07 35.945 ;
    END
  END w_data_i[23]
  PIN w_data_i[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 80.675 0.07 80.745 ;
    END
  END w_data_i[240]
  PIN w_data_i[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 42.315 94.11 42.385 ;
    END
  END w_data_i[241]
  PIN w_data_i[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 84.315 0.07 84.385 ;
    END
  END w_data_i[242]
  PIN w_data_i[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 91.875 94.11 91.945 ;
    END
  END w_data_i[243]
  PIN w_data_i[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 99.995 0.07 100.065 ;
    END
  END w_data_i[244]
  PIN w_data_i[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 113.435 94.11 113.505 ;
    END
  END w_data_i[245]
  PIN w_data_i[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 129.675 0.07 129.745 ;
    END
  END w_data_i[246]
  PIN w_data_i[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 81.795 0.07 81.865 ;
    END
  END w_data_i[247]
  PIN w_data_i[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  76.745 0 76.885 0.14 ;
    END
  END w_data_i[248]
  PIN w_data_i[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 110.355 0.07 110.425 ;
    END
  END w_data_i[249]
  PIN w_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  40.345 0 40.485 0.14 ;
    END
  END w_data_i[24]
  PIN w_data_i[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  55.465 140.02 55.605 140.16 ;
    END
  END w_data_i[250]
  PIN w_data_i[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 68.075 0.07 68.145 ;
    END
  END w_data_i[251]
  PIN w_data_i[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  36.985 140.02 37.125 140.16 ;
    END
  END w_data_i[252]
  PIN w_data_i[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  87.945 140.02 88.085 140.16 ;
    END
  END w_data_i[253]
  PIN w_data_i[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 51.555 94.11 51.625 ;
    END
  END w_data_i[254]
  PIN w_data_i[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 2.275 0.07 2.345 ;
    END
  END w_data_i[255]
  PIN w_data_i[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  49.865 140.02 50.005 140.16 ;
    END
  END w_data_i[256]
  PIN w_data_i[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  29.145 140.02 29.285 140.16 ;
    END
  END w_data_i[257]
  PIN w_data_i[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  53.225 140.02 53.365 140.16 ;
    END
  END w_data_i[258]
  PIN w_data_i[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.675 0.07 31.745 ;
    END
  END w_data_i[259]
  PIN w_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 124.355 94.11 124.425 ;
    END
  END w_data_i[25]
  PIN w_data_i[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 111.195 0.07 111.265 ;
    END
  END w_data_i[260]
  PIN w_data_i[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 22.155 94.11 22.225 ;
    END
  END w_data_i[261]
  PIN w_data_i[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 16.275 0.07 16.345 ;
    END
  END w_data_i[262]
  PIN w_data_i[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 43.995 0.07 44.065 ;
    END
  END w_data_i[263]
  PIN w_data_i[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 109.235 94.11 109.305 ;
    END
  END w_data_i[264]
  PIN w_data_i[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  30.825 140.02 30.965 140.16 ;
    END
  END w_data_i[265]
  PIN w_data_i[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 125.195 0.07 125.265 ;
    END
  END w_data_i[266]
  PIN w_data_i[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 91.315 94.11 91.385 ;
    END
  END w_data_i[267]
  PIN w_data_i[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  21.865 140.02 22.005 140.16 ;
    END
  END w_data_i[268]
  PIN w_data_i[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 133.315 0.07 133.385 ;
    END
  END w_data_i[269]
  PIN w_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 71.715 0.07 71.785 ;
    END
  END w_data_i[26]
  PIN w_data_i[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 124.635 0.07 124.705 ;
    END
  END w_data_i[270]
  PIN w_data_i[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 14.035 94.11 14.105 ;
    END
  END w_data_i[271]
  PIN w_data_i[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 120.435 0.07 120.505 ;
    END
  END w_data_i[272]
  PIN w_data_i[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 64.155 0.07 64.225 ;
    END
  END w_data_i[273]
  PIN w_data_i[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 82.635 94.11 82.705 ;
    END
  END w_data_i[274]
  PIN w_data_i[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 28.875 0.07 28.945 ;
    END
  END w_data_i[275]
  PIN w_data_i[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 126.315 0.07 126.385 ;
    END
  END w_data_i[276]
  PIN w_data_i[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  56.025 140.02 56.165 140.16 ;
    END
  END w_data_i[277]
  PIN w_data_i[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  87.385 0 87.525 0.14 ;
    END
  END w_data_i[278]
  PIN w_data_i[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 119.315 94.11 119.385 ;
    END
  END w_data_i[279]
  PIN w_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 4.235 0.07 4.305 ;
    END
  END w_data_i[27]
  PIN w_data_i[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 87.955 0.07 88.025 ;
    END
  END w_data_i[280]
  PIN w_data_i[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 128.555 94.11 128.625 ;
    END
  END w_data_i[281]
  PIN w_data_i[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  22.425 140.02 22.565 140.16 ;
    END
  END w_data_i[282]
  PIN w_data_i[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 90.195 94.11 90.265 ;
    END
  END w_data_i[283]
  PIN w_data_i[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 138.075 0.07 138.145 ;
    END
  END w_data_i[284]
  PIN w_data_i[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 6.755 94.11 6.825 ;
    END
  END w_data_i[285]
  PIN w_data_i[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  57.705 0 57.845 0.14 ;
    END
  END w_data_i[286]
  PIN w_data_i[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  91.865 140.02 92.005 140.16 ;
    END
  END w_data_i[287]
  PIN w_data_i[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 72.555 0.07 72.625 ;
    END
  END w_data_i[288]
  PIN w_data_i[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 125.475 94.11 125.545 ;
    END
  END w_data_i[289]
  PIN w_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  70.025 0 70.165 0.14 ;
    END
  END w_data_i[28]
  PIN w_data_i[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  38.105 140.02 38.245 140.16 ;
    END
  END w_data_i[290]
  PIN w_data_i[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 20.755 0.07 20.825 ;
    END
  END w_data_i[291]
  PIN w_data_i[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 85.995 94.11 86.065 ;
    END
  END w_data_i[292]
  PIN w_data_i[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 52.675 94.11 52.745 ;
    END
  END w_data_i[293]
  PIN w_data_i[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 83.195 0.07 83.265 ;
    END
  END w_data_i[294]
  PIN w_data_i[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 130.795 94.11 130.865 ;
    END
  END w_data_i[295]
  PIN w_data_i[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 129.955 0.07 130.025 ;
    END
  END w_data_i[296]
  PIN w_data_i[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  89.065 0 89.205 0.14 ;
    END
  END w_data_i[297]
  PIN w_data_i[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  49.865 0 50.005 0.14 ;
    END
  END w_data_i[298]
  PIN w_data_i[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 119.875 94.11 119.945 ;
    END
  END w_data_i[299]
  PIN w_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 40.635 0.07 40.705 ;
    END
  END w_data_i[29]
  PIN w_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 12.355 94.11 12.425 ;
    END
  END w_data_i[2]
  PIN w_data_i[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  45.945 140.02 46.085 140.16 ;
    END
  END w_data_i[300]
  PIN w_data_i[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 86.275 94.11 86.345 ;
    END
  END w_data_i[301]
  PIN w_data_i[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 138.075 94.11 138.145 ;
    END
  END w_data_i[302]
  PIN w_data_i[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  8.985 0 9.125 0.14 ;
    END
  END w_data_i[303]
  PIN w_data_i[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 10.955 94.11 11.025 ;
    END
  END w_data_i[304]
  PIN w_data_i[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 130.235 94.11 130.305 ;
    END
  END w_data_i[305]
  PIN w_data_i[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 38.955 94.11 39.025 ;
    END
  END w_data_i[306]
  PIN w_data_i[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 107.835 94.11 107.905 ;
    END
  END w_data_i[307]
  PIN w_data_i[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 61.075 0.07 61.145 ;
    END
  END w_data_i[308]
  PIN w_data_i[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 33.075 0.07 33.145 ;
    END
  END w_data_i[309]
  PIN w_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 136.115 94.11 136.185 ;
    END
  END w_data_i[30]
  PIN w_data_i[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 2.835 94.11 2.905 ;
    END
  END w_data_i[310]
  PIN w_data_i[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 87.395 94.11 87.465 ;
    END
  END w_data_i[311]
  PIN w_data_i[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 38.395 94.11 38.465 ;
    END
  END w_data_i[312]
  PIN w_data_i[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 99.715 0.07 99.785 ;
    END
  END w_data_i[313]
  PIN w_data_i[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 3.395 0.07 3.465 ;
    END
  END w_data_i[314]
  PIN w_data_i[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  43.145 140.02 43.285 140.16 ;
    END
  END w_data_i[315]
  PIN w_data_i[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 50.995 0.07 51.065 ;
    END
  END w_data_i[316]
  PIN w_data_i[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  33.065 140.02 33.205 140.16 ;
    END
  END w_data_i[317]
  PIN w_data_i[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 95.795 94.11 95.865 ;
    END
  END w_data_i[318]
  PIN w_data_i[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 24.395 0.07 24.465 ;
    END
  END w_data_i[319]
  PIN w_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 95.795 0.07 95.865 ;
    END
  END w_data_i[31]
  PIN w_data_i[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 110.075 0.07 110.145 ;
    END
  END w_data_i[320]
  PIN w_data_i[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 5.355 0.07 5.425 ;
    END
  END w_data_i[321]
  PIN w_data_i[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 79.275 94.11 79.345 ;
    END
  END w_data_i[322]
  PIN w_data_i[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 52.115 94.11 52.185 ;
    END
  END w_data_i[323]
  PIN w_data_i[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  35.305 140.02 35.445 140.16 ;
    END
  END w_data_i[324]
  PIN w_data_i[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 50.715 0.07 50.785 ;
    END
  END w_data_i[325]
  PIN w_data_i[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 18.795 94.11 18.865 ;
    END
  END w_data_i[326]
  PIN w_data_i[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 85.995 0.07 86.065 ;
    END
  END w_data_i[327]
  PIN w_data_i[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 52.955 94.11 53.025 ;
    END
  END w_data_i[328]
  PIN w_data_i[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  54.905 140.02 55.045 140.16 ;
    END
  END w_data_i[329]
  PIN w_data_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  43.145 0 43.285 0.14 ;
    END
  END w_data_i[32]
  PIN w_data_i[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 134.715 94.11 134.785 ;
    END
  END w_data_i[330]
  PIN w_data_i[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 113.715 94.11 113.785 ;
    END
  END w_data_i[331]
  PIN w_data_i[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 91.315 0.07 91.385 ;
    END
  END w_data_i[332]
  PIN w_data_i[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 103.355 94.11 103.425 ;
    END
  END w_data_i[333]
  PIN w_data_i[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 104.755 0.07 104.825 ;
    END
  END w_data_i[334]
  PIN w_data_i[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 75.355 94.11 75.425 ;
    END
  END w_data_i[335]
  PIN w_data_i[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 35.035 0.07 35.105 ;
    END
  END w_data_i[336]
  PIN w_data_i[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 98.035 94.11 98.105 ;
    END
  END w_data_i[337]
  PIN w_data_i[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  78.985 0 79.125 0.14 ;
    END
  END w_data_i[338]
  PIN w_data_i[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 138.915 94.11 138.985 ;
    END
  END w_data_i[339]
  PIN w_data_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 19.075 94.11 19.145 ;
    END
  END w_data_i[33]
  PIN w_data_i[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 126.875 94.11 126.945 ;
    END
  END w_data_i[340]
  PIN w_data_i[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 83.475 0.07 83.545 ;
    END
  END w_data_i[341]
  PIN w_data_i[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 48.475 94.11 48.545 ;
    END
  END w_data_i[342]
  PIN w_data_i[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 30.275 94.11 30.345 ;
    END
  END w_data_i[343]
  PIN w_data_i[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.945 0 18.085 0.14 ;
    END
  END w_data_i[344]
  PIN w_data_i[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  28.025 0 28.165 0.14 ;
    END
  END w_data_i[345]
  PIN w_data_i[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 66.955 94.11 67.025 ;
    END
  END w_data_i[346]
  PIN w_data_i[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 58.275 0.07 58.345 ;
    END
  END w_data_i[347]
  PIN w_data_i[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 91.875 0.07 91.945 ;
    END
  END w_data_i[348]
  PIN w_data_i[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 121.835 94.11 121.905 ;
    END
  END w_data_i[349]
  PIN w_data_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 27.755 94.11 27.825 ;
    END
  END w_data_i[34]
  PIN w_data_i[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  20.185 0 20.325 0.14 ;
    END
  END w_data_i[350]
  PIN w_data_i[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 95.235 0.07 95.305 ;
    END
  END w_data_i[351]
  PIN w_data_i[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 32.795 94.11 32.865 ;
    END
  END w_data_i[352]
  PIN w_data_i[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  82.345 0 82.485 0.14 ;
    END
  END w_data_i[353]
  PIN w_data_i[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 26.075 0.07 26.145 ;
    END
  END w_data_i[354]
  PIN w_data_i[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 89.915 0.07 89.985 ;
    END
  END w_data_i[355]
  PIN w_data_i[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 92.155 94.11 92.225 ;
    END
  END w_data_i[356]
  PIN w_data_i[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 66.675 0.07 66.745 ;
    END
  END w_data_i[357]
  PIN w_data_i[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 24.395 94.11 24.465 ;
    END
  END w_data_i[358]
  PIN w_data_i[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 22.995 94.11 23.065 ;
    END
  END w_data_i[359]
  PIN w_data_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 102.235 0.07 102.305 ;
    END
  END w_data_i[35]
  PIN w_data_i[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 24.955 94.11 25.025 ;
    END
  END w_data_i[360]
  PIN w_data_i[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 99.155 0.07 99.225 ;
    END
  END w_data_i[361]
  PIN w_data_i[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  36.425 0 36.565 0.14 ;
    END
  END w_data_i[362]
  PIN w_data_i[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 56.315 94.11 56.385 ;
    END
  END w_data_i[363]
  PIN w_data_i[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 67.515 94.11 67.585 ;
    END
  END w_data_i[364]
  PIN w_data_i[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  68.345 140.02 68.485 140.16 ;
    END
  END w_data_i[365]
  PIN w_data_i[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 111.195 94.11 111.265 ;
    END
  END w_data_i[366]
  PIN w_data_i[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 84.875 0.07 84.945 ;
    END
  END w_data_i[367]
  PIN w_data_i[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 15.995 94.11 16.065 ;
    END
  END w_data_i[368]
  PIN w_data_i[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 45.395 94.11 45.465 ;
    END
  END w_data_i[369]
  PIN w_data_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 1.715 94.11 1.785 ;
    END
  END w_data_i[36]
  PIN w_data_i[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 103.915 0.07 103.985 ;
    END
  END w_data_i[370]
  PIN w_data_i[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 23.555 94.11 23.625 ;
    END
  END w_data_i[371]
  PIN w_data_i[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 50.155 94.11 50.225 ;
    END
  END w_data_i[372]
  PIN w_data_i[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 30.555 94.11 30.625 ;
    END
  END w_data_i[373]
  PIN w_data_i[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  68.345 0 68.485 0.14 ;
    END
  END w_data_i[374]
  PIN w_data_i[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  69.465 140.02 69.605 140.16 ;
    END
  END w_data_i[375]
  PIN w_data_i[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 17.675 94.11 17.745 ;
    END
  END w_data_i[376]
  PIN w_data_i[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 1.155 0.07 1.225 ;
    END
  END w_data_i[377]
  PIN w_data_i[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 59.115 0.07 59.185 ;
    END
  END w_data_i[378]
  PIN w_data_i[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 106.995 94.11 107.065 ;
    END
  END w_data_i[379]
  PIN w_data_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 100.275 94.11 100.345 ;
    END
  END w_data_i[37]
  PIN w_data_i[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 1.435 94.11 1.505 ;
    END
  END w_data_i[380]
  PIN w_data_i[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  3.945 0 4.085 0.14 ;
    END
  END w_data_i[381]
  PIN w_data_i[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 51.275 0.07 51.345 ;
    END
  END w_data_i[382]
  PIN w_data_i[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 50.435 0.07 50.505 ;
    END
  END w_data_i[383]
  PIN w_data_i[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 55.475 94.11 55.545 ;
    END
  END w_data_i[384]
  PIN w_data_i[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 78.995 0.07 79.065 ;
    END
  END w_data_i[385]
  PIN w_data_i[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 9.835 0.07 9.905 ;
    END
  END w_data_i[386]
  PIN w_data_i[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 70.035 0.07 70.105 ;
    END
  END w_data_i[387]
  PIN w_data_i[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 75.075 0.07 75.145 ;
    END
  END w_data_i[388]
  PIN w_data_i[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 10.675 0.07 10.745 ;
    END
  END w_data_i[389]
  PIN w_data_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 62.475 0.07 62.545 ;
    END
  END w_data_i[38]
  PIN w_data_i[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 16.835 0.07 16.905 ;
    END
  END w_data_i[390]
  PIN w_data_i[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 107.555 0.07 107.625 ;
    END
  END w_data_i[391]
  PIN w_data_i[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 42.595 0.07 42.665 ;
    END
  END w_data_i[392]
  PIN w_data_i[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 57.715 94.11 57.785 ;
    END
  END w_data_i[393]
  PIN w_data_i[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 34.195 0.07 34.265 ;
    END
  END w_data_i[394]
  PIN w_data_i[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  71.145 0 71.285 0.14 ;
    END
  END w_data_i[395]
  PIN w_data_i[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 135.275 0.07 135.345 ;
    END
  END w_data_i[396]
  PIN w_data_i[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 47.355 0.07 47.425 ;
    END
  END w_data_i[397]
  PIN w_data_i[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 112.035 94.11 112.105 ;
    END
  END w_data_i[398]
  PIN w_data_i[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 112.035 0.07 112.105 ;
    END
  END w_data_i[399]
  PIN w_data_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 8.435 0.07 8.505 ;
    END
  END w_data_i[39]
  PIN w_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 76.475 94.11 76.545 ;
    END
  END w_data_i[3]
  PIN w_data_i[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 8.995 94.11 9.065 ;
    END
  END w_data_i[400]
  PIN w_data_i[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 47.075 0.07 47.145 ;
    END
  END w_data_i[401]
  PIN w_data_i[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.315 0.07 7.385 ;
    END
  END w_data_i[402]
  PIN w_data_i[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 64.995 0.07 65.065 ;
    END
  END w_data_i[403]
  PIN w_data_i[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 113.435 0.07 113.505 ;
    END
  END w_data_i[404]
  PIN w_data_i[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  62.745 0 62.885 0.14 ;
    END
  END w_data_i[405]
  PIN w_data_i[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 13.755 0.07 13.825 ;
    END
  END w_data_i[406]
  PIN w_data_i[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 41.475 94.11 41.545 ;
    END
  END w_data_i[407]
  PIN w_data_i[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 131.355 0.07 131.425 ;
    END
  END w_data_i[408]
  PIN w_data_i[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 57.155 0.07 57.225 ;
    END
  END w_data_i[409]
  PIN w_data_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 94.675 0.07 94.745 ;
    END
  END w_data_i[40]
  PIN w_data_i[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 44.555 0.07 44.625 ;
    END
  END w_data_i[410]
  PIN w_data_i[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 2.275 94.11 2.345 ;
    END
  END w_data_i[411]
  PIN w_data_i[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  49.305 140.02 49.445 140.16 ;
    END
  END w_data_i[412]
  PIN w_data_i[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 40.635 94.11 40.705 ;
    END
  END w_data_i[413]
  PIN w_data_i[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 133.035 94.11 133.105 ;
    END
  END w_data_i[414]
  PIN w_data_i[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  45.945 0 46.085 0.14 ;
    END
  END w_data_i[415]
  PIN w_data_i[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 88.515 0.07 88.585 ;
    END
  END w_data_i[416]
  PIN w_data_i[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 22.715 94.11 22.785 ;
    END
  END w_data_i[417]
  PIN w_data_i[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 14.875 94.11 14.945 ;
    END
  END w_data_i[418]
  PIN w_data_i[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  9.545 140.02 9.685 140.16 ;
    END
  END w_data_i[419]
  PIN w_data_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 116.515 94.11 116.585 ;
    END
  END w_data_i[41]
  PIN w_data_i[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 77.595 94.11 77.665 ;
    END
  END w_data_i[420]
  PIN w_data_i[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 136.395 94.11 136.465 ;
    END
  END w_data_i[421]
  PIN w_data_i[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 29.155 94.11 29.225 ;
    END
  END w_data_i[422]
  PIN w_data_i[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 26.915 0.07 26.985 ;
    END
  END w_data_i[423]
  PIN w_data_i[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 52.955 0.07 53.025 ;
    END
  END w_data_i[424]
  PIN w_data_i[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  42.585 140.02 42.725 140.16 ;
    END
  END w_data_i[425]
  PIN w_data_i[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 108.395 94.11 108.465 ;
    END
  END w_data_i[426]
  PIN w_data_i[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 124.915 94.11 124.985 ;
    END
  END w_data_i[427]
  PIN w_data_i[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 49.595 94.11 49.665 ;
    END
  END w_data_i[428]
  PIN w_data_i[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 9.275 0.07 9.345 ;
    END
  END w_data_i[429]
  PIN w_data_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  76.185 140.02 76.325 140.16 ;
    END
  END w_data_i[42]
  PIN w_data_i[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 41.195 0.07 41.265 ;
    END
  END w_data_i[430]
  PIN w_data_i[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  19.065 0 19.205 0.14 ;
    END
  END w_data_i[431]
  PIN w_data_i[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 15.715 94.11 15.785 ;
    END
  END w_data_i[432]
  PIN w_data_i[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  66.105 0 66.245 0.14 ;
    END
  END w_data_i[433]
  PIN w_data_i[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 88.795 94.11 88.865 ;
    END
  END w_data_i[434]
  PIN w_data_i[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.595 0.07 7.665 ;
    END
  END w_data_i[435]
  PIN w_data_i[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 24.955 0.07 25.025 ;
    END
  END w_data_i[436]
  PIN w_data_i[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 85.435 94.11 85.505 ;
    END
  END w_data_i[437]
  PIN w_data_i[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  26.905 140.02 27.045 140.16 ;
    END
  END w_data_i[438]
  PIN w_data_i[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 115.115 94.11 115.185 ;
    END
  END w_data_i[439]
  PIN w_data_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  25.225 0 25.365 0.14 ;
    END
  END w_data_i[43]
  PIN w_data_i[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 106.435 94.11 106.505 ;
    END
  END w_data_i[440]
  PIN w_data_i[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 33.075 94.11 33.145 ;
    END
  END w_data_i[441]
  PIN w_data_i[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 132.755 0.07 132.825 ;
    END
  END w_data_i[442]
  PIN w_data_i[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 26.915 94.11 26.985 ;
    END
  END w_data_i[443]
  PIN w_data_i[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 127.995 94.11 128.065 ;
    END
  END w_data_i[444]
  PIN w_data_i[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  16.265 140.02 16.405 140.16 ;
    END
  END w_data_i[445]
  PIN w_data_i[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 134.715 0.07 134.785 ;
    END
  END w_data_i[446]
  PIN w_data_i[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 107.275 0.07 107.345 ;
    END
  END w_data_i[447]
  PIN w_data_i[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  19.625 140.02 19.765 140.16 ;
    END
  END w_data_i[448]
  PIN w_data_i[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 68.635 0.07 68.705 ;
    END
  END w_data_i[449]
  PIN w_data_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  74.505 0 74.645 0.14 ;
    END
  END w_data_i[44]
  PIN w_data_i[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 73.395 94.11 73.465 ;
    END
  END w_data_i[450]
  PIN w_data_i[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 101.675 94.11 101.745 ;
    END
  END w_data_i[451]
  PIN w_data_i[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 129.675 94.11 129.745 ;
    END
  END w_data_i[452]
  PIN w_data_i[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 17.395 0.07 17.465 ;
    END
  END w_data_i[453]
  PIN w_data_i[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 40.355 94.11 40.425 ;
    END
  END w_data_i[454]
  PIN w_data_i[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  63.865 140.02 64.005 140.16 ;
    END
  END w_data_i[455]
  PIN w_data_i[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  92.425 140.02 92.565 140.16 ;
    END
  END w_data_i[456]
  PIN w_data_i[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  5.065 140.02 5.205 140.16 ;
    END
  END w_data_i[457]
  PIN w_data_i[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 27.475 0.07 27.545 ;
    END
  END w_data_i[458]
  PIN w_data_i[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 56.595 94.11 56.665 ;
    END
  END w_data_i[459]
  PIN w_data_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  42.025 140.02 42.165 140.16 ;
    END
  END w_data_i[45]
  PIN w_data_i[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 52.395 94.11 52.465 ;
    END
  END w_data_i[460]
  PIN w_data_i[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 71.155 94.11 71.225 ;
    END
  END w_data_i[461]
  PIN w_data_i[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  39.785 0 39.925 0.14 ;
    END
  END w_data_i[462]
  PIN w_data_i[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  60.505 0 60.645 0.14 ;
    END
  END w_data_i[463]
  PIN w_data_i[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 58.835 94.11 58.905 ;
    END
  END w_data_i[464]
  PIN w_data_i[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 14.315 0.07 14.385 ;
    END
  END w_data_i[465]
  PIN w_data_i[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  67.785 140.02 67.925 140.16 ;
    END
  END w_data_i[466]
  PIN w_data_i[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 100.835 0.07 100.905 ;
    END
  END w_data_i[467]
  PIN w_data_i[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 96.635 0.07 96.705 ;
    END
  END w_data_i[468]
  PIN w_data_i[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 79.555 0.07 79.625 ;
    END
  END w_data_i[469]
  PIN w_data_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  73.945 0 74.085 0.14 ;
    END
  END w_data_i[46]
  PIN w_data_i[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  47.625 140.02 47.765 140.16 ;
    END
  END w_data_i[470]
  PIN w_data_i[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 68.635 94.11 68.705 ;
    END
  END w_data_i[471]
  PIN w_data_i[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 74.795 0.07 74.865 ;
    END
  END w_data_i[472]
  PIN w_data_i[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  47.625 0 47.765 0.14 ;
    END
  END w_data_i[473]
  PIN w_data_i[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  75.065 140.02 75.205 140.16 ;
    END
  END w_data_i[474]
  PIN w_data_i[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 123.515 0.07 123.585 ;
    END
  END w_data_i[475]
  PIN w_data_i[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 117.355 0.07 117.425 ;
    END
  END w_data_i[476]
  PIN w_data_i[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 136.675 0.07 136.745 ;
    END
  END w_data_i[477]
  PIN w_data_i[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  6.185 140.02 6.325 140.16 ;
    END
  END w_data_i[478]
  PIN w_data_i[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  8.425 140.02 8.565 140.16 ;
    END
  END w_data_i[479]
  PIN w_data_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 18.235 94.11 18.305 ;
    END
  END w_data_i[47]
  PIN w_data_i[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 107.835 0.07 107.905 ;
    END
  END w_data_i[480]
  PIN w_data_i[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 22.155 0.07 22.225 ;
    END
  END w_data_i[481]
  PIN w_data_i[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  3.385 0 3.525 0.14 ;
    END
  END w_data_i[482]
  PIN w_data_i[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 49.035 94.11 49.105 ;
    END
  END w_data_i[483]
  PIN w_data_i[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 18.515 94.11 18.585 ;
    END
  END w_data_i[484]
  PIN w_data_i[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 82.075 94.11 82.145 ;
    END
  END w_data_i[485]
  PIN w_data_i[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 120.155 0.07 120.225 ;
    END
  END w_data_i[486]
  PIN w_data_i[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 91.595 94.11 91.665 ;
    END
  END w_data_i[487]
  PIN w_data_i[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 50.155 0.07 50.225 ;
    END
  END w_data_i[488]
  PIN w_data_i[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.105 0 10.245 0.14 ;
    END
  END w_data_i[489]
  PIN w_data_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  48.185 0 48.325 0.14 ;
    END
  END w_data_i[48]
  PIN w_data_i[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 8.155 94.11 8.225 ;
    END
  END w_data_i[490]
  PIN w_data_i[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 108.955 0.07 109.025 ;
    END
  END w_data_i[491]
  PIN w_data_i[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 50.995 94.11 51.065 ;
    END
  END w_data_i[492]
  PIN w_data_i[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  92.425 0 92.565 0.14 ;
    END
  END w_data_i[493]
  PIN w_data_i[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 44.555 94.11 44.625 ;
    END
  END w_data_i[494]
  PIN w_data_i[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 40.915 0.07 40.985 ;
    END
  END w_data_i[495]
  PIN w_data_i[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  65.545 140.02 65.685 140.16 ;
    END
  END w_data_i[496]
  PIN w_data_i[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 46.515 94.11 46.585 ;
    END
  END w_data_i[497]
  PIN w_data_i[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 53.795 0.07 53.865 ;
    END
  END w_data_i[498]
  PIN w_data_i[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 71.435 94.11 71.505 ;
    END
  END w_data_i[499]
  PIN w_data_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  77.305 140.02 77.445 140.16 ;
    END
  END w_data_i[49]
  PIN w_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 97.755 0.07 97.825 ;
    END
  END w_data_i[4]
  PIN w_data_i[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 132.195 94.11 132.265 ;
    END
  END w_data_i[500]
  PIN w_data_i[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 43.995 94.11 44.065 ;
    END
  END w_data_i[501]
  PIN w_data_i[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 123.795 0.07 123.865 ;
    END
  END w_data_i[502]
  PIN w_data_i[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 82.915 94.11 82.985 ;
    END
  END w_data_i[503]
  PIN w_data_i[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 91.035 0.07 91.105 ;
    END
  END w_data_i[504]
  PIN w_data_i[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 62.195 94.11 62.265 ;
    END
  END w_data_i[505]
  PIN w_data_i[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 51.835 0.07 51.905 ;
    END
  END w_data_i[506]
  PIN w_data_i[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  30.265 0 30.405 0.14 ;
    END
  END w_data_i[507]
  PIN w_data_i[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 127.435 94.11 127.505 ;
    END
  END w_data_i[508]
  PIN w_data_i[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 19.635 94.11 19.705 ;
    END
  END w_data_i[509]
  PIN w_data_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  83.465 140.02 83.605 140.16 ;
    END
  END w_data_i[50]
  PIN w_data_i[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  58.825 0 58.965 0.14 ;
    END
  END w_data_i[510]
  PIN w_data_i[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 63.315 94.11 63.385 ;
    END
  END w_data_i[511]
  PIN w_data_i[512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 62.755 0.07 62.825 ;
    END
  END w_data_i[512]
  PIN w_data_i[513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 127.715 0.07 127.785 ;
    END
  END w_data_i[513]
  PIN w_data_i[514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  62.745 140.02 62.885 140.16 ;
    END
  END w_data_i[514]
  PIN w_data_i[515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 60.235 0.07 60.305 ;
    END
  END w_data_i[515]
  PIN w_data_i[516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 70.595 0.07 70.665 ;
    END
  END w_data_i[516]
  PIN w_data_i[517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 86.835 94.11 86.905 ;
    END
  END w_data_i[517]
  PIN w_data_i[518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 54.915 0.07 54.985 ;
    END
  END w_data_i[518]
  PIN w_data_i[519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 105.595 94.11 105.665 ;
    END
  END w_data_i[519]
  PIN w_data_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 109.795 0.07 109.865 ;
    END
  END w_data_i[51]
  PIN w_data_i[520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 86.835 0.07 86.905 ;
    END
  END w_data_i[520]
  PIN w_data_i[521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 43.715 0.07 43.785 ;
    END
  END w_data_i[521]
  PIN w_data_i[522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  21.305 0 21.445 0.14 ;
    END
  END w_data_i[522]
  PIN w_data_i[523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 16.555 94.11 16.625 ;
    END
  END w_data_i[523]
  PIN w_data_i[524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  78.985 140.02 79.125 140.16 ;
    END
  END w_data_i[524]
  PIN w_data_i[525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  92.985 140.02 93.125 140.16 ;
    END
  END w_data_i[525]
  PIN w_data_i[526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 17.955 0.07 18.025 ;
    END
  END w_data_i[526]
  PIN w_data_i[527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 130.515 94.11 130.585 ;
    END
  END w_data_i[527]
  PIN w_data_i[528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 98.875 94.11 98.945 ;
    END
  END w_data_i[528]
  PIN w_data_i[529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 60.235 94.11 60.305 ;
    END
  END w_data_i[529]
  PIN w_data_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 113.715 0.07 113.785 ;
    END
  END w_data_i[52]
  PIN w_data_i[530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.345 140.02 12.485 140.16 ;
    END
  END w_data_i[530]
  PIN w_data_i[531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 16.275 94.11 16.345 ;
    END
  END w_data_i[531]
  PIN w_data_i[532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 42.595 94.11 42.665 ;
    END
  END w_data_i[532]
  PIN w_data_i[533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 87.675 94.11 87.745 ;
    END
  END w_data_i[533]
  PIN w_data_i[534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 59.955 0.07 60.025 ;
    END
  END w_data_i[534]
  PIN w_data_i[535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 13.475 94.11 13.545 ;
    END
  END w_data_i[535]
  PIN w_data_i[536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  23.545 0 23.685 0.14 ;
    END
  END w_data_i[536]
  PIN w_data_i[537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 85.155 0.07 85.225 ;
    END
  END w_data_i[537]
  PIN w_data_i[538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 124.075 94.11 124.145 ;
    END
  END w_data_i[538]
  PIN w_data_i[539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  44.825 140.02 44.965 140.16 ;
    END
  END w_data_i[539]
  PIN w_data_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  84.025 0 84.165 0.14 ;
    END
  END w_data_i[53]
  PIN w_data_i[540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 135.835 0.07 135.905 ;
    END
  END w_data_i[540]
  PIN w_data_i[541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 105.875 94.11 105.945 ;
    END
  END w_data_i[541]
  PIN w_data_i[542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 37.275 94.11 37.345 ;
    END
  END w_data_i[542]
  PIN w_data_i[543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 134.435 0.07 134.505 ;
    END
  END w_data_i[543]
  PIN w_data_i[544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 33.915 94.11 33.985 ;
    END
  END w_data_i[544]
  PIN w_data_i[545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  67.785 0 67.925 0.14 ;
    END
  END w_data_i[545]
  PIN w_data_i[546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  11.225 0 11.365 0.14 ;
    END
  END w_data_i[546]
  PIN w_data_i[547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 59.675 94.11 59.745 ;
    END
  END w_data_i[547]
  PIN w_data_i[548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 87.955 94.11 88.025 ;
    END
  END w_data_i[548]
  PIN w_data_i[549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 90.475 0.07 90.545 ;
    END
  END w_data_i[549]
  PIN w_data_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  71.705 140.02 71.845 140.16 ;
    END
  END w_data_i[54]
  PIN w_data_i[550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 34.755 0.07 34.825 ;
    END
  END w_data_i[550]
  PIN w_data_i[551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 42.875 0.07 42.945 ;
    END
  END w_data_i[551]
  PIN w_data_i[552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 40.075 0.07 40.145 ;
    END
  END w_data_i[552]
  PIN w_data_i[553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  9.545 0 9.685 0.14 ;
    END
  END w_data_i[553]
  PIN w_data_i[554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  45.385 0 45.525 0.14 ;
    END
  END w_data_i[554]
  PIN w_data_i[555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 111.755 94.11 111.825 ;
    END
  END w_data_i[555]
  PIN w_data_i[556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 13.755 94.11 13.825 ;
    END
  END w_data_i[556]
  PIN w_data_i[557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 132.475 0.07 132.545 ;
    END
  END w_data_i[557]
  PIN w_data_i[558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  37.545 140.02 37.685 140.16 ;
    END
  END w_data_i[558]
  PIN w_data_i[559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 8.715 0.07 8.785 ;
    END
  END w_data_i[559]
  PIN w_data_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  32.505 0 32.645 0.14 ;
    END
  END w_data_i[55]
  PIN w_data_i[560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 118.195 94.11 118.265 ;
    END
  END w_data_i[560]
  PIN w_data_i[561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  46.505 140.02 46.645 140.16 ;
    END
  END w_data_i[561]
  PIN w_data_i[562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 15.715 0.07 15.785 ;
    END
  END w_data_i[562]
  PIN w_data_i[563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 135.555 94.11 135.625 ;
    END
  END w_data_i[563]
  PIN w_data_i[564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 89.075 94.11 89.145 ;
    END
  END w_data_i[564]
  PIN w_data_i[565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 24.675 94.11 24.745 ;
    END
  END w_data_i[565]
  PIN w_data_i[566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 14.035 0.07 14.105 ;
    END
  END w_data_i[566]
  PIN w_data_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 93.275 0.07 93.345 ;
    END
  END w_data_i[56]
  PIN w_data_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  63.865 0 64.005 0.14 ;
    END
  END w_data_i[57]
  PIN w_data_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 115.955 94.11 116.025 ;
    END
  END w_data_i[58]
  PIN w_data_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 36.715 94.11 36.785 ;
    END
  END w_data_i[59]
  PIN w_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 84.035 94.11 84.105 ;
    END
  END w_data_i[5]
  PIN w_data_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 24.675 0.07 24.745 ;
    END
  END w_data_i[60]
  PIN w_data_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 13.475 0.07 13.545 ;
    END
  END w_data_i[61]
  PIN w_data_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  33.625 0 33.765 0.14 ;
    END
  END w_data_i[62]
  PIN w_data_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 3.955 94.11 4.025 ;
    END
  END w_data_i[63]
  PIN w_data_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 96.915 94.11 96.985 ;
    END
  END w_data_i[64]
  PIN w_data_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  26.345 140.02 26.485 140.16 ;
    END
  END w_data_i[65]
  PIN w_data_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  88.505 140.02 88.645 140.16 ;
    END
  END w_data_i[66]
  PIN w_data_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 58.275 94.11 58.345 ;
    END
  END w_data_i[67]
  PIN w_data_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  16.265 0 16.405 0.14 ;
    END
  END w_data_i[68]
  PIN w_data_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 108.675 94.11 108.745 ;
    END
  END w_data_i[69]
  PIN w_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  5.065 0 5.205 0.14 ;
    END
  END w_data_i[6]
  PIN w_data_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  86.825 140.02 86.965 140.16 ;
    END
  END w_data_i[70]
  PIN w_data_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  23.545 140.02 23.685 140.16 ;
    END
  END w_data_i[71]
  PIN w_data_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 63.595 94.11 63.665 ;
    END
  END w_data_i[72]
  PIN w_data_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  19.065 140.02 19.205 140.16 ;
    END
  END w_data_i[73]
  PIN w_data_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 20.195 94.11 20.265 ;
    END
  END w_data_i[74]
  PIN w_data_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 13.195 0.07 13.265 ;
    END
  END w_data_i[75]
  PIN w_data_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 19.915 94.11 19.985 ;
    END
  END w_data_i[76]
  PIN w_data_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END w_data_i[77]
  PIN w_data_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 30.835 94.11 30.905 ;
    END
  END w_data_i[78]
  PIN w_data_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.395 0.07 31.465 ;
    END
  END w_data_i[79]
  PIN w_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 69.195 0.07 69.265 ;
    END
  END w_data_i[7]
  PIN w_data_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 109.235 0.07 109.305 ;
    END
  END w_data_i[80]
  PIN w_data_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 18.795 0.07 18.865 ;
    END
  END w_data_i[81]
  PIN w_data_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  41.465 0 41.605 0.14 ;
    END
  END w_data_i[82]
  PIN w_data_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  15.145 0 15.285 0.14 ;
    END
  END w_data_i[83]
  PIN w_data_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 134.155 0.07 134.225 ;
    END
  END w_data_i[84]
  PIN w_data_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 113.155 0.07 113.225 ;
    END
  END w_data_i[85]
  PIN w_data_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 6.195 94.11 6.265 ;
    END
  END w_data_i[86]
  PIN w_data_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  25.225 140.02 25.365 140.16 ;
    END
  END w_data_i[87]
  PIN w_data_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 75.915 94.11 75.985 ;
    END
  END w_data_i[88]
  PIN w_data_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 54.355 0.07 54.425 ;
    END
  END w_data_i[89]
  PIN w_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 122.115 94.11 122.185 ;
    END
  END w_data_i[8]
  PIN w_data_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  42.585 0 42.725 0.14 ;
    END
  END w_data_i[90]
  PIN w_data_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  72.825 0 72.965 0.14 ;
    END
  END w_data_i[91]
  PIN w_data_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 3.675 0.07 3.745 ;
    END
  END w_data_i[92]
  PIN w_data_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 117.915 94.11 117.985 ;
    END
  END w_data_i[93]
  PIN w_data_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 11.515 94.11 11.585 ;
    END
  END w_data_i[94]
  PIN w_data_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  24.665 140.02 24.805 140.16 ;
    END
  END w_data_i[95]
  PIN w_data_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  22.985 140.02 23.125 140.16 ;
    END
  END w_data_i[96]
  PIN w_data_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 83.755 0.07 83.825 ;
    END
  END w_data_i[97]
  PIN w_data_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 101.115 0.07 101.185 ;
    END
  END w_data_i[98]
  PIN w_data_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 21.875 94.11 21.945 ;
    END
  END w_data_i[99]
  PIN w_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 19.915 0.07 19.985 ;
    END
  END w_data_i[9]
  PIN w_reset_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 76.475 0.07 76.545 ;
    END
  END w_reset_i
  PIN w_v_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  94.04 92.715 94.11 92.785 ;
    END
  END w_v_i
  OBS
    LAYER metal1 ;
     RECT  0 -0.085 3.23 140.16 ;
     RECT  3.23 0 94.11 140.16 ;
    LAYER metal2 ;
     RECT  0 0 94.11 140.16 ;
    LAYER metal3 ;
     RECT  0 0 94.11 140.16 ;
    LAYER metal4 ;
     RECT  0 0 94.11 140.16 ;
  END
END bsg_mem_p567
END LIBRARY
