VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MACRO spram_12x4
  FOREIGN spram_12x4 0 0 ;
  CLASS BLOCK ;
  SIZE 12.69 BY 66.14 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 62.915 11.59 63.085 ;
        RECT  1.14 60.115 11.59 60.285 ;
        RECT  1.14 57.315 11.59 57.485 ;
        RECT  1.14 54.515 11.59 54.685 ;
        RECT  1.14 51.715 11.59 51.885 ;
        RECT  1.14 48.915 11.59 49.085 ;
        RECT  1.14 46.115 11.59 46.285 ;
        RECT  1.14 43.315 11.59 43.485 ;
        RECT  1.14 40.515 11.59 40.685 ;
        RECT  1.14 37.715 11.59 37.885 ;
        RECT  1.14 34.915 11.59 35.085 ;
        RECT  1.14 32.115 11.59 32.285 ;
        RECT  1.14 29.315 11.59 29.485 ;
        RECT  1.14 26.515 11.59 26.685 ;
        RECT  1.14 23.715 11.59 23.885 ;
        RECT  1.14 20.915 11.59 21.085 ;
        RECT  1.14 18.115 11.59 18.285 ;
        RECT  1.14 15.315 11.59 15.485 ;
        RECT  1.14 12.515 11.59 12.685 ;
        RECT  1.14 9.715 11.59 9.885 ;
        RECT  1.14 6.915 11.59 7.085 ;
        RECT  1.14 4.115 11.59 4.285 ;
        RECT  1.14 1.315 11.59 1.485 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 64.315 11.59 64.485 ;
        RECT  1.14 61.515 11.59 61.685 ;
        RECT  1.14 58.715 11.59 58.885 ;
        RECT  1.14 55.915 11.59 56.085 ;
        RECT  1.14 53.115 11.59 53.285 ;
        RECT  1.14 50.315 11.59 50.485 ;
        RECT  1.14 47.515 11.59 47.685 ;
        RECT  1.14 44.715 11.59 44.885 ;
        RECT  1.14 41.915 11.59 42.085 ;
        RECT  1.14 39.115 11.59 39.285 ;
        RECT  1.14 36.315 11.59 36.485 ;
        RECT  1.14 33.515 11.59 33.685 ;
        RECT  1.14 30.715 11.59 30.885 ;
        RECT  1.14 27.915 11.59 28.085 ;
        RECT  1.14 25.115 11.59 25.285 ;
        RECT  1.14 22.315 11.59 22.485 ;
        RECT  1.14 19.515 11.59 19.685 ;
        RECT  1.14 16.715 11.59 16.885 ;
        RECT  1.14 13.915 11.59 14.085 ;
        RECT  1.14 11.115 11.59 11.285 ;
        RECT  1.14 8.315 11.59 8.485 ;
        RECT  1.14 5.515 11.59 5.685 ;
        RECT  1.14 2.715 11.59 2.885 ;
    END
  END VDD
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 44.835 0.07 44.905 ;
    END
  END clk
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 64.995 0.07 65.065 ;
    END
  END din[0]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 36.995 0.07 37.065 ;
    END
  END din[1]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 28.875 0.07 28.945 ;
    END
  END din[2]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  12.62 22.995 12.69 23.065 ;
    END
  END din[3]
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.915 0.07 12.985 ;
    END
  END dout[0]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 61.075 0.07 61.145 ;
    END
  END dout[1]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 4.795 0.07 4.865 ;
    END
  END dout[2]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 20.755 0.07 20.825 ;
    END
  END dout[3]
  PIN raddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  12.62 55.195 12.69 55.265 ;
    END
  END raddr[0]
  PIN raddr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  12.62 31.115 12.69 31.185 ;
    END
  END raddr[10]
  PIN raddr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  12.62 26.915 12.69 26.985 ;
    END
  END raddr[11]
  PIN raddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 8.715 0.07 8.785 ;
    END
  END raddr[1]
  PIN raddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  12.62 50.995 12.69 51.065 ;
    END
  END raddr[2]
  PIN raddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END raddr[3]
  PIN raddr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 56.875 0.07 56.945 ;
    END
  END raddr[4]
  PIN raddr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  12.62 43.155 12.69 43.225 ;
    END
  END raddr[5]
  PIN raddr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 24.955 0.07 25.025 ;
    END
  END raddr[6]
  PIN raddr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 40.915 0.07 40.985 ;
    END
  END raddr[7]
  PIN raddr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  12.62 19.075 12.69 19.145 ;
    END
  END raddr[8]
  PIN raddr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.865 66 8.005 66.14 ;
    END
  END raddr[9]
  PIN re
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  12.62 35.035 12.69 35.105 ;
    END
  END re
  PIN waddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  8.425 0 8.565 0.14 ;
    END
  END waddr[0]
  PIN waddr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  12.62 2.835 12.69 2.905 ;
    END
  END waddr[10]
  PIN waddr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  12.62 7.035 12.69 7.105 ;
    END
  END waddr[11]
  PIN waddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  12.62 38.955 12.69 39.025 ;
    END
  END waddr[1]
  PIN waddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  12.62 10.955 12.69 11.025 ;
    END
  END waddr[2]
  PIN waddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  12.62 59.115 12.69 59.185 ;
    END
  END waddr[3]
  PIN waddr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  12.62 63.035 12.69 63.105 ;
    END
  END waddr[4]
  PIN waddr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 49.035 0.07 49.105 ;
    END
  END waddr[5]
  PIN waddr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 52.955 0.07 53.025 ;
    END
  END waddr[6]
  PIN waddr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  12.62 14.875 12.69 14.945 ;
    END
  END waddr[7]
  PIN waddr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 16.835 0.07 16.905 ;
    END
  END waddr[8]
  PIN waddr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 32.795 0.07 32.865 ;
    END
  END waddr[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  12.62 47.075 12.69 47.145 ;
    END
  END we
  OBS
    LAYER metal1 ;
     RECT  0 -0.085 3.23 66.14 ;
     RECT  3.23 0 12.69 66.14 ;
    LAYER metal2 ;
     RECT  0 0 12.69 66.14 ;
    LAYER metal3 ;
     RECT  0 0 12.69 66.14 ;
    LAYER metal4 ;
     RECT  0 0 12.69 66.14 ;
  END
END spram_12x4
END LIBRARY
