VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MACRO fifo_v3_8
  FOREIGN fifo_v3_8 0 0 ;
  CLASS BLOCK ;
  SIZE 123.245 BY 147.49 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 144.115 122.17 144.285 ;
        RECT  1.14 141.315 122.17 141.485 ;
        RECT  1.14 138.515 122.17 138.685 ;
        RECT  1.14 135.715 122.17 135.885 ;
        RECT  1.14 132.915 122.17 133.085 ;
        RECT  1.14 130.115 122.17 130.285 ;
        RECT  1.14 127.315 122.17 127.485 ;
        RECT  1.14 124.515 122.17 124.685 ;
        RECT  1.14 121.715 122.17 121.885 ;
        RECT  1.14 118.915 122.17 119.085 ;
        RECT  1.14 116.115 122.17 116.285 ;
        RECT  1.14 113.315 122.17 113.485 ;
        RECT  1.14 110.515 122.17 110.685 ;
        RECT  1.14 107.715 122.17 107.885 ;
        RECT  1.14 104.915 122.17 105.085 ;
        RECT  1.14 102.115 122.17 102.285 ;
        RECT  1.14 99.315 122.17 99.485 ;
        RECT  1.14 96.515 122.17 96.685 ;
        RECT  1.14 93.715 122.17 93.885 ;
        RECT  1.14 90.915 122.17 91.085 ;
        RECT  1.14 88.115 122.17 88.285 ;
        RECT  1.14 85.315 122.17 85.485 ;
        RECT  1.14 82.515 122.17 82.685 ;
        RECT  1.14 79.715 122.17 79.885 ;
        RECT  1.14 76.915 122.17 77.085 ;
        RECT  1.14 74.115 122.17 74.285 ;
        RECT  1.14 71.315 122.17 71.485 ;
        RECT  1.14 68.515 122.17 68.685 ;
        RECT  1.14 65.715 122.17 65.885 ;
        RECT  1.14 62.915 122.17 63.085 ;
        RECT  1.14 60.115 122.17 60.285 ;
        RECT  1.14 57.315 122.17 57.485 ;
        RECT  1.14 54.515 122.17 54.685 ;
        RECT  1.14 51.715 122.17 51.885 ;
        RECT  1.14 48.915 122.17 49.085 ;
        RECT  1.14 46.115 122.17 46.285 ;
        RECT  1.14 43.315 122.17 43.485 ;
        RECT  1.14 40.515 122.17 40.685 ;
        RECT  1.14 37.715 122.17 37.885 ;
        RECT  1.14 34.915 122.17 35.085 ;
        RECT  1.14 32.115 122.17 32.285 ;
        RECT  1.14 29.315 122.17 29.485 ;
        RECT  1.14 26.515 122.17 26.685 ;
        RECT  1.14 23.715 122.17 23.885 ;
        RECT  1.14 20.915 122.17 21.085 ;
        RECT  1.14 18.115 122.17 18.285 ;
        RECT  1.14 15.315 122.17 15.485 ;
        RECT  1.14 12.515 122.17 12.685 ;
        RECT  1.14 9.715 122.17 9.885 ;
        RECT  1.14 6.915 122.17 7.085 ;
        RECT  1.14 4.115 122.17 4.285 ;
        RECT  1.14 1.315 122.17 1.485 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 145.515 122.17 145.685 ;
        RECT  1.14 142.715 122.17 142.885 ;
        RECT  1.14 139.915 122.17 140.085 ;
        RECT  1.14 137.115 122.17 137.285 ;
        RECT  1.14 134.315 122.17 134.485 ;
        RECT  1.14 131.515 122.17 131.685 ;
        RECT  1.14 128.715 122.17 128.885 ;
        RECT  1.14 125.915 122.17 126.085 ;
        RECT  1.14 123.115 122.17 123.285 ;
        RECT  1.14 120.315 122.17 120.485 ;
        RECT  1.14 117.515 122.17 117.685 ;
        RECT  1.14 114.715 122.17 114.885 ;
        RECT  1.14 111.915 122.17 112.085 ;
        RECT  1.14 109.115 122.17 109.285 ;
        RECT  1.14 106.315 122.17 106.485 ;
        RECT  1.14 103.515 122.17 103.685 ;
        RECT  1.14 100.715 122.17 100.885 ;
        RECT  1.14 97.915 122.17 98.085 ;
        RECT  1.14 95.115 122.17 95.285 ;
        RECT  1.14 92.315 122.17 92.485 ;
        RECT  1.14 89.515 122.17 89.685 ;
        RECT  1.14 86.715 122.17 86.885 ;
        RECT  1.14 83.915 122.17 84.085 ;
        RECT  1.14 81.115 122.17 81.285 ;
        RECT  1.14 78.315 122.17 78.485 ;
        RECT  1.14 75.515 122.17 75.685 ;
        RECT  1.14 72.715 122.17 72.885 ;
        RECT  1.14 69.915 122.17 70.085 ;
        RECT  1.14 67.115 122.17 67.285 ;
        RECT  1.14 64.315 122.17 64.485 ;
        RECT  1.14 61.515 122.17 61.685 ;
        RECT  1.14 58.715 122.17 58.885 ;
        RECT  1.14 55.915 122.17 56.085 ;
        RECT  1.14 53.115 122.17 53.285 ;
        RECT  1.14 50.315 122.17 50.485 ;
        RECT  1.14 47.515 122.17 47.685 ;
        RECT  1.14 44.715 122.17 44.885 ;
        RECT  1.14 41.915 122.17 42.085 ;
        RECT  1.14 39.115 122.17 39.285 ;
        RECT  1.14 36.315 122.17 36.485 ;
        RECT  1.14 33.515 122.17 33.685 ;
        RECT  1.14 30.715 122.17 30.885 ;
        RECT  1.14 27.915 122.17 28.085 ;
        RECT  1.14 25.115 122.17 25.285 ;
        RECT  1.14 22.315 122.17 22.485 ;
        RECT  1.14 19.515 122.17 19.685 ;
        RECT  1.14 16.715 122.17 16.885 ;
        RECT  1.14 13.915 122.17 14.085 ;
        RECT  1.14 11.115 122.17 11.285 ;
        RECT  1.14 8.315 122.17 8.485 ;
        RECT  1.14 5.515 122.17 5.685 ;
        RECT  1.14 2.715 122.17 2.885 ;
    END
  END VDD
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 38.115 123.245 38.185 ;
    END
  END clk_i
  PIN data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 87.115 123.245 87.185 ;
    END
  END data_i[0]
  PIN data_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 58.555 123.245 58.625 ;
    END
  END data_i[100]
  PIN data_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 87.115 0.07 87.185 ;
    END
  END data_i[101]
  PIN data_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  75.625 147.35 75.765 147.49 ;
    END
  END data_i[102]
  PIN data_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.875 0.07 7.945 ;
    END
  END data_i[103]
  PIN data_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 61.915 123.245 61.985 ;
    END
  END data_i[104]
  PIN data_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  61.065 147.35 61.205 147.49 ;
    END
  END data_i[105]
  PIN data_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 45.115 123.245 45.185 ;
    END
  END data_i[106]
  PIN data_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 133.875 0.07 133.945 ;
    END
  END data_i[107]
  PIN data_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 6.755 0.07 6.825 ;
    END
  END data_i[108]
  PIN data_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 12.915 123.245 12.985 ;
    END
  END data_i[109]
  PIN data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 131.355 0.07 131.425 ;
    END
  END data_i[10]
  PIN data_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  74.505 0 74.645 0.14 ;
    END
  END data_i[110]
  PIN data_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 41.755 123.245 41.825 ;
    END
  END data_i[111]
  PIN data_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 89.635 123.245 89.705 ;
    END
  END data_i[112]
  PIN data_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  113.145 0 113.285 0.14 ;
    END
  END data_i[113]
  PIN data_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 75.355 123.245 75.425 ;
    END
  END data_i[114]
  PIN data_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  104.185 147.35 104.325 147.49 ;
    END
  END data_i[115]
  PIN data_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 67.795 0.07 67.865 ;
    END
  END data_i[116]
  PIN data_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  15.705 147.35 15.845 147.49 ;
    END
  END data_i[117]
  PIN data_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 84.595 0.07 84.665 ;
    END
  END data_i[118]
  PIN data_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 3.395 123.245 3.465 ;
    END
  END data_i[119]
  PIN data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 111.195 123.245 111.265 ;
    END
  END data_i[11]
  PIN data_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 45.115 0.07 45.185 ;
    END
  END data_i[120]
  PIN data_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 70.315 0.07 70.385 ;
    END
  END data_i[121]
  PIN data_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 64.435 123.245 64.505 ;
    END
  END data_i[122]
  PIN data_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  98.585 0 98.725 0.14 ;
    END
  END data_i[123]
  PIN data_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 75.075 0.07 75.145 ;
    END
  END data_i[124]
  PIN data_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  109.225 147.35 109.365 147.49 ;
    END
  END data_i[125]
  PIN data_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  55.465 0 55.605 0.14 ;
    END
  END data_i[126]
  PIN data_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 76.195 0.07 76.265 ;
    END
  END data_i[127]
  PIN data_i[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 81.235 123.245 81.305 ;
    END
  END data_i[128]
  PIN data_i[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 105.315 123.245 105.385 ;
    END
  END data_i[129]
  PIN data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 66.955 123.245 67.025 ;
    END
  END data_i[12]
  PIN data_i[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  91.305 0 91.445 0.14 ;
    END
  END data_i[130]
  PIN data_i[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 105.035 0.07 105.105 ;
    END
  END data_i[131]
  PIN data_i[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 56.035 0.07 56.105 ;
    END
  END data_i[132]
  PIN data_i[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 31.955 123.245 32.025 ;
    END
  END data_i[133]
  PIN data_i[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 17.395 0.07 17.465 ;
    END
  END data_i[134]
  PIN data_i[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.345 0 12.485 0.14 ;
    END
  END data_i[135]
  PIN data_i[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 58.275 0.07 58.345 ;
    END
  END data_i[136]
  PIN data_i[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 114.555 0.07 114.625 ;
    END
  END data_i[137]
  PIN data_i[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  42.025 147.35 42.165 147.49 ;
    END
  END data_i[138]
  PIN data_i[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  20.185 147.35 20.325 147.49 ;
    END
  END data_i[139]
  PIN data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 119.595 123.245 119.665 ;
    END
  END data_i[13]
  PIN data_i[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 18.795 0.07 18.865 ;
    END
  END data_i[140]
  PIN data_i[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  56.585 147.35 56.725 147.49 ;
    END
  END data_i[141]
  PIN data_i[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 61.915 0.07 61.985 ;
    END
  END data_i[142]
  PIN data_i[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 19.915 0.07 19.985 ;
    END
  END data_i[143]
  PIN data_i[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 21.315 123.245 21.385 ;
    END
  END data_i[144]
  PIN data_i[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  120.425 0 120.565 0.14 ;
    END
  END data_i[145]
  PIN data_i[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  70.585 147.35 70.725 147.49 ;
    END
  END data_i[146]
  PIN data_i[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 122.955 0.07 123.025 ;
    END
  END data_i[147]
  PIN data_i[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  58.825 147.35 58.965 147.49 ;
    END
  END data_i[148]
  PIN data_i[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  114.265 147.35 114.405 147.49 ;
    END
  END data_i[149]
  PIN data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  111.465 147.35 111.605 147.49 ;
    END
  END data_i[14]
  PIN data_i[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 102.795 0.07 102.865 ;
    END
  END data_i[150]
  PIN data_i[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  106.985 147.35 107.125 147.49 ;
    END
  END data_i[151]
  PIN data_i[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 52.395 0.07 52.465 ;
    END
  END data_i[152]
  PIN data_i[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 24.675 0.07 24.745 ;
    END
  END data_i[153]
  PIN data_i[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  103.625 0 103.765 0.14 ;
    END
  END data_i[154]
  PIN data_i[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 137.515 123.245 137.585 ;
    END
  END data_i[155]
  PIN data_i[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 114.835 123.245 114.905 ;
    END
  END data_i[156]
  PIN data_i[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 121.835 0.07 121.905 ;
    END
  END data_i[157]
  PIN data_i[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 126.595 0.07 126.665 ;
    END
  END data_i[158]
  PIN data_i[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 115.955 123.245 116.025 ;
    END
  END data_i[159]
  PIN data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 112.315 123.245 112.385 ;
    END
  END data_i[15]
  PIN data_i[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  60.505 0 60.645 0.14 ;
    END
  END data_i[160]
  PIN data_i[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  67.225 0 67.365 0.14 ;
    END
  END data_i[161]
  PIN data_i[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  117.625 0 117.765 0.14 ;
    END
  END data_i[162]
  PIN data_i[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 88.235 0.07 88.305 ;
    END
  END data_i[163]
  PIN data_i[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 127.995 123.245 128.065 ;
    END
  END data_i[164]
  PIN data_i[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 109.795 0.07 109.865 ;
    END
  END data_i[165]
  PIN data_i[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 65.555 0.07 65.625 ;
    END
  END data_i[166]
  PIN data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 63.315 123.245 63.385 ;
    END
  END data_i[16]
  PIN data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 26.075 123.245 26.145 ;
    END
  END data_i[17]
  PIN data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 48.755 0.07 48.825 ;
    END
  END data_i[18]
  PIN data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 120.715 123.245 120.785 ;
    END
  END data_i[19]
  PIN data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 49.875 0.07 49.945 ;
    END
  END data_i[1]
  PIN data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 145.915 123.245 145.985 ;
    END
  END data_i[20]
  PIN data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  118.745 147.35 118.885 147.49 ;
    END
  END data_i[21]
  PIN data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 59.395 0.07 59.465 ;
    END
  END data_i[22]
  PIN data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  1.145 147.35 1.285 147.49 ;
    END
  END data_i[23]
  PIN data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  84.025 0 84.165 0.14 ;
    END
  END data_i[24]
  PIN data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  92.425 147.35 92.565 147.49 ;
    END
  END data_i[25]
  PIN data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 118.195 0.07 118.265 ;
    END
  END data_i[26]
  PIN data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 144.795 0.07 144.865 ;
    END
  END data_i[27]
  PIN data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 51.275 123.245 51.345 ;
    END
  END data_i[28]
  PIN data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  64.985 0 65.125 0.14 ;
    END
  END data_i[29]
  PIN data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  68.345 147.35 68.485 147.49 ;
    END
  END data_i[2]
  PIN data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  99.705 147.35 99.845 147.49 ;
    END
  END data_i[30]
  PIN data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 124.355 123.245 124.425 ;
    END
  END data_i[31]
  PIN data_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 34.195 0.07 34.265 ;
    END
  END data_i[32]
  PIN data_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 8.995 0.07 9.065 ;
    END
  END data_i[33]
  PIN data_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  30.265 147.35 30.405 147.49 ;
    END
  END data_i[34]
  PIN data_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  53.225 0 53.365 0.14 ;
    END
  END data_i[35]
  PIN data_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 142.275 0.07 142.345 ;
    END
  END data_i[36]
  PIN data_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 141.155 0.07 141.225 ;
    END
  END data_i[37]
  PIN data_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 77.595 0.07 77.665 ;
    END
  END data_i[38]
  PIN data_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 81.235 0.07 81.305 ;
    END
  END data_i[39]
  PIN data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 117.075 0.07 117.145 ;
    END
  END data_i[3]
  PIN data_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 50.155 123.245 50.225 ;
    END
  END data_i[40]
  PIN data_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 42.595 0.07 42.665 ;
    END
  END data_i[41]
  PIN data_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 40.355 123.245 40.425 ;
    END
  END data_i[42]
  PIN data_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  82.905 147.35 83.045 147.49 ;
    END
  END data_i[43]
  PIN data_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 37.835 0.07 37.905 ;
    END
  END data_i[44]
  PIN data_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 99.155 0.07 99.225 ;
    END
  END data_i[45]
  PIN data_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 56.035 123.245 56.105 ;
    END
  END data_i[46]
  PIN data_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 138.635 0.07 138.705 ;
    END
  END data_i[47]
  PIN data_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 29.435 0.07 29.505 ;
    END
  END data_i[48]
  PIN data_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  57.705 0 57.845 0.14 ;
    END
  END data_i[49]
  PIN data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 47.635 123.245 47.705 ;
    END
  END data_i[4]
  PIN data_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 14.035 0.07 14.105 ;
    END
  END data_i[50]
  PIN data_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 106.155 0.07 106.225 ;
    END
  END data_i[51]
  PIN data_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  29.145 0 29.285 0.14 ;
    END
  END data_i[52]
  PIN data_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  6.185 147.35 6.325 147.49 ;
    END
  END data_i[53]
  PIN data_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.745 147.35 34.885 147.49 ;
    END
  END data_i[54]
  PIN data_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 54.915 123.245 54.985 ;
    END
  END data_i[55]
  PIN data_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 28.595 123.245 28.665 ;
    END
  END data_i[56]
  PIN data_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 73.955 123.245 74.025 ;
    END
  END data_i[57]
  PIN data_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 113.435 0.07 113.505 ;
    END
  END data_i[58]
  PIN data_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 136.395 123.245 136.465 ;
    END
  END data_i[59]
  PIN data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 42.875 123.245 42.945 ;
    END
  END data_i[5]
  PIN data_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  86.825 0 86.965 0.14 ;
    END
  END data_i[60]
  PIN data_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 29.715 123.245 29.785 ;
    END
  END data_i[61]
  PIN data_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  21.865 0 22.005 0.14 ;
    END
  END data_i[62]
  PIN data_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 83.755 123.245 83.825 ;
    END
  END data_i[63]
  PIN data_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 113.715 123.245 113.785 ;
    END
  END data_i[64]
  PIN data_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 90.755 0.07 90.825 ;
    END
  END data_i[65]
  PIN data_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 57.155 123.245 57.225 ;
    END
  END data_i[66]
  PIN data_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 24.955 123.245 25.025 ;
    END
  END data_i[67]
  PIN data_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 4.515 123.245 4.585 ;
    END
  END data_i[68]
  PIN data_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  49.305 147.35 49.445 147.49 ;
    END
  END data_i[69]
  PIN data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 15.155 0.07 15.225 ;
    END
  END data_i[6]
  PIN data_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 78.715 0.07 78.785 ;
    END
  END data_i[70]
  PIN data_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 88.515 123.245 88.585 ;
    END
  END data_i[71]
  PIN data_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 40.355 0.07 40.425 ;
    END
  END data_i[72]
  PIN data_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 23.555 123.245 23.625 ;
    END
  END data_i[73]
  PIN data_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 138.915 123.245 138.985 ;
    END
  END data_i[74]
  PIN data_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  105.865 0 106.005 0.14 ;
    END
  END data_i[75]
  PIN data_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 124.355 0.07 124.425 ;
    END
  END data_i[76]
  PIN data_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 48.755 123.245 48.825 ;
    END
  END data_i[77]
  PIN data_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 93.275 123.245 93.345 ;
    END
  END data_i[78]
  PIN data_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 89.635 0.07 89.705 ;
    END
  END data_i[79]
  PIN data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  70.025 0 70.165 0.14 ;
    END
  END data_i[7]
  PIN data_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  36.985 147.35 37.125 147.49 ;
    END
  END data_i[80]
  PIN data_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 17.675 123.245 17.745 ;
    END
  END data_i[81]
  PIN data_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  39.785 147.35 39.925 147.49 ;
    END
  END data_i[82]
  PIN data_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  38.665 0 38.805 0.14 ;
    END
  END data_i[83]
  PIN data_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 83.475 0.07 83.545 ;
    END
  END data_i[84]
  PIN data_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 125.475 0.07 125.545 ;
    END
  END data_i[85]
  PIN data_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 34.475 123.245 34.545 ;
    END
  END data_i[86]
  PIN data_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 25.795 0.07 25.865 ;
    END
  END data_i[87]
  PIN data_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 134.995 0.07 135.065 ;
    END
  END data_i[88]
  PIN data_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.035 0.07 21.105 ;
    END
  END data_i[89]
  PIN data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 50.995 0.07 51.065 ;
    END
  END data_i[8]
  PIN data_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  89.065 0 89.205 0.14 ;
    END
  END data_i[90]
  PIN data_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 47.635 0.07 47.705 ;
    END
  END data_i[91]
  PIN data_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 73.955 0.07 74.025 ;
    END
  END data_i[92]
  PIN data_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  87.385 147.35 87.525 147.49 ;
    END
  END data_i[93]
  PIN data_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 103.915 123.245 103.985 ;
    END
  END data_i[94]
  PIN data_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 111.195 0.07 111.265 ;
    END
  END data_i[95]
  PIN data_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 92.995 0.07 93.065 ;
    END
  END data_i[96]
  PIN data_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 16.275 0.07 16.345 ;
    END
  END data_i[97]
  PIN data_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 15.155 123.245 15.225 ;
    END
  END data_i[98]
  PIN data_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 82.355 0.07 82.425 ;
    END
  END data_i[99]
  PIN data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 127.995 0.07 128.065 ;
    END
  END data_i[9]
  PIN data_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 66.675 0.07 66.745 ;
    END
  END data_o[0]
  PIN data_o[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 108.675 0.07 108.745 ;
    END
  END data_o[100]
  PIN data_o[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 57.155 0.07 57.225 ;
    END
  END data_o[101]
  PIN data_o[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 60.795 123.245 60.865 ;
    END
  END data_o[102]
  PIN data_o[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 90.755 123.245 90.825 ;
    END
  END data_o[103]
  PIN data_o[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 77.595 123.245 77.665 ;
    END
  END data_o[104]
  PIN data_o[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 6.755 123.245 6.825 ;
    END
  END data_o[105]
  PIN data_o[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 95.515 0.07 95.585 ;
    END
  END data_o[106]
  PIN data_o[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 5.635 123.245 5.705 ;
    END
  END data_o[107]
  PIN data_o[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 107.555 0.07 107.625 ;
    END
  END data_o[108]
  PIN data_o[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  26.905 0 27.045 0.14 ;
    END
  END data_o[109]
  PIN data_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  40.905 0 41.045 0.14 ;
    END
  END data_o[10]
  PIN data_o[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 10.395 0.07 10.465 ;
    END
  END data_o[110]
  PIN data_o[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 36.995 123.245 37.065 ;
    END
  END data_o[111]
  PIN data_o[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 76.475 123.245 76.545 ;
    END
  END data_o[112]
  PIN data_o[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 126.875 123.245 126.945 ;
    END
  END data_o[113]
  PIN data_o[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 130.515 123.245 130.585 ;
    END
  END data_o[114]
  PIN data_o[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 143.675 123.245 143.745 ;
    END
  END data_o[115]
  PIN data_o[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  50.425 0 50.565 0.14 ;
    END
  END data_o[116]
  PIN data_o[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 85.995 123.245 86.065 ;
    END
  END data_o[117]
  PIN data_o[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 33.075 0.07 33.145 ;
    END
  END data_o[118]
  PIN data_o[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  116.505 147.35 116.645 147.49 ;
    END
  END data_o[119]
  PIN data_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 53.515 0.07 53.585 ;
    END
  END data_o[11]
  PIN data_o[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  22.985 147.35 23.125 147.49 ;
    END
  END data_o[120]
  PIN data_o[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 117.355 123.245 117.425 ;
    END
  END data_o[121]
  PIN data_o[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 123.235 123.245 123.305 ;
    END
  END data_o[122]
  PIN data_o[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 110.075 123.245 110.145 ;
    END
  END data_o[123]
  PIN data_o[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  66.105 147.35 66.245 147.49 ;
    END
  END data_o[124]
  PIN data_o[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 106.435 123.245 106.505 ;
    END
  END data_o[125]
  PIN data_o[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  94.105 0 94.245 0.14 ;
    END
  END data_o[126]
  PIN data_o[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 134.155 123.245 134.225 ;
    END
  END data_o[127]
  PIN data_o[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 43.995 0.07 44.065 ;
    END
  END data_o[128]
  PIN data_o[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  2.825 0 2.965 0.14 ;
    END
  END data_o[129]
  PIN data_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 129.115 0.07 129.185 ;
    END
  END data_o[12]
  PIN data_o[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  96.345 0 96.485 0.14 ;
    END
  END data_o[130]
  PIN data_o[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 35.595 123.245 35.665 ;
    END
  END data_o[131]
  PIN data_o[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 129.115 123.245 129.185 ;
    END
  END data_o[132]
  PIN data_o[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 145.915 0.07 145.985 ;
    END
  END data_o[133]
  PIN data_o[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  47.065 147.35 47.205 147.49 ;
    END
  END data_o[134]
  PIN data_o[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 79.835 0.07 79.905 ;
    END
  END data_o[135]
  PIN data_o[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  36.425 0 36.565 0.14 ;
    END
  END data_o[136]
  PIN data_o[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  81.785 0 81.925 0.14 ;
    END
  END data_o[137]
  PIN data_o[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 142.555 123.245 142.625 ;
    END
  END data_o[138]
  PIN data_o[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 91.875 0.07 91.945 ;
    END
  END data_o[139]
  PIN data_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  72.265 0 72.405 0.14 ;
    END
  END data_o[13]
  PIN data_o[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 10.395 123.245 10.465 ;
    END
  END data_o[140]
  PIN data_o[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 78.715 123.245 78.785 ;
    END
  END data_o[141]
  PIN data_o[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 96.915 123.245 96.985 ;
    END
  END data_o[142]
  PIN data_o[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 3.115 0.07 3.185 ;
    END
  END data_o[143]
  PIN data_o[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  32.505 147.35 32.645 147.49 ;
    END
  END data_o[144]
  PIN data_o[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 112.315 0.07 112.385 ;
    END
  END data_o[145]
  PIN data_o[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 1.995 0.07 2.065 ;
    END
  END data_o[146]
  PIN data_o[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  97.465 147.35 97.605 147.49 ;
    END
  END data_o[147]
  PIN data_o[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 139.755 0.07 139.825 ;
    END
  END data_o[148]
  PIN data_o[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 11.795 123.245 11.865 ;
    END
  END data_o[149]
  PIN data_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 140.035 123.245 140.105 ;
    END
  END data_o[14]
  PIN data_o[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.955 0.07 32.025 ;
    END
  END data_o[150]
  PIN data_o[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 41.475 0.07 41.545 ;
    END
  END data_o[151]
  PIN data_o[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 27.195 123.245 27.265 ;
    END
  END data_o[152]
  PIN data_o[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.665 147.35 10.805 147.49 ;
    END
  END data_o[153]
  PIN data_o[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  24.105 0 24.245 0.14 ;
    END
  END data_o[154]
  PIN data_o[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 82.355 123.245 82.425 ;
    END
  END data_o[155]
  PIN data_o[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 119.595 0.07 119.665 ;
    END
  END data_o[156]
  PIN data_o[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 98.035 123.245 98.105 ;
    END
  END data_o[157]
  PIN data_o[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  48.185 0 48.325 0.14 ;
    END
  END data_o[158]
  PIN data_o[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 30.835 123.245 30.905 ;
    END
  END data_o[159]
  PIN data_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.945 147.35 18.085 147.49 ;
    END
  END data_o[15]
  PIN data_o[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 69.195 0.07 69.265 ;
    END
  END data_o[160]
  PIN data_o[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 108.955 123.245 109.025 ;
    END
  END data_o[161]
  PIN data_o[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  8.425 147.35 8.565 147.49 ;
    END
  END data_o[162]
  PIN data_o[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  25.225 147.35 25.365 147.49 ;
    END
  END data_o[163]
  PIN data_o[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 52.395 123.245 52.465 ;
    END
  END data_o[164]
  PIN data_o[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 143.395 0.07 143.465 ;
    END
  END data_o[165]
  PIN data_o[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 69.195 123.245 69.265 ;
    END
  END data_o[166]
  PIN data_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  85.145 147.35 85.285 147.49 ;
    END
  END data_o[16]
  PIN data_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  44.265 147.35 44.405 147.49 ;
    END
  END data_o[17]
  PIN data_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 130.235 0.07 130.305 ;
    END
  END data_o[18]
  PIN data_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 46.235 0.07 46.305 ;
    END
  END data_o[19]
  PIN data_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 103.915 0.07 103.985 ;
    END
  END data_o[1]
  PIN data_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 107.555 123.245 107.625 ;
    END
  END data_o[20]
  PIN data_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 102.795 123.245 102.865 ;
    END
  END data_o[21]
  PIN data_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 0.875 123.245 0.945 ;
    END
  END data_o[22]
  PIN data_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 100.275 0.07 100.345 ;
    END
  END data_o[23]
  PIN data_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 68.075 123.245 68.145 ;
    END
  END data_o[24]
  PIN data_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 33.355 123.245 33.425 ;
    END
  END data_o[25]
  PIN data_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  77.865 147.35 78.005 147.49 ;
    END
  END data_o[26]
  PIN data_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 141.155 123.245 141.225 ;
    END
  END data_o[27]
  PIN data_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 22.435 0.07 22.505 ;
    END
  END data_o[28]
  PIN data_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 18.795 123.245 18.865 ;
    END
  END data_o[29]
  PIN data_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 59.675 123.245 59.745 ;
    END
  END data_o[2]
  PIN data_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 132.755 0.07 132.825 ;
    END
  END data_o[30]
  PIN data_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  108.105 0 108.245 0.14 ;
    END
  END data_o[31]
  PIN data_o[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  19.625 0 19.765 0.14 ;
    END
  END data_o[32]
  PIN data_o[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  13.465 147.35 13.605 147.49 ;
    END
  END data_o[33]
  PIN data_o[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 95.515 123.245 95.585 ;
    END
  END data_o[34]
  PIN data_o[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 132.755 123.245 132.825 ;
    END
  END data_o[35]
  PIN data_o[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  77.305 0 77.445 0.14 ;
    END
  END data_o[36]
  PIN data_o[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 63.035 0.07 63.105 ;
    END
  END data_o[37]
  PIN data_o[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 80.115 123.245 80.185 ;
    END
  END data_o[38]
  PIN data_o[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 16.555 123.245 16.625 ;
    END
  END data_o[39]
  PIN data_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  94.665 147.35 94.805 147.49 ;
    END
  END data_o[3]
  PIN data_o[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 5.635 0.07 5.705 ;
    END
  END data_o[40]
  PIN data_o[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 60.795 0.07 60.865 ;
    END
  END data_o[41]
  PIN data_o[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.105 0 10.245 0.14 ;
    END
  END data_o[42]
  PIN data_o[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 39.235 123.245 39.305 ;
    END
  END data_o[43]
  PIN data_o[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 65.555 123.245 65.625 ;
    END
  END data_o[44]
  PIN data_o[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  3.385 147.35 3.525 147.49 ;
    END
  END data_o[45]
  PIN data_o[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 125.755 123.245 125.825 ;
    END
  END data_o[46]
  PIN data_o[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 30.835 0.07 30.905 ;
    END
  END data_o[47]
  PIN data_o[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 101.395 0.07 101.465 ;
    END
  END data_o[48]
  PIN data_o[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 98.035 0.07 98.105 ;
    END
  END data_o[49]
  PIN data_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.305 0 7.445 0.14 ;
    END
  END data_o[4]
  PIN data_o[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 27.195 0.07 27.265 ;
    END
  END data_o[50]
  PIN data_o[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 92.155 123.245 92.225 ;
    END
  END data_o[51]
  PIN data_o[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  115.385 0 115.525 0.14 ;
    END
  END data_o[52]
  PIN data_o[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 36.715 0.07 36.785 ;
    END
  END data_o[53]
  PIN data_o[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  120.985 147.35 121.125 147.49 ;
    END
  END data_o[54]
  PIN data_o[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 120.715 0.07 120.785 ;
    END
  END data_o[55]
  PIN data_o[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.385 0 31.525 0.14 ;
    END
  END data_o[56]
  PIN data_o[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 100.555 123.245 100.625 ;
    END
  END data_o[57]
  PIN data_o[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 144.795 123.245 144.865 ;
    END
  END data_o[58]
  PIN data_o[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 72.835 0.07 72.905 ;
    END
  END data_o[59]
  PIN data_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.635 0.07 12.705 ;
    END
  END data_o[5]
  PIN data_o[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 72.835 123.245 72.905 ;
    END
  END data_o[60]
  PIN data_o[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 9.275 123.245 9.345 ;
    END
  END data_o[61]
  PIN data_o[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  101.945 147.35 102.085 147.49 ;
    END
  END data_o[62]
  PIN data_o[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 4.235 0.07 4.305 ;
    END
  END data_o[63]
  PIN data_o[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  62.745 0 62.885 0.14 ;
    END
  END data_o[64]
  PIN data_o[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 101.675 123.245 101.745 ;
    END
  END data_o[65]
  PIN data_o[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 22.435 123.245 22.505 ;
    END
  END data_o[66]
  PIN data_o[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 70.315 123.245 70.385 ;
    END
  END data_o[67]
  PIN data_o[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 64.435 0.07 64.505 ;
    END
  END data_o[68]
  PIN data_o[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 43.995 123.245 44.065 ;
    END
  END data_o[69]
  PIN data_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  33.625 0 33.765 0.14 ;
    END
  END data_o[6]
  PIN data_o[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  100.825 0 100.965 0.14 ;
    END
  END data_o[70]
  PIN data_o[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 84.875 123.245 84.945 ;
    END
  END data_o[71]
  PIN data_o[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  90.185 147.35 90.325 147.49 ;
    END
  END data_o[72]
  PIN data_o[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 131.635 123.245 131.705 ;
    END
  END data_o[73]
  PIN data_o[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 46.515 123.245 46.585 ;
    END
  END data_o[74]
  PIN data_o[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  16.825 0 16.965 0.14 ;
    END
  END data_o[75]
  PIN data_o[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 99.155 123.245 99.225 ;
    END
  END data_o[76]
  PIN data_o[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  5.065 0 5.205 0.14 ;
    END
  END data_o[77]
  PIN data_o[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 135.275 123.245 135.345 ;
    END
  END data_o[78]
  PIN data_o[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  80.665 147.35 80.805 147.49 ;
    END
  END data_o[79]
  PIN data_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 53.515 123.245 53.585 ;
    END
  END data_o[7]
  PIN data_o[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  73.385 147.35 73.525 147.49 ;
    END
  END data_o[80]
  PIN data_o[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 35.595 0.07 35.665 ;
    END
  END data_o[81]
  PIN data_o[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 28.315 0.07 28.385 ;
    END
  END data_o[82]
  PIN data_o[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 8.155 123.245 8.225 ;
    END
  END data_o[83]
  PIN data_o[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END data_o[84]
  PIN data_o[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 20.195 123.245 20.265 ;
    END
  END data_o[85]
  PIN data_o[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 54.635 0.07 54.705 ;
    END
  END data_o[86]
  PIN data_o[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 94.395 0.07 94.465 ;
    END
  END data_o[87]
  PIN data_o[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 136.395 0.07 136.465 ;
    END
  END data_o[88]
  PIN data_o[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 39.235 0.07 39.305 ;
    END
  END data_o[89]
  PIN data_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  43.705 0 43.845 0.14 ;
    END
  END data_o[8]
  PIN data_o[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.585 0 14.725 0.14 ;
    END
  END data_o[90]
  PIN data_o[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  27.465 147.35 27.605 147.49 ;
    END
  END data_o[91]
  PIN data_o[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 137.515 0.07 137.585 ;
    END
  END data_o[92]
  PIN data_o[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  110.905 0 111.045 0.14 ;
    END
  END data_o[93]
  PIN data_o[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  63.865 147.35 64.005 147.49 ;
    END
  END data_o[94]
  PIN data_o[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 71.715 123.245 71.785 ;
    END
  END data_o[95]
  PIN data_o[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 71.435 0.07 71.505 ;
    END
  END data_o[96]
  PIN data_o[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 122.115 123.245 122.185 ;
    END
  END data_o[97]
  PIN data_o[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  45.945 0 46.085 0.14 ;
    END
  END data_o[98]
  PIN data_o[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  79.545 0 79.685 0.14 ;
    END
  END data_o[99]
  PIN data_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 11.515 0.07 11.585 ;
    END
  END data_o[9]
  PIN empty_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 118.475 123.245 118.545 ;
    END
  END empty_o
  PIN flush_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 1.995 123.245 2.065 ;
    END
  END flush_i
  PIN full_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  53.785 147.35 53.925 147.49 ;
    END
  END full_o
  PIN pop_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  51.545 147.35 51.685 147.49 ;
    END
  END pop_i
  PIN push_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 96.635 0.07 96.705 ;
    END
  END push_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 115.955 0.07 116.025 ;
    END
  END rst_ni
  PIN testmode_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 14.035 123.245 14.105 ;
    END
  END testmode_i
  PIN usage_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 23.555 0.07 23.625 ;
    END
  END usage_o[0]
  PIN usage_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 85.995 0.07 86.065 ;
    END
  END usage_o[1]
  PIN usage_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  123.175 94.395 123.245 94.465 ;
    END
  END usage_o[2]
  OBS
    LAYER metal1 ;
     RECT  0 -0.085 3.8 147.49 ;
     RECT  3.8 0 123.245 147.49 ;
    LAYER metal2 ;
     RECT  0 0 123.245 147.49 ;
    LAYER metal3 ;
     RECT  0 0 123.245 147.49 ;
    LAYER metal4 ;
     RECT  0 0 123.245 147.49 ;
  END
END fifo_v3_8
END LIBRARY
