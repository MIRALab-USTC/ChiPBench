VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MACRO memory_block_64x8
  FOREIGN memory_block_64x8 0 0 ;
  CLASS BLOCK ;
  SIZE 43.585 BY 126.755 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 124.515 42.56 124.685 ;
        RECT  1.14 121.715 42.56 121.885 ;
        RECT  1.14 118.915 42.56 119.085 ;
        RECT  1.14 116.115 42.56 116.285 ;
        RECT  1.14 113.315 42.56 113.485 ;
        RECT  1.14 110.515 42.56 110.685 ;
        RECT  1.14 107.715 42.56 107.885 ;
        RECT  1.14 104.915 42.56 105.085 ;
        RECT  1.14 102.115 42.56 102.285 ;
        RECT  1.14 99.315 42.56 99.485 ;
        RECT  1.14 96.515 42.56 96.685 ;
        RECT  1.14 93.715 42.56 93.885 ;
        RECT  1.14 90.915 42.56 91.085 ;
        RECT  1.14 88.115 42.56 88.285 ;
        RECT  1.14 85.315 42.56 85.485 ;
        RECT  1.14 82.515 42.56 82.685 ;
        RECT  1.14 79.715 42.56 79.885 ;
        RECT  1.14 76.915 42.56 77.085 ;
        RECT  1.14 74.115 42.56 74.285 ;
        RECT  1.14 71.315 42.56 71.485 ;
        RECT  1.14 68.515 42.56 68.685 ;
        RECT  1.14 65.715 42.56 65.885 ;
        RECT  1.14 62.915 42.56 63.085 ;
        RECT  1.14 60.115 42.56 60.285 ;
        RECT  1.14 57.315 42.56 57.485 ;
        RECT  1.14 54.515 42.56 54.685 ;
        RECT  1.14 51.715 42.56 51.885 ;
        RECT  1.14 48.915 42.56 49.085 ;
        RECT  1.14 46.115 42.56 46.285 ;
        RECT  1.14 43.315 42.56 43.485 ;
        RECT  1.14 40.515 42.56 40.685 ;
        RECT  1.14 37.715 42.56 37.885 ;
        RECT  1.14 34.915 42.56 35.085 ;
        RECT  1.14 32.115 42.56 32.285 ;
        RECT  1.14 29.315 42.56 29.485 ;
        RECT  1.14 26.515 42.56 26.685 ;
        RECT  1.14 23.715 42.56 23.885 ;
        RECT  1.14 20.915 42.56 21.085 ;
        RECT  1.14 18.115 42.56 18.285 ;
        RECT  1.14 15.315 42.56 15.485 ;
        RECT  1.14 12.515 42.56 12.685 ;
        RECT  1.14 9.715 42.56 9.885 ;
        RECT  1.14 6.915 42.56 7.085 ;
        RECT  1.14 4.115 42.56 4.285 ;
        RECT  1.14 1.315 42.56 1.485 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 123.115 42.56 123.285 ;
        RECT  1.14 120.315 42.56 120.485 ;
        RECT  1.14 117.515 42.56 117.685 ;
        RECT  1.14 114.715 42.56 114.885 ;
        RECT  1.14 111.915 42.56 112.085 ;
        RECT  1.14 109.115 42.56 109.285 ;
        RECT  1.14 106.315 42.56 106.485 ;
        RECT  1.14 103.515 42.56 103.685 ;
        RECT  1.14 100.715 42.56 100.885 ;
        RECT  1.14 97.915 42.56 98.085 ;
        RECT  1.14 95.115 42.56 95.285 ;
        RECT  1.14 92.315 42.56 92.485 ;
        RECT  1.14 89.515 42.56 89.685 ;
        RECT  1.14 86.715 42.56 86.885 ;
        RECT  1.14 83.915 42.56 84.085 ;
        RECT  1.14 81.115 42.56 81.285 ;
        RECT  1.14 78.315 42.56 78.485 ;
        RECT  1.14 75.515 42.56 75.685 ;
        RECT  1.14 72.715 42.56 72.885 ;
        RECT  1.14 69.915 42.56 70.085 ;
        RECT  1.14 67.115 42.56 67.285 ;
        RECT  1.14 64.315 42.56 64.485 ;
        RECT  1.14 61.515 42.56 61.685 ;
        RECT  1.14 58.715 42.56 58.885 ;
        RECT  1.14 55.915 42.56 56.085 ;
        RECT  1.14 53.115 42.56 53.285 ;
        RECT  1.14 50.315 42.56 50.485 ;
        RECT  1.14 47.515 42.56 47.685 ;
        RECT  1.14 44.715 42.56 44.885 ;
        RECT  1.14 41.915 42.56 42.085 ;
        RECT  1.14 39.115 42.56 39.285 ;
        RECT  1.14 36.315 42.56 36.485 ;
        RECT  1.14 33.515 42.56 33.685 ;
        RECT  1.14 30.715 42.56 30.885 ;
        RECT  1.14 27.915 42.56 28.085 ;
        RECT  1.14 25.115 42.56 25.285 ;
        RECT  1.14 22.315 42.56 22.485 ;
        RECT  1.14 19.515 42.56 19.685 ;
        RECT  1.14 16.715 42.56 16.885 ;
        RECT  1.14 13.915 42.56 14.085 ;
        RECT  1.14 11.115 42.56 11.285 ;
        RECT  1.14 8.315 42.56 8.485 ;
        RECT  1.14 5.515 42.56 5.685 ;
        RECT  1.14 2.715 42.56 2.885 ;
    END
  END VDD
  PIN di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 92.715 0.07 92.785 ;
    END
  END di[0]
  PIN di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.945 126.615 18.085 126.755 ;
    END
  END di[1]
  PIN di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 75.915 0.07 75.985 ;
    END
  END di[2]
  PIN di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 59.395 0.07 59.465 ;
    END
  END di[3]
  PIN di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.515 38.115 43.585 38.185 ;
    END
  END di[4]
  PIN di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 25.795 0.07 25.865 ;
    END
  END di[5]
  PIN di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  1.145 126.615 1.285 126.755 ;
    END
  END di[6]
  PIN di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 8.995 0.07 9.065 ;
    END
  END di[7]
  PIN do_slice[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 42.595 0.07 42.665 ;
    END
  END do_slice[0]
  PIN do_slice[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.515 105.035 43.585 105.105 ;
    END
  END do_slice[1]
  PIN do_slice[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.515 54.635 43.585 54.705 ;
    END
  END do_slice[2]
  PIN do_slice[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.515 46.515 43.585 46.585 ;
    END
  END do_slice[3]
  PIN do_slice[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 17.395 0.07 17.465 ;
    END
  END do_slice[4]
  PIN do_slice[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.515 96.635 43.585 96.705 ;
    END
  END do_slice[5]
  PIN do_slice[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END do_slice[6]
  PIN do_slice[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 117.915 0.07 117.985 ;
    END
  END do_slice[7]
  PIN raddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.515 79.835 43.585 79.905 ;
    END
  END raddr[0]
  PIN raddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 50.995 0.07 51.065 ;
    END
  END raddr[1]
  PIN raddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 84.315 0.07 84.385 ;
    END
  END raddr[2]
  PIN raddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.515 29.715 43.585 29.785 ;
    END
  END raddr[3]
  PIN raddr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.745 126.615 34.885 126.755 ;
    END
  END raddr[4]
  PIN raddr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.515 63.035 43.585 63.105 ;
    END
  END raddr[5]
  PIN rce
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  16.825 0 16.965 0.14 ;
    END
  END rce
  PIN rclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  33.625 0 33.765 0.14 ;
    END
  END rclk
  PIN rrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.515 4.515 43.585 4.585 ;
    END
  END rrst
  PIN waddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.515 71.435 43.585 71.505 ;
    END
  END waddr[0]
  PIN waddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.515 12.915 43.585 12.985 ;
    END
  END waddr[1]
  PIN waddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.515 113.435 43.585 113.505 ;
    END
  END waddr[2]
  PIN waddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.515 121.835 43.585 121.905 ;
    END
  END waddr[3]
  PIN waddr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 101.115 0.07 101.185 ;
    END
  END waddr[4]
  PIN waddr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 109.515 0.07 109.585 ;
    END
  END waddr[5]
  PIN wce
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.515 21.315 43.585 21.385 ;
    END
  END wce
  PIN wclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 34.195 0.07 34.265 ;
    END
  END wclk
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 67.795 0.07 67.865 ;
    END
  END we
  PIN wrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.515 88.235 43.585 88.305 ;
    END
  END wrst
  OBS
    LAYER metal1 ;
     RECT  0 -0.085 3.42 126.755 ;
     RECT  3.42 0 43.585 126.755 ;
    LAYER metal2 ;
     RECT  0 0 43.585 126.755 ;
    LAYER metal3 ;
     RECT  0 0 43.585 126.755 ;
    LAYER metal4 ;
     RECT  0 0 43.585 126.755 ;
  END
END memory_block_64x8
END LIBRARY
