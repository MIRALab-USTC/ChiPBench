VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MACRO small_mem_block
  FOREIGN small_mem_block 0 0 ;
  CLASS BLOCK ;
  SIZE 210.39 BY 418.78 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 417.115 209.38 417.285 ;
        RECT  1.14 414.315 209.38 414.485 ;
        RECT  1.14 411.515 209.38 411.685 ;
        RECT  1.14 408.715 209.38 408.885 ;
        RECT  1.14 405.915 209.38 406.085 ;
        RECT  1.14 403.115 209.38 403.285 ;
        RECT  1.14 400.315 209.38 400.485 ;
        RECT  1.14 397.515 209.38 397.685 ;
        RECT  1.14 394.715 209.38 394.885 ;
        RECT  1.14 391.915 209.38 392.085 ;
        RECT  1.14 389.115 209.38 389.285 ;
        RECT  1.14 386.315 209.38 386.485 ;
        RECT  1.14 383.515 209.38 383.685 ;
        RECT  1.14 380.715 209.38 380.885 ;
        RECT  1.14 377.915 209.38 378.085 ;
        RECT  1.14 375.115 209.38 375.285 ;
        RECT  1.14 372.315 209.38 372.485 ;
        RECT  1.14 369.515 209.38 369.685 ;
        RECT  1.14 366.715 209.38 366.885 ;
        RECT  1.14 363.915 209.38 364.085 ;
        RECT  1.14 361.115 209.38 361.285 ;
        RECT  1.14 358.315 209.38 358.485 ;
        RECT  1.14 355.515 209.38 355.685 ;
        RECT  1.14 352.715 209.38 352.885 ;
        RECT  1.14 349.915 209.38 350.085 ;
        RECT  1.14 347.115 209.38 347.285 ;
        RECT  1.14 344.315 209.38 344.485 ;
        RECT  1.14 341.515 209.38 341.685 ;
        RECT  1.14 338.715 209.38 338.885 ;
        RECT  1.14 335.915 209.38 336.085 ;
        RECT  1.14 333.115 209.38 333.285 ;
        RECT  1.14 330.315 209.38 330.485 ;
        RECT  1.14 327.515 209.38 327.685 ;
        RECT  1.14 324.715 209.38 324.885 ;
        RECT  1.14 321.915 209.38 322.085 ;
        RECT  1.14 319.115 209.38 319.285 ;
        RECT  1.14 316.315 209.38 316.485 ;
        RECT  1.14 313.515 209.38 313.685 ;
        RECT  1.14 310.715 209.38 310.885 ;
        RECT  1.14 307.915 209.38 308.085 ;
        RECT  1.14 305.115 209.38 305.285 ;
        RECT  1.14 302.315 209.38 302.485 ;
        RECT  1.14 299.515 209.38 299.685 ;
        RECT  1.14 296.715 209.38 296.885 ;
        RECT  1.14 293.915 209.38 294.085 ;
        RECT  1.14 291.115 209.38 291.285 ;
        RECT  1.14 288.315 209.38 288.485 ;
        RECT  1.14 285.515 209.38 285.685 ;
        RECT  1.14 282.715 209.38 282.885 ;
        RECT  1.14 279.915 209.38 280.085 ;
        RECT  1.14 277.115 209.38 277.285 ;
        RECT  1.14 274.315 209.38 274.485 ;
        RECT  1.14 271.515 209.38 271.685 ;
        RECT  1.14 268.715 209.38 268.885 ;
        RECT  1.14 265.915 209.38 266.085 ;
        RECT  1.14 263.115 209.38 263.285 ;
        RECT  1.14 260.315 209.38 260.485 ;
        RECT  1.14 257.515 209.38 257.685 ;
        RECT  1.14 254.715 209.38 254.885 ;
        RECT  1.14 251.915 209.38 252.085 ;
        RECT  1.14 249.115 209.38 249.285 ;
        RECT  1.14 246.315 209.38 246.485 ;
        RECT  1.14 243.515 209.38 243.685 ;
        RECT  1.14 240.715 209.38 240.885 ;
        RECT  1.14 237.915 209.38 238.085 ;
        RECT  1.14 235.115 209.38 235.285 ;
        RECT  1.14 232.315 209.38 232.485 ;
        RECT  1.14 229.515 209.38 229.685 ;
        RECT  1.14 226.715 209.38 226.885 ;
        RECT  1.14 223.915 209.38 224.085 ;
        RECT  1.14 221.115 209.38 221.285 ;
        RECT  1.14 218.315 209.38 218.485 ;
        RECT  1.14 215.515 209.38 215.685 ;
        RECT  1.14 212.715 209.38 212.885 ;
        RECT  1.14 209.915 209.38 210.085 ;
        RECT  1.14 207.115 209.38 207.285 ;
        RECT  1.14 204.315 209.38 204.485 ;
        RECT  1.14 201.515 209.38 201.685 ;
        RECT  1.14 198.715 209.38 198.885 ;
        RECT  1.14 195.915 209.38 196.085 ;
        RECT  1.14 193.115 209.38 193.285 ;
        RECT  1.14 190.315 209.38 190.485 ;
        RECT  1.14 187.515 209.38 187.685 ;
        RECT  1.14 184.715 209.38 184.885 ;
        RECT  1.14 181.915 209.38 182.085 ;
        RECT  1.14 179.115 209.38 179.285 ;
        RECT  1.14 176.315 209.38 176.485 ;
        RECT  1.14 173.515 209.38 173.685 ;
        RECT  1.14 170.715 209.38 170.885 ;
        RECT  1.14 167.915 209.38 168.085 ;
        RECT  1.14 165.115 209.38 165.285 ;
        RECT  1.14 162.315 209.38 162.485 ;
        RECT  1.14 159.515 209.38 159.685 ;
        RECT  1.14 156.715 209.38 156.885 ;
        RECT  1.14 153.915 209.38 154.085 ;
        RECT  1.14 151.115 209.38 151.285 ;
        RECT  1.14 148.315 209.38 148.485 ;
        RECT  1.14 145.515 209.38 145.685 ;
        RECT  1.14 142.715 209.38 142.885 ;
        RECT  1.14 139.915 209.38 140.085 ;
        RECT  1.14 137.115 209.38 137.285 ;
        RECT  1.14 134.315 209.38 134.485 ;
        RECT  1.14 131.515 209.38 131.685 ;
        RECT  1.14 128.715 209.38 128.885 ;
        RECT  1.14 125.915 209.38 126.085 ;
        RECT  1.14 123.115 209.38 123.285 ;
        RECT  1.14 120.315 209.38 120.485 ;
        RECT  1.14 117.515 209.38 117.685 ;
        RECT  1.14 114.715 209.38 114.885 ;
        RECT  1.14 111.915 209.38 112.085 ;
        RECT  1.14 109.115 209.38 109.285 ;
        RECT  1.14 106.315 209.38 106.485 ;
        RECT  1.14 103.515 209.38 103.685 ;
        RECT  1.14 100.715 209.38 100.885 ;
        RECT  1.14 97.915 209.38 98.085 ;
        RECT  1.14 95.115 209.38 95.285 ;
        RECT  1.14 92.315 209.38 92.485 ;
        RECT  1.14 89.515 209.38 89.685 ;
        RECT  1.14 86.715 209.38 86.885 ;
        RECT  1.14 83.915 209.38 84.085 ;
        RECT  1.14 81.115 209.38 81.285 ;
        RECT  1.14 78.315 209.38 78.485 ;
        RECT  1.14 75.515 209.38 75.685 ;
        RECT  1.14 72.715 209.38 72.885 ;
        RECT  1.14 69.915 209.38 70.085 ;
        RECT  1.14 67.115 209.38 67.285 ;
        RECT  1.14 64.315 209.38 64.485 ;
        RECT  1.14 61.515 209.38 61.685 ;
        RECT  1.14 58.715 209.38 58.885 ;
        RECT  1.14 55.915 209.38 56.085 ;
        RECT  1.14 53.115 209.38 53.285 ;
        RECT  1.14 50.315 209.38 50.485 ;
        RECT  1.14 47.515 209.38 47.685 ;
        RECT  1.14 44.715 209.38 44.885 ;
        RECT  1.14 41.915 209.38 42.085 ;
        RECT  1.14 39.115 209.38 39.285 ;
        RECT  1.14 36.315 209.38 36.485 ;
        RECT  1.14 33.515 209.38 33.685 ;
        RECT  1.14 30.715 209.38 30.885 ;
        RECT  1.14 27.915 209.38 28.085 ;
        RECT  1.14 25.115 209.38 25.285 ;
        RECT  1.14 22.315 209.38 22.485 ;
        RECT  1.14 19.515 209.38 19.685 ;
        RECT  1.14 16.715 209.38 16.885 ;
        RECT  1.14 13.915 209.38 14.085 ;
        RECT  1.14 11.115 209.38 11.285 ;
        RECT  1.14 8.315 209.38 8.485 ;
        RECT  1.14 5.515 209.38 5.685 ;
        RECT  1.14 2.715 209.38 2.885 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 415.715 209.38 415.885 ;
        RECT  1.14 412.915 209.38 413.085 ;
        RECT  1.14 410.115 209.38 410.285 ;
        RECT  1.14 407.315 209.38 407.485 ;
        RECT  1.14 404.515 209.38 404.685 ;
        RECT  1.14 401.715 209.38 401.885 ;
        RECT  1.14 398.915 209.38 399.085 ;
        RECT  1.14 396.115 209.38 396.285 ;
        RECT  1.14 393.315 209.38 393.485 ;
        RECT  1.14 390.515 209.38 390.685 ;
        RECT  1.14 387.715 209.38 387.885 ;
        RECT  1.14 384.915 209.38 385.085 ;
        RECT  1.14 382.115 209.38 382.285 ;
        RECT  1.14 379.315 209.38 379.485 ;
        RECT  1.14 376.515 209.38 376.685 ;
        RECT  1.14 373.715 209.38 373.885 ;
        RECT  1.14 370.915 209.38 371.085 ;
        RECT  1.14 368.115 209.38 368.285 ;
        RECT  1.14 365.315 209.38 365.485 ;
        RECT  1.14 362.515 209.38 362.685 ;
        RECT  1.14 359.715 209.38 359.885 ;
        RECT  1.14 356.915 209.38 357.085 ;
        RECT  1.14 354.115 209.38 354.285 ;
        RECT  1.14 351.315 209.38 351.485 ;
        RECT  1.14 348.515 209.38 348.685 ;
        RECT  1.14 345.715 209.38 345.885 ;
        RECT  1.14 342.915 209.38 343.085 ;
        RECT  1.14 340.115 209.38 340.285 ;
        RECT  1.14 337.315 209.38 337.485 ;
        RECT  1.14 334.515 209.38 334.685 ;
        RECT  1.14 331.715 209.38 331.885 ;
        RECT  1.14 328.915 209.38 329.085 ;
        RECT  1.14 326.115 209.38 326.285 ;
        RECT  1.14 323.315 209.38 323.485 ;
        RECT  1.14 320.515 209.38 320.685 ;
        RECT  1.14 317.715 209.38 317.885 ;
        RECT  1.14 314.915 209.38 315.085 ;
        RECT  1.14 312.115 209.38 312.285 ;
        RECT  1.14 309.315 209.38 309.485 ;
        RECT  1.14 306.515 209.38 306.685 ;
        RECT  1.14 303.715 209.38 303.885 ;
        RECT  1.14 300.915 209.38 301.085 ;
        RECT  1.14 298.115 209.38 298.285 ;
        RECT  1.14 295.315 209.38 295.485 ;
        RECT  1.14 292.515 209.38 292.685 ;
        RECT  1.14 289.715 209.38 289.885 ;
        RECT  1.14 286.915 209.38 287.085 ;
        RECT  1.14 284.115 209.38 284.285 ;
        RECT  1.14 281.315 209.38 281.485 ;
        RECT  1.14 278.515 209.38 278.685 ;
        RECT  1.14 275.715 209.38 275.885 ;
        RECT  1.14 272.915 209.38 273.085 ;
        RECT  1.14 270.115 209.38 270.285 ;
        RECT  1.14 267.315 209.38 267.485 ;
        RECT  1.14 264.515 209.38 264.685 ;
        RECT  1.14 261.715 209.38 261.885 ;
        RECT  1.14 258.915 209.38 259.085 ;
        RECT  1.14 256.115 209.38 256.285 ;
        RECT  1.14 253.315 209.38 253.485 ;
        RECT  1.14 250.515 209.38 250.685 ;
        RECT  1.14 247.715 209.38 247.885 ;
        RECT  1.14 244.915 209.38 245.085 ;
        RECT  1.14 242.115 209.38 242.285 ;
        RECT  1.14 239.315 209.38 239.485 ;
        RECT  1.14 236.515 209.38 236.685 ;
        RECT  1.14 233.715 209.38 233.885 ;
        RECT  1.14 230.915 209.38 231.085 ;
        RECT  1.14 228.115 209.38 228.285 ;
        RECT  1.14 225.315 209.38 225.485 ;
        RECT  1.14 222.515 209.38 222.685 ;
        RECT  1.14 219.715 209.38 219.885 ;
        RECT  1.14 216.915 209.38 217.085 ;
        RECT  1.14 214.115 209.38 214.285 ;
        RECT  1.14 211.315 209.38 211.485 ;
        RECT  1.14 208.515 209.38 208.685 ;
        RECT  1.14 205.715 209.38 205.885 ;
        RECT  1.14 202.915 209.38 203.085 ;
        RECT  1.14 200.115 209.38 200.285 ;
        RECT  1.14 197.315 209.38 197.485 ;
        RECT  1.14 194.515 209.38 194.685 ;
        RECT  1.14 191.715 209.38 191.885 ;
        RECT  1.14 188.915 209.38 189.085 ;
        RECT  1.14 186.115 209.38 186.285 ;
        RECT  1.14 183.315 209.38 183.485 ;
        RECT  1.14 180.515 209.38 180.685 ;
        RECT  1.14 177.715 209.38 177.885 ;
        RECT  1.14 174.915 209.38 175.085 ;
        RECT  1.14 172.115 209.38 172.285 ;
        RECT  1.14 169.315 209.38 169.485 ;
        RECT  1.14 166.515 209.38 166.685 ;
        RECT  1.14 163.715 209.38 163.885 ;
        RECT  1.14 160.915 209.38 161.085 ;
        RECT  1.14 158.115 209.38 158.285 ;
        RECT  1.14 155.315 209.38 155.485 ;
        RECT  1.14 152.515 209.38 152.685 ;
        RECT  1.14 149.715 209.38 149.885 ;
        RECT  1.14 146.915 209.38 147.085 ;
        RECT  1.14 144.115 209.38 144.285 ;
        RECT  1.14 141.315 209.38 141.485 ;
        RECT  1.14 138.515 209.38 138.685 ;
        RECT  1.14 135.715 209.38 135.885 ;
        RECT  1.14 132.915 209.38 133.085 ;
        RECT  1.14 130.115 209.38 130.285 ;
        RECT  1.14 127.315 209.38 127.485 ;
        RECT  1.14 124.515 209.38 124.685 ;
        RECT  1.14 121.715 209.38 121.885 ;
        RECT  1.14 118.915 209.38 119.085 ;
        RECT  1.14 116.115 209.38 116.285 ;
        RECT  1.14 113.315 209.38 113.485 ;
        RECT  1.14 110.515 209.38 110.685 ;
        RECT  1.14 107.715 209.38 107.885 ;
        RECT  1.14 104.915 209.38 105.085 ;
        RECT  1.14 102.115 209.38 102.285 ;
        RECT  1.14 99.315 209.38 99.485 ;
        RECT  1.14 96.515 209.38 96.685 ;
        RECT  1.14 93.715 209.38 93.885 ;
        RECT  1.14 90.915 209.38 91.085 ;
        RECT  1.14 88.115 209.38 88.285 ;
        RECT  1.14 85.315 209.38 85.485 ;
        RECT  1.14 82.515 209.38 82.685 ;
        RECT  1.14 79.715 209.38 79.885 ;
        RECT  1.14 76.915 209.38 77.085 ;
        RECT  1.14 74.115 209.38 74.285 ;
        RECT  1.14 71.315 209.38 71.485 ;
        RECT  1.14 68.515 209.38 68.685 ;
        RECT  1.14 65.715 209.38 65.885 ;
        RECT  1.14 62.915 209.38 63.085 ;
        RECT  1.14 60.115 209.38 60.285 ;
        RECT  1.14 57.315 209.38 57.485 ;
        RECT  1.14 54.515 209.38 54.685 ;
        RECT  1.14 51.715 209.38 51.885 ;
        RECT  1.14 48.915 209.38 49.085 ;
        RECT  1.14 46.115 209.38 46.285 ;
        RECT  1.14 43.315 209.38 43.485 ;
        RECT  1.14 40.515 209.38 40.685 ;
        RECT  1.14 37.715 209.38 37.885 ;
        RECT  1.14 34.915 209.38 35.085 ;
        RECT  1.14 32.115 209.38 32.285 ;
        RECT  1.14 29.315 209.38 29.485 ;
        RECT  1.14 26.515 209.38 26.685 ;
        RECT  1.14 23.715 209.38 23.885 ;
        RECT  1.14 20.915 209.38 21.085 ;
        RECT  1.14 18.115 209.38 18.285 ;
        RECT  1.14 15.315 209.38 15.485 ;
        RECT  1.14 12.515 209.38 12.685 ;
        RECT  1.14 9.715 209.38 9.885 ;
        RECT  1.14 6.915 209.38 7.085 ;
        RECT  1.14 4.115 209.38 4.285 ;
        RECT  1.14 1.315 209.38 1.485 ;
    END
  END VSS
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 135.835 210.39 135.905 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 206.395 210.39 206.465 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 319.235 210.39 319.305 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 183.995 0.07 184.065 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 99.435 0.07 99.505 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  141.145 0 141.285 0.14 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  68.905 418.64 69.045 418.78 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  209.465 418.64 209.605 418.78 ;
    END
  END addr[7]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 155.995 0.07 156.065 ;
    END
  END clk
  PIN rd_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 107.555 210.39 107.625 ;
    END
  END rd_data[0]
  PIN rd_data[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 192.115 210.39 192.185 ;
    END
  END rd_data[10]
  PIN rd_data[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 234.675 210.39 234.745 ;
    END
  END rd_data[11]
  PIN rd_data[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 347.515 210.39 347.585 ;
    END
  END rd_data[12]
  PIN rd_data[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 361.515 210.39 361.585 ;
    END
  END rd_data[13]
  PIN rd_data[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 353.395 0.07 353.465 ;
    END
  END rd_data[14]
  PIN rd_data[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 212.275 0.07 212.345 ;
    END
  END rd_data[15]
  PIN rd_data[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  197.705 0 197.845 0.14 ;
    END
  END rd_data[16]
  PIN rd_data[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 28.875 0.07 28.945 ;
    END
  END rd_data[17]
  PIN rd_data[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 220.395 210.39 220.465 ;
    END
  END rd_data[18]
  PIN rd_data[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 14.875 0.07 14.945 ;
    END
  END rd_data[19]
  PIN rd_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 304.955 210.39 305.025 ;
    END
  END rd_data[1]
  PIN rd_data[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 333.235 210.39 333.305 ;
    END
  END rd_data[20]
  PIN rd_data[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 93.555 210.39 93.625 ;
    END
  END rd_data[21]
  PIN rd_data[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 240.555 0.07 240.625 ;
    END
  END rd_data[22]
  PIN rd_data[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 311.115 0.07 311.185 ;
    END
  END rd_data[23]
  PIN rd_data[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 51.275 210.39 51.345 ;
    END
  END rd_data[24]
  PIN rd_data[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 169.995 0.07 170.065 ;
    END
  END rd_data[25]
  PIN rd_data[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 282.835 0.07 282.905 ;
    END
  END rd_data[26]
  PIN rd_data[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 198.275 0.07 198.345 ;
    END
  END rd_data[27]
  PIN rd_data[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  40.345 418.64 40.485 418.78 ;
    END
  END rd_data[28]
  PIN rd_data[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 43.155 0.07 43.225 ;
    END
  END rd_data[29]
  PIN rd_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  113.145 0 113.285 0.14 ;
    END
  END rd_data[2]
  PIN rd_data[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 57.155 0.07 57.225 ;
    END
  END rd_data[30]
  PIN rd_data[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 268.835 0.07 268.905 ;
    END
  END rd_data[31]
  PIN rd_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 149.835 210.39 149.905 ;
    END
  END rd_data[3]
  PIN rd_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 381.675 0.07 381.745 ;
    END
  END rd_data[4]
  PIN rd_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  181.465 418.64 181.605 418.78 ;
    END
  END rd_data[5]
  PIN rd_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 121.835 210.39 121.905 ;
    END
  END rd_data[6]
  PIN rd_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 395.675 0.07 395.745 ;
    END
  END rd_data[7]
  PIN rd_data[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 178.115 210.39 178.185 ;
    END
  END rd_data[8]
  PIN rd_data[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 248.675 210.39 248.745 ;
    END
  END rd_data[9]
  PIN wr_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 65.275 210.39 65.345 ;
    END
  END wr_data[0]
  PIN wr_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 262.675 210.39 262.745 ;
    END
  END wr_data[10]
  PIN wr_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 367.395 0.07 367.465 ;
    END
  END wr_data[11]
  PIN wr_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.345 418.64 12.485 418.78 ;
    END
  END wr_data[12]
  PIN wr_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 254.555 0.07 254.625 ;
    END
  END wr_data[13]
  PIN wr_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END wr_data[14]
  PIN wr_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 127.715 0.07 127.785 ;
    END
  END wr_data[15]
  PIN wr_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 409.675 0.07 409.745 ;
    END
  END wr_data[16]
  PIN wr_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  96.905 418.64 97.045 418.78 ;
    END
  END wr_data[17]
  PIN wr_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 403.795 210.39 403.865 ;
    END
  END wr_data[18]
  PIN wr_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 339.395 0.07 339.465 ;
    END
  END wr_data[19]
  PIN wr_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  56.585 0 56.725 0.14 ;
    END
  END wr_data[1]
  PIN wr_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  28.585 0 28.725 0.14 ;
    END
  END wr_data[20]
  PIN wr_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 389.795 210.39 389.865 ;
    END
  END wr_data[21]
  PIN wr_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 113.715 0.07 113.785 ;
    END
  END wr_data[22]
  PIN wr_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 8.995 210.39 9.065 ;
    END
  END wr_data[23]
  PIN wr_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 375.515 210.39 375.585 ;
    END
  END wr_data[24]
  PIN wr_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 164.115 210.39 164.185 ;
    END
  END wr_data[25]
  PIN wr_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 71.155 0.07 71.225 ;
    END
  END wr_data[26]
  PIN wr_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 141.715 0.07 141.785 ;
    END
  END wr_data[27]
  PIN wr_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  85.145 0 85.285 0.14 ;
    END
  END wr_data[28]
  PIN wr_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  169.705 0 169.845 0.14 ;
    END
  END wr_data[29]
  PIN wr_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 22.995 210.39 23.065 ;
    END
  END wr_data[2]
  PIN wr_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 290.955 210.39 291.025 ;
    END
  END wr_data[30]
  PIN wr_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 36.995 210.39 37.065 ;
    END
  END wr_data[31]
  PIN wr_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  153.465 418.64 153.605 418.78 ;
    END
  END wr_data[3]
  PIN wr_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  124.905 418.64 125.045 418.78 ;
    END
  END wr_data[4]
  PIN wr_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 296.835 0.07 296.905 ;
    END
  END wr_data[5]
  PIN wr_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 325.115 0.07 325.185 ;
    END
  END wr_data[6]
  PIN wr_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 79.275 210.39 79.345 ;
    END
  END wr_data[7]
  PIN wr_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 85.435 0.07 85.505 ;
    END
  END wr_data[8]
  PIN wr_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 226.555 0.07 226.625 ;
    END
  END wr_data[9]
  PIN wr_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  210.32 276.955 210.39 277.025 ;
    END
  END wr_en
  OBS
    LAYER metal1 ;
     RECT  0 -0.085 4.75 418.78 ;
     RECT  4.75 0 210.39 418.78 ;
    LAYER metal2 ;
     RECT  0 0 210.39 418.78 ;
    LAYER metal3 ;
     RECT  0 0 210.39 418.78 ;
    LAYER metal4 ;
     RECT  0 0 210.39 418.78 ;
  END
END small_mem_block
END LIBRARY
