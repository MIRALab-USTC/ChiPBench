// Name: Black Parrot
//
// Description: 64-bit RISC-V Core with Cache Coherence Directory.
//
// Top Module: bp_multi_top
//
// GitHub: https://github.com/black-parrot/pre-alpha-release
//    commit: dbe4def684cbaf836b675ec480119d198f168c4e
//

module instr_scan_eaddr_width_p64_instr_width_p32
(
  instr_i,
  scan_o
);

  input [31:0] instr_i;
  output [68:0] scan_o;
  wire [68:0] scan_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,
  N23,N24,N25,N26,N27,N28,N29,N30;
  assign scan_o[66] = 1'b0;
  assign scan_o[67] = 1'b0;
  assign N7 = instr_i[0] & instr_i[1];
  assign scan_o[68] = ~N7;
  assign N9 = ~instr_i[6];
  assign N10 = ~instr_i[5];
  assign N11 = ~instr_i[3];
  assign N12 = ~instr_i[2];
  assign N13 = ~instr_i[1];
  assign N14 = ~instr_i[0];
  assign N15 = N10 | N9;
  assign N16 = instr_i[4] | N15;
  assign N17 = N11 | N16;
  assign N18 = N12 | N17;
  assign N19 = N13 | N18;
  assign N20 = N14 | N19;
  assign N21 = ~N20;
  assign N22 = instr_i[3] | N16;
  assign N23 = N12 | N22;
  assign N24 = N13 | N23;
  assign N25 = N14 | N24;
  assign N26 = ~N25;
  assign N27 = instr_i[2] | N22;
  assign N28 = N13 | N27;
  assign N29 = N14 | N28;
  assign N30 = ~N29;
  assign scan_o[65:64] = (N0)? { 1'b0, 1'b0 } :
                         (N1)? { 1'b0, 1'b1 } :
                         (N4)? { 1'b1, N20 } : 1'b0;
  assign N0 = N30;
  assign N1 = N26;
  assign scan_o[63:0] = (N0)? { instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[7:7], instr_i[30:25], instr_i[11:8], 1'b0 } :
                        (N1)? { instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:20] } :
                        (N2)? { instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[31:31], instr_i[19:12], instr_i[20:20], instr_i[30:21], 1'b0 } :
                        (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2 = N21;
  assign N3 = N26 | N30;
  assign N4 = ~N3;
  assign N5 = N21 | N3;
  assign N6 = ~N5;

endmodule



module bp_fe_bht_bht_indx_width_p5
(
  clk_i,
  en_i,
  reset_i,
  idx_r_i,
  idx_w_i,
  r_v_i,
  w_v_i,
  correct_i,
  predict_o
);

  input [4:0] idx_r_i;
  input [4:0] idx_w_i;
  input clk_i;
  input en_i;
  input reset_i;
  input r_v_i;
  input w_v_i;
  input correct_i;
  output predict_o;
  wire predict_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,
  N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,
  N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,
  N404,N405,N406,N407,N408,N409,N410,N411,N412,N413;
  reg [63:0] mem;
  assign predict_o = (N52)? mem[1] :
                     (N54)? mem[3] :
                     (N56)? mem[5] :
                     (N58)? mem[7] :
                     (N60)? mem[9] :
                     (N62)? mem[11] :
                     (N64)? mem[13] :
                     (N66)? mem[15] :
                     (N68)? mem[17] :
                     (N70)? mem[19] :
                     (N72)? mem[21] :
                     (N74)? mem[23] :
                     (N76)? mem[25] :
                     (N78)? mem[27] :
                     (N80)? mem[29] :
                     (N82)? mem[31] :
                     (N53)? mem[33] :
                     (N55)? mem[35] :
                     (N57)? mem[37] :
                     (N59)? mem[39] :
                     (N61)? mem[41] :
                     (N63)? mem[43] :
                     (N65)? mem[45] :
                     (N67)? mem[47] :
                     (N69)? mem[49] :
                     (N71)? mem[51] :
                     (N73)? mem[53] :
                     (N75)? mem[55] :
                     (N77)? mem[57] :
                     (N79)? mem[59] :
                     (N81)? mem[61] :
                     (N83)? mem[63] : 1'b0;
  assign N87 = (N147)? mem[1] :
               (N148)? mem[3] :
               (N149)? mem[5] :
               (N150)? mem[7] :
               (N151)? mem[9] :
               (N152)? mem[11] :
               (N153)? mem[13] :
               (N154)? mem[15] :
               (N155)? mem[17] :
               (N156)? mem[19] :
               (N157)? mem[21] :
               (N158)? mem[23] :
               (N159)? mem[25] :
               (N160)? mem[27] :
               (N161)? mem[29] :
               (N162)? mem[31] :
               (N123)? mem[33] :
               (N125)? mem[35] :
               (N127)? mem[37] :
               (N129)? mem[39] :
               (N131)? mem[41] :
               (N133)? mem[43] :
               (N135)? mem[45] :
               (N137)? mem[47] :
               (N272)? mem[49] :
               (N274)? mem[51] :
               (N276)? mem[53] :
               (N278)? mem[55] :
               (N280)? mem[57] :
               (N282)? mem[59] :
               (N284)? mem[61] :
               (N286)? mem[63] : 1'b0;
  assign N88 = (N147)? mem[0] :
               (N148)? mem[2] :
               (N149)? mem[4] :
               (N150)? mem[6] :
               (N151)? mem[8] :
               (N152)? mem[10] :
               (N153)? mem[12] :
               (N154)? mem[14] :
               (N155)? mem[16] :
               (N156)? mem[18] :
               (N157)? mem[20] :
               (N158)? mem[22] :
               (N159)? mem[24] :
               (N160)? mem[26] :
               (N161)? mem[28] :
               (N162)? mem[30] :
               (N123)? mem[32] :
               (N125)? mem[34] :
               (N127)? mem[36] :
               (N129)? mem[38] :
               (N131)? mem[40] :
               (N133)? mem[42] :
               (N135)? mem[44] :
               (N137)? mem[46] :
               (N272)? mem[48] :
               (N274)? mem[50] :
               (N276)? mem[52] :
               (N278)? mem[54] :
               (N280)? mem[56] :
               (N282)? mem[58] :
               (N284)? mem[60] :
               (N286)? mem[62] : 1'b0;
  assign N92 = N89 & N90;
  assign N93 = N92 & N91;
  assign N94 = correct_i | N87;
  assign N95 = N94 | N91;
  assign N97 = correct_i | N90;
  assign N98 = N97 | N88;
  assign N100 = N97 | N91;
  assign N102 = N89 | N87;
  assign N103 = N102 | N88;
  assign N105 = N102 | N91;
  assign N107 = N89 | N90;
  assign N108 = N107 | N88;
  assign N110 = correct_i & N87;
  assign N111 = N110 & N88;
  assign N146 = (N122)? mem[1] :
                (N124)? mem[3] :
                (N126)? mem[5] :
                (N128)? mem[7] :
                (N130)? mem[9] :
                (N132)? mem[11] :
                (N134)? mem[13] :
                (N136)? mem[15] :
                (N138)? mem[17] :
                (N139)? mem[19] :
                (N140)? mem[21] :
                (N141)? mem[23] :
                (N142)? mem[25] :
                (N143)? mem[27] :
                (N144)? mem[29] :
                (N145)? mem[31] :
                (N123)? mem[33] :
                (N125)? mem[35] :
                (N127)? mem[37] :
                (N129)? mem[39] :
                (N131)? mem[41] :
                (N133)? mem[43] :
                (N135)? mem[45] :
                (N137)? mem[47] :
                (N272)? mem[49] :
                (N274)? mem[51] :
                (N276)? mem[53] :
                (N278)? mem[55] :
                (N280)? mem[57] :
                (N282)? mem[59] :
                (N284)? mem[61] :
                (N286)? mem[63] : 1'b0;
  assign N163 = (N147)? mem[0] :
                (N148)? mem[2] :
                (N149)? mem[4] :
                (N150)? mem[6] :
                (N151)? mem[8] :
                (N152)? mem[10] :
                (N153)? mem[12] :
                (N154)? mem[14] :
                (N155)? mem[16] :
                (N156)? mem[18] :
                (N157)? mem[20] :
                (N158)? mem[22] :
                (N159)? mem[24] :
                (N160)? mem[26] :
                (N161)? mem[28] :
                (N162)? mem[30] :
                (N123)? mem[32] :
                (N125)? mem[34] :
                (N127)? mem[36] :
                (N129)? mem[38] :
                (N131)? mem[40] :
                (N133)? mem[42] :
                (N135)? mem[44] :
                (N137)? mem[46] :
                (N272)? mem[48] :
                (N274)? mem[50] :
                (N276)? mem[52] :
                (N278)? mem[54] :
                (N280)? mem[56] :
                (N282)? mem[58] :
                (N284)? mem[60] :
                (N286)? mem[62] : 1'b0;
  assign N205 = (N197)? mem[1] :
                (N198)? mem[3] :
                (N199)? mem[5] :
                (N200)? mem[7] :
                (N201)? mem[9] :
                (N202)? mem[11] :
                (N203)? mem[13] :
                (N204)? mem[15] :
                (N155)? mem[17] :
                (N156)? mem[19] :
                (N157)? mem[21] :
                (N158)? mem[23] :
                (N159)? mem[25] :
                (N160)? mem[27] :
                (N161)? mem[29] :
                (N162)? mem[31] :
                (N256)? mem[33] :
                (N258)? mem[35] :
                (N260)? mem[37] :
                (N262)? mem[39] :
                (N264)? mem[41] :
                (N266)? mem[43] :
                (N268)? mem[45] :
                (N270)? mem[47] :
                (N272)? mem[49] :
                (N274)? mem[51] :
                (N276)? mem[53] :
                (N278)? mem[55] :
                (N280)? mem[57] :
                (N282)? mem[59] :
                (N284)? mem[61] :
                (N286)? mem[63] : 1'b0;
  assign N214 = (N206)? mem[0] :
                (N207)? mem[2] :
                (N208)? mem[4] :
                (N209)? mem[6] :
                (N210)? mem[8] :
                (N211)? mem[10] :
                (N212)? mem[12] :
                (N213)? mem[14] :
                (N138)? mem[16] :
                (N139)? mem[18] :
                (N140)? mem[20] :
                (N141)? mem[22] :
                (N142)? mem[24] :
                (N143)? mem[26] :
                (N144)? mem[28] :
                (N145)? mem[30] :
                (N256)? mem[32] :
                (N258)? mem[34] :
                (N260)? mem[36] :
                (N262)? mem[38] :
                (N264)? mem[40] :
                (N266)? mem[42] :
                (N268)? mem[44] :
                (N270)? mem[46] :
                (N272)? mem[48] :
                (N274)? mem[50] :
                (N276)? mem[52] :
                (N278)? mem[54] :
                (N280)? mem[56] :
                (N282)? mem[58] :
                (N284)? mem[60] :
                (N286)? mem[62] : 1'b0;
  assign N216 = (N206)? mem[1] :
                (N207)? mem[3] :
                (N208)? mem[5] :
                (N209)? mem[7] :
                (N210)? mem[9] :
                (N211)? mem[11] :
                (N212)? mem[13] :
                (N213)? mem[15] :
                (N138)? mem[17] :
                (N139)? mem[19] :
                (N140)? mem[21] :
                (N141)? mem[23] :
                (N142)? mem[25] :
                (N143)? mem[27] :
                (N144)? mem[29] :
                (N145)? mem[31] :
                (N256)? mem[33] :
                (N258)? mem[35] :
                (N260)? mem[37] :
                (N262)? mem[39] :
                (N264)? mem[41] :
                (N266)? mem[43] :
                (N268)? mem[45] :
                (N270)? mem[47] :
                (N272)? mem[49] :
                (N274)? mem[51] :
                (N276)? mem[53] :
                (N278)? mem[55] :
                (N280)? mem[57] :
                (N282)? mem[59] :
                (N284)? mem[61] :
                (N286)? mem[63] : 1'b0;
  assign N217 = (N206)? mem[0] :
                (N207)? mem[2] :
                (N208)? mem[4] :
                (N209)? mem[6] :
                (N210)? mem[8] :
                (N211)? mem[10] :
                (N212)? mem[12] :
                (N213)? mem[14] :
                (N138)? mem[16] :
                (N139)? mem[18] :
                (N140)? mem[20] :
                (N141)? mem[22] :
                (N142)? mem[24] :
                (N143)? mem[26] :
                (N144)? mem[28] :
                (N145)? mem[30] :
                (N256)? mem[32] :
                (N258)? mem[34] :
                (N260)? mem[36] :
                (N262)? mem[38] :
                (N264)? mem[40] :
                (N266)? mem[42] :
                (N268)? mem[44] :
                (N270)? mem[46] :
                (N272)? mem[48] :
                (N274)? mem[50] :
                (N276)? mem[52] :
                (N278)? mem[54] :
                (N280)? mem[56] :
                (N282)? mem[58] :
                (N284)? mem[60] :
                (N286)? mem[62] : 1'b0;
  assign N219 = (N206)? mem[1] :
                (N207)? mem[3] :
                (N208)? mem[5] :
                (N209)? mem[7] :
                (N210)? mem[9] :
                (N211)? mem[11] :
                (N212)? mem[13] :
                (N213)? mem[15] :
                (N138)? mem[17] :
                (N139)? mem[19] :
                (N140)? mem[21] :
                (N141)? mem[23] :
                (N142)? mem[25] :
                (N143)? mem[27] :
                (N144)? mem[29] :
                (N145)? mem[31] :
                (N256)? mem[33] :
                (N258)? mem[35] :
                (N260)? mem[37] :
                (N262)? mem[39] :
                (N264)? mem[41] :
                (N266)? mem[43] :
                (N268)? mem[45] :
                (N270)? mem[47] :
                (N272)? mem[49] :
                (N274)? mem[51] :
                (N276)? mem[53] :
                (N278)? mem[55] :
                (N280)? mem[57] :
                (N282)? mem[59] :
                (N284)? mem[61] :
                (N286)? mem[63] : 1'b0;
  assign N220 = (N206)? mem[0] :
                (N207)? mem[2] :
                (N208)? mem[4] :
                (N209)? mem[6] :
                (N210)? mem[8] :
                (N211)? mem[10] :
                (N212)? mem[12] :
                (N213)? mem[14] :
                (N138)? mem[16] :
                (N139)? mem[18] :
                (N140)? mem[20] :
                (N141)? mem[22] :
                (N142)? mem[24] :
                (N143)? mem[26] :
                (N144)? mem[28] :
                (N145)? mem[30] :
                (N256)? mem[32] :
                (N258)? mem[34] :
                (N260)? mem[36] :
                (N262)? mem[38] :
                (N264)? mem[40] :
                (N266)? mem[42] :
                (N268)? mem[44] :
                (N270)? mem[46] :
                (N272)? mem[48] :
                (N274)? mem[50] :
                (N276)? mem[52] :
                (N278)? mem[54] :
                (N280)? mem[56] :
                (N282)? mem[58] :
                (N284)? mem[60] :
                (N286)? mem[62] : 1'b0;
  assign N222 = (N255)? mem[1] :
                (N257)? mem[3] :
                (N259)? mem[5] :
                (N261)? mem[7] :
                (N263)? mem[9] :
                (N265)? mem[11] :
                (N267)? mem[13] :
                (N269)? mem[15] :
                (N271)? mem[17] :
                (N273)? mem[19] :
                (N275)? mem[21] :
                (N277)? mem[23] :
                (N279)? mem[25] :
                (N281)? mem[27] :
                (N283)? mem[29] :
                (N285)? mem[31] :
                (N256)? mem[33] :
                (N258)? mem[35] :
                (N260)? mem[37] :
                (N262)? mem[39] :
                (N264)? mem[41] :
                (N266)? mem[43] :
                (N268)? mem[45] :
                (N270)? mem[47] :
                (N272)? mem[49] :
                (N274)? mem[51] :
                (N276)? mem[53] :
                (N278)? mem[55] :
                (N280)? mem[57] :
                (N282)? mem[59] :
                (N284)? mem[61] :
                (N286)? mem[63] : 1'b0;
  assign N223 = (N255)? mem[0] :
                (N257)? mem[2] :
                (N259)? mem[4] :
                (N261)? mem[6] :
                (N263)? mem[8] :
                (N265)? mem[10] :
                (N267)? mem[12] :
                (N269)? mem[14] :
                (N271)? mem[16] :
                (N273)? mem[18] :
                (N275)? mem[20] :
                (N277)? mem[22] :
                (N279)? mem[24] :
                (N281)? mem[26] :
                (N283)? mem[28] :
                (N285)? mem[30] :
                (N256)? mem[32] :
                (N258)? mem[34] :
                (N260)? mem[36] :
                (N262)? mem[38] :
                (N264)? mem[40] :
                (N266)? mem[42] :
                (N268)? mem[44] :
                (N270)? mem[46] :
                (N272)? mem[48] :
                (N274)? mem[50] :
                (N276)? mem[52] :
                (N278)? mem[54] :
                (N280)? mem[56] :
                (N282)? mem[58] :
                (N284)? mem[60] :
                (N286)? mem[62] : 1'b0;
  assign N287 = (N255)? mem[1] :
                (N257)? mem[3] :
                (N259)? mem[5] :
                (N261)? mem[7] :
                (N263)? mem[9] :
                (N265)? mem[11] :
                (N267)? mem[13] :
                (N269)? mem[15] :
                (N271)? mem[17] :
                (N273)? mem[19] :
                (N275)? mem[21] :
                (N277)? mem[23] :
                (N279)? mem[25] :
                (N281)? mem[27] :
                (N283)? mem[29] :
                (N285)? mem[31] :
                (N256)? mem[33] :
                (N258)? mem[35] :
                (N260)? mem[37] :
                (N262)? mem[39] :
                (N264)? mem[41] :
                (N266)? mem[43] :
                (N268)? mem[45] :
                (N270)? mem[47] :
                (N272)? mem[49] :
                (N274)? mem[51] :
                (N276)? mem[53] :
                (N278)? mem[55] :
                (N280)? mem[57] :
                (N282)? mem[59] :
                (N284)? mem[61] :
                (N286)? mem[63] : 1'b0;
  assign N288 = (N255)? mem[0] :
                (N257)? mem[2] :
                (N259)? mem[4] :
                (N261)? mem[6] :
                (N263)? mem[8] :
                (N265)? mem[10] :
                (N267)? mem[12] :
                (N269)? mem[14] :
                (N271)? mem[16] :
                (N273)? mem[18] :
                (N275)? mem[20] :
                (N277)? mem[22] :
                (N279)? mem[24] :
                (N281)? mem[26] :
                (N283)? mem[28] :
                (N285)? mem[30] :
                (N256)? mem[32] :
                (N258)? mem[34] :
                (N260)? mem[36] :
                (N262)? mem[38] :
                (N264)? mem[40] :
                (N266)? mem[42] :
                (N268)? mem[44] :
                (N270)? mem[46] :
                (N272)? mem[48] :
                (N274)? mem[50] :
                (N276)? mem[52] :
                (N278)? mem[54] :
                (N280)? mem[56] :
                (N282)? mem[58] :
                (N284)? mem[60] :
                (N286)? mem[62] : 1'b0;
  assign N290 = (N255)? mem[1] :
                (N257)? mem[3] :
                (N259)? mem[5] :
                (N261)? mem[7] :
                (N263)? mem[9] :
                (N265)? mem[11] :
                (N267)? mem[13] :
                (N269)? mem[15] :
                (N271)? mem[17] :
                (N273)? mem[19] :
                (N275)? mem[21] :
                (N277)? mem[23] :
                (N279)? mem[25] :
                (N281)? mem[27] :
                (N283)? mem[29] :
                (N285)? mem[31] :
                (N256)? mem[33] :
                (N258)? mem[35] :
                (N260)? mem[37] :
                (N262)? mem[39] :
                (N264)? mem[41] :
                (N266)? mem[43] :
                (N268)? mem[45] :
                (N270)? mem[47] :
                (N272)? mem[49] :
                (N274)? mem[51] :
                (N276)? mem[53] :
                (N278)? mem[55] :
                (N280)? mem[57] :
                (N282)? mem[59] :
                (N284)? mem[61] :
                (N286)? mem[63] : 1'b0;
  assign N291 = (N255)? mem[0] :
                (N257)? mem[2] :
                (N259)? mem[4] :
                (N261)? mem[6] :
                (N263)? mem[8] :
                (N265)? mem[10] :
                (N267)? mem[12] :
                (N269)? mem[14] :
                (N271)? mem[16] :
                (N273)? mem[18] :
                (N275)? mem[20] :
                (N277)? mem[22] :
                (N279)? mem[24] :
                (N281)? mem[26] :
                (N283)? mem[28] :
                (N285)? mem[30] :
                (N256)? mem[32] :
                (N258)? mem[34] :
                (N260)? mem[36] :
                (N262)? mem[38] :
                (N264)? mem[40] :
                (N266)? mem[42] :
                (N268)? mem[44] :
                (N270)? mem[46] :
                (N272)? mem[48] :
                (N274)? mem[50] :
                (N276)? mem[52] :
                (N278)? mem[54] :
                (N280)? mem[56] :
                (N282)? mem[58] :
                (N284)? mem[60] :
                (N286)? mem[62] : 1'b0;
  assign N292 = (N255)? mem[1] :
                (N257)? mem[3] :
                (N259)? mem[5] :
                (N261)? mem[7] :
                (N263)? mem[9] :
                (N265)? mem[11] :
                (N267)? mem[13] :
                (N269)? mem[15] :
                (N271)? mem[17] :
                (N273)? mem[19] :
                (N275)? mem[21] :
                (N277)? mem[23] :
                (N279)? mem[25] :
                (N281)? mem[27] :
                (N283)? mem[29] :
                (N285)? mem[31] :
                (N256)? mem[33] :
                (N258)? mem[35] :
                (N260)? mem[37] :
                (N262)? mem[39] :
                (N264)? mem[41] :
                (N266)? mem[43] :
                (N268)? mem[45] :
                (N270)? mem[47] :
                (N272)? mem[49] :
                (N274)? mem[51] :
                (N276)? mem[53] :
                (N278)? mem[55] :
                (N280)? mem[57] :
                (N282)? mem[59] :
                (N284)? mem[61] :
                (N286)? mem[63] : 1'b0;
  assign N293 = (N255)? mem[0] :
                (N257)? mem[2] :
                (N259)? mem[4] :
                (N261)? mem[6] :
                (N263)? mem[8] :
                (N265)? mem[10] :
                (N267)? mem[12] :
                (N269)? mem[14] :
                (N271)? mem[16] :
                (N273)? mem[18] :
                (N275)? mem[20] :
                (N277)? mem[22] :
                (N279)? mem[24] :
                (N281)? mem[26] :
                (N283)? mem[28] :
                (N285)? mem[30] :
                (N256)? mem[32] :
                (N258)? mem[34] :
                (N260)? mem[36] :
                (N262)? mem[38] :
                (N264)? mem[40] :
                (N266)? mem[42] :
                (N268)? mem[44] :
                (N270)? mem[46] :
                (N272)? mem[48] :
                (N274)? mem[50] :
                (N276)? mem[52] :
                (N278)? mem[54] :
                (N280)? mem[56] :
                (N282)? mem[58] :
                (N284)? mem[60] :
                (N286)? mem[62] : 1'b0;
  assign N397 = idx_w_i[3] & idx_w_i[4];
  assign N398 = N0 & idx_w_i[4];
  assign N0 = ~idx_w_i[3];
  assign N399 = idx_w_i[3] & N1;
  assign N1 = ~idx_w_i[4];
  assign N400 = N2 & N3;
  assign N2 = ~idx_w_i[3];
  assign N3 = ~idx_w_i[4];
  assign N401 = ~idx_w_i[2];
  assign N402 = idx_w_i[0] & idx_w_i[1];
  assign N403 = N4 & idx_w_i[1];
  assign N4 = ~idx_w_i[0];
  assign N404 = idx_w_i[0] & N5;
  assign N5 = ~idx_w_i[1];
  assign N405 = N6 & N7;
  assign N6 = ~idx_w_i[0];
  assign N7 = ~idx_w_i[1];
  assign N406 = idx_w_i[2] & N402;
  assign N407 = idx_w_i[2] & N403;
  assign N408 = idx_w_i[2] & N404;
  assign N409 = idx_w_i[2] & N405;
  assign N410 = N401 & N402;
  assign N411 = N401 & N403;
  assign N412 = N401 & N404;
  assign N413 = N401 & N405;
  assign N195 = N397 & N406;
  assign N194 = N397 & N407;
  assign N193 = N397 & N408;
  assign N192 = N397 & N409;
  assign N191 = N397 & N410;
  assign N190 = N397 & N411;
  assign N189 = N397 & N412;
  assign N188 = N397 & N413;
  assign N187 = N398 & N406;
  assign N186 = N398 & N407;
  assign N185 = N398 & N408;
  assign N184 = N398 & N409;
  assign N183 = N398 & N410;
  assign N182 = N398 & N411;
  assign N181 = N398 & N412;
  assign N180 = N398 & N413;
  assign N179 = N399 & N406;
  assign N178 = N399 & N407;
  assign N177 = N399 & N408;
  assign N176 = N399 & N409;
  assign N175 = N399 & N410;
  assign N174 = N399 & N411;
  assign N173 = N399 & N412;
  assign N172 = N399 & N413;
  assign N171 = N400 & N406;
  assign N170 = N400 & N407;
  assign N169 = N400 & N408;
  assign N168 = N400 & N409;
  assign N167 = N400 & N410;
  assign N166 = N400 & N411;
  assign N165 = N400 & N412;
  assign N164 = N400 & N413;
  assign { N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N295 } = (N8)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } :
                                                                                                                                                                                                              (N9)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } :
                                                                                                                                                                                                              (N10)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } :
                                                                                                                                                                                                              (N11)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } :
                                                                                                                                                                                                              (N12)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } :
                                                                                                                                                                                                              (N13)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } :
                                                                                                                                                                                                              (N14)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } :
                                                                                                                                                                                                              (N15)? { N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164 } : 1'b0;
  assign N8 = N93;
  assign N9 = N96;
  assign N10 = N99;
  assign N11 = N101;
  assign N12 = N104;
  assign N13 = N106;
  assign N14 = N109;
  assign N15 = N111;
  assign { N297, N296 } = (N8)? { N196, 1'b1 } :
                          (N9)? { N215, 1'b1 } :
                          (N10)? { N218, 1'b1 } :
                          (N11)? { N221, 1'b1 } :
                          (N12)? { N222, N223 } :
                          (N13)? { N287, N289 } :
                          (N14)? { N290, N291 } :
                          (N15)? { N292, N294 } : 1'b0;
  assign { N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N329 } = (N16)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } :
                                                                                                                                                                                                              (N396)? { N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N295 } :
                                                                                                                                                                                                              (N86)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = reset_i;
  assign { N331, N330 } = (N16)? { 1'b0, 1'b1 } :
                          (N396)? { N297, N296 } : 1'b0;
  assign { N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363 } = (N17)? { N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N329 } :
                                                                                                                                                                                                              (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N17 = en_i;
  assign N18 = N84;
  assign N19 = ~idx_r_i[0];
  assign N20 = ~idx_r_i[1];
  assign N21 = N19 & N20;
  assign N22 = N19 & idx_r_i[1];
  assign N23 = idx_r_i[0] & N20;
  assign N24 = idx_r_i[0] & idx_r_i[1];
  assign N25 = ~idx_r_i[2];
  assign N26 = N21 & N25;
  assign N27 = N21 & idx_r_i[2];
  assign N28 = N23 & N25;
  assign N29 = N23 & idx_r_i[2];
  assign N30 = N22 & N25;
  assign N31 = N22 & idx_r_i[2];
  assign N32 = N24 & N25;
  assign N33 = N24 & idx_r_i[2];
  assign N34 = ~idx_r_i[3];
  assign N35 = N26 & N34;
  assign N36 = N26 & idx_r_i[3];
  assign N37 = N28 & N34;
  assign N38 = N28 & idx_r_i[3];
  assign N39 = N30 & N34;
  assign N40 = N30 & idx_r_i[3];
  assign N41 = N32 & N34;
  assign N42 = N32 & idx_r_i[3];
  assign N43 = N27 & N34;
  assign N44 = N27 & idx_r_i[3];
  assign N45 = N29 & N34;
  assign N46 = N29 & idx_r_i[3];
  assign N47 = N31 & N34;
  assign N48 = N31 & idx_r_i[3];
  assign N49 = N33 & N34;
  assign N50 = N33 & idx_r_i[3];
  assign N51 = ~idx_r_i[4];
  assign N52 = N35 & N51;
  assign N53 = N35 & idx_r_i[4];
  assign N54 = N37 & N51;
  assign N55 = N37 & idx_r_i[4];
  assign N56 = N39 & N51;
  assign N57 = N39 & idx_r_i[4];
  assign N58 = N41 & N51;
  assign N59 = N41 & idx_r_i[4];
  assign N60 = N43 & N51;
  assign N61 = N43 & idx_r_i[4];
  assign N62 = N45 & N51;
  assign N63 = N45 & idx_r_i[4];
  assign N64 = N47 & N51;
  assign N65 = N47 & idx_r_i[4];
  assign N66 = N49 & N51;
  assign N67 = N49 & idx_r_i[4];
  assign N68 = N36 & N51;
  assign N69 = N36 & idx_r_i[4];
  assign N70 = N38 & N51;
  assign N71 = N38 & idx_r_i[4];
  assign N72 = N40 & N51;
  assign N73 = N40 & idx_r_i[4];
  assign N74 = N42 & N51;
  assign N75 = N42 & idx_r_i[4];
  assign N76 = N44 & N51;
  assign N77 = N44 & idx_r_i[4];
  assign N78 = N46 & N51;
  assign N79 = N46 & idx_r_i[4];
  assign N80 = N48 & N51;
  assign N81 = N48 & idx_r_i[4];
  assign N82 = N50 & N51;
  assign N83 = N50 & idx_r_i[4];
  assign N84 = ~en_i;
  assign N85 = w_v_i | reset_i;
  assign N86 = ~N85;
  assign N89 = ~correct_i;
  assign N90 = ~N87;
  assign N91 = ~N88;
  assign N96 = ~N95;
  assign N99 = ~N98;
  assign N101 = ~N100;
  assign N104 = ~N103;
  assign N106 = ~N105;
  assign N109 = ~N108;
  assign N112 = ~idx_w_i[3];
  assign N113 = N231 & N112;
  assign N114 = N233 & N112;
  assign N115 = N235 & N112;
  assign N116 = N237 & N112;
  assign N117 = N232 & N112;
  assign N118 = N234 & N112;
  assign N119 = N236 & N112;
  assign N120 = N238 & N112;
  assign N121 = ~idx_w_i[4];
  assign N122 = N113 & N121;
  assign N123 = N113 & idx_w_i[4];
  assign N124 = N114 & N121;
  assign N125 = N114 & idx_w_i[4];
  assign N126 = N115 & N121;
  assign N127 = N115 & idx_w_i[4];
  assign N128 = N116 & N121;
  assign N129 = N116 & idx_w_i[4];
  assign N130 = N117 & N121;
  assign N131 = N117 & idx_w_i[4];
  assign N132 = N118 & N121;
  assign N133 = N118 & idx_w_i[4];
  assign N134 = N119 & N121;
  assign N135 = N119 & idx_w_i[4];
  assign N136 = N120 & N121;
  assign N137 = N120 & idx_w_i[4];
  assign N138 = N240 & N121;
  assign N139 = N242 & N121;
  assign N140 = N244 & N121;
  assign N141 = N246 & N121;
  assign N142 = N248 & N121;
  assign N143 = N250 & N121;
  assign N144 = N252 & N121;
  assign N145 = N254 & N121;
  assign N147 = N113 & N121;
  assign N148 = N114 & N121;
  assign N149 = N115 & N121;
  assign N150 = N116 & N121;
  assign N151 = N117 & N121;
  assign N152 = N118 & N121;
  assign N153 = N119 & N121;
  assign N154 = N120 & N121;
  assign N155 = N240 & N121;
  assign N156 = N242 & N121;
  assign N157 = N244 & N121;
  assign N158 = N246 & N121;
  assign N159 = N248 & N121;
  assign N160 = N250 & N121;
  assign N161 = N252 & N121;
  assign N162 = N254 & N121;
  assign N196 = N146 ^ N163;
  assign N197 = N239 & N121;
  assign N198 = N241 & N121;
  assign N199 = N243 & N121;
  assign N200 = N245 & N121;
  assign N201 = N247 & N121;
  assign N202 = N249 & N121;
  assign N203 = N251 & N121;
  assign N204 = N253 & N121;
  assign N206 = N239 & N121;
  assign N207 = N241 & N121;
  assign N208 = N243 & N121;
  assign N209 = N245 & N121;
  assign N210 = N247 & N121;
  assign N211 = N249 & N121;
  assign N212 = N251 & N121;
  assign N213 = N253 & N121;
  assign N215 = N205 ^ N214;
  assign N218 = N216 ^ N217;
  assign N221 = N219 ^ N220;
  assign N224 = ~idx_w_i[0];
  assign N225 = ~idx_w_i[1];
  assign N226 = N224 & N225;
  assign N227 = N224 & idx_w_i[1];
  assign N228 = idx_w_i[0] & N225;
  assign N229 = idx_w_i[0] & idx_w_i[1];
  assign N230 = ~idx_w_i[2];
  assign N231 = N226 & N230;
  assign N232 = N226 & idx_w_i[2];
  assign N233 = N228 & N230;
  assign N234 = N228 & idx_w_i[2];
  assign N235 = N227 & N230;
  assign N236 = N227 & idx_w_i[2];
  assign N237 = N229 & N230;
  assign N238 = N229 & idx_w_i[2];
  assign N239 = N231 & N112;
  assign N240 = N231 & idx_w_i[3];
  assign N241 = N233 & N112;
  assign N242 = N233 & idx_w_i[3];
  assign N243 = N235 & N112;
  assign N244 = N235 & idx_w_i[3];
  assign N245 = N237 & N112;
  assign N246 = N237 & idx_w_i[3];
  assign N247 = N232 & N112;
  assign N248 = N232 & idx_w_i[3];
  assign N249 = N234 & N112;
  assign N250 = N234 & idx_w_i[3];
  assign N251 = N236 & N112;
  assign N252 = N236 & idx_w_i[3];
  assign N253 = N238 & N112;
  assign N254 = N238 & idx_w_i[3];
  assign N255 = N239 & N121;
  assign N256 = N239 & idx_w_i[4];
  assign N257 = N241 & N121;
  assign N258 = N241 & idx_w_i[4];
  assign N259 = N243 & N121;
  assign N260 = N243 & idx_w_i[4];
  assign N261 = N245 & N121;
  assign N262 = N245 & idx_w_i[4];
  assign N263 = N247 & N121;
  assign N264 = N247 & idx_w_i[4];
  assign N265 = N249 & N121;
  assign N266 = N249 & idx_w_i[4];
  assign N267 = N251 & N121;
  assign N268 = N251 & idx_w_i[4];
  assign N269 = N253 & N121;
  assign N270 = N253 & idx_w_i[4];
  assign N271 = N240 & N121;
  assign N272 = N240 & idx_w_i[4];
  assign N273 = N242 & N121;
  assign N274 = N242 & idx_w_i[4];
  assign N275 = N244 & N121;
  assign N276 = N244 & idx_w_i[4];
  assign N277 = N246 & N121;
  assign N278 = N246 & idx_w_i[4];
  assign N279 = N248 & N121;
  assign N280 = N248 & idx_w_i[4];
  assign N281 = N250 & N121;
  assign N282 = N250 & idx_w_i[4];
  assign N283 = N252 & N121;
  assign N284 = N252 & idx_w_i[4];
  assign N285 = N254 & N121;
  assign N286 = N254 & idx_w_i[4];
  assign N289 = ~N288;
  assign N294 = ~N293;
  assign N395 = ~reset_i;
  assign N396 = w_v_i & N395;

  always @(posedge clk_i) begin
    if(N394) begin
      { mem[63:62] } <= { N331, N330 };
    end
    if(N393) begin
      { mem[61:60] } <= { N331, N330 };
    end
    if(N392) begin
      { mem[59:58] } <= { N331, N330 };
    end
    if(N391) begin
      { mem[57:56] } <= { N331, N330 };
    end
    if(N390) begin
      { mem[55:54] } <= { N331, N330 };
    end
    if(N389) begin
      { mem[53:52] } <= { N331, N330 };
    end
    if(N388) begin
      { mem[51:50] } <= { N331, N330 };
    end
    if(N387) begin
      { mem[49:48] } <= { N331, N330 };
    end
    if(N386) begin
      { mem[47:46] } <= { N331, N330 };
    end
    if(N385) begin
      { mem[45:44] } <= { N331, N330 };
    end
    if(N384) begin
      { mem[43:42] } <= { N331, N330 };
    end
    if(N383) begin
      { mem[41:40] } <= { N331, N330 };
    end
    if(N382) begin
      { mem[39:38] } <= { N331, N330 };
    end
    if(N381) begin
      { mem[37:36] } <= { N331, N330 };
    end
    if(N380) begin
      { mem[35:34] } <= { N331, N330 };
    end
    if(N379) begin
      { mem[33:32] } <= { N331, N330 };
    end
    if(N378) begin
      { mem[31:30] } <= { N331, N330 };
    end
    if(N377) begin
      { mem[29:28] } <= { N331, N330 };
    end
    if(N376) begin
      { mem[27:26] } <= { N331, N330 };
    end
    if(N375) begin
      { mem[25:24] } <= { N331, N330 };
    end
    if(N374) begin
      { mem[23:22] } <= { N331, N330 };
    end
    if(N373) begin
      { mem[21:20] } <= { N331, N330 };
    end
    if(N372) begin
      { mem[19:18] } <= { N331, N330 };
    end
    if(N371) begin
      { mem[17:16] } <= { N331, N330 };
    end
    if(N370) begin
      { mem[15:14] } <= { N331, N330 };
    end
    if(N369) begin
      { mem[13:12] } <= { N331, N330 };
    end
    if(N368) begin
      { mem[11:10] } <= { N331, N330 };
    end
    if(N367) begin
      { mem[9:8] } <= { N331, N330 };
    end
    if(N366) begin
      { mem[7:6] } <= { N331, N330 };
    end
    if(N365) begin
      { mem[5:4] } <= { N331, N330 };
    end
    if(N364) begin
      { mem[3:2] } <= { N331, N330 };
    end
    if(N363) begin
      { mem[1:0] } <= { N331, N330 };
    end
  end


endmodule



module bsg_mem_1rw_sync_width_p64_els_p512_addr_width_lp9
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_i,
  data_o
);

  input [63:0] data_i;
  input [8:0] addr_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [63:0] data_o;

  hard_mem_1rw_d512_w64_wrapper
  macro_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bp_fe_btb_bp_fe_pc_gen_btb_idx_width_lp9_eaddr_width_p64
(
  clk_i,
  reset_i,
  idx_w_i,
  idx_r_i,
  r_v_i,
  w_v_i,
  branch_target_i,
  branch_target_o,
  read_valid_o
);

  input [8:0] idx_w_i;
  input [8:0] idx_r_i;
  input [63:0] branch_target_i;
  output [63:0] branch_target_o;
  input clk_i;
  input reset_i;
  input r_v_i;
  input w_v_i;
  output read_valid_o;
  wire [63:0] branch_target_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,
  N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,
  N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,
  N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,
  N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,
  N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,
  N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,
  N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,
  N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,
  N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,
  N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,
  N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,
  N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,
  N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,
  N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,
  N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,
  N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,
  N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,
  N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,
  N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,
  N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,
  N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,
  N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,
  N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,
  N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,
  N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,
  N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,
  N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,
  N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,
  N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,
  N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,
  N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,
  N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,
  N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,
  N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,
  N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,
  N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,
  N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,
  N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,
  N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,
  N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,
  N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,
  N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,
  N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,
  N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,
  N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,
  N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,
  N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,
  N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,
  N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,
  N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,
  N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,
  N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,
  N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,
  N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,
  N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,
  N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,
  N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,
  N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,
  N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,
  N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,
  N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,
  N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,
  N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,
  N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,
  N2078,N2079,N2080,n_0_net_,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,
  N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,
  N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,
  N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,
  N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,
  N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153;
  wire [8:0] addr;
  reg [511:0] valid;
  reg read_valid_o;
  assign N2080 = (N1568)? valid[0] :
                 (N1570)? valid[1] :
                 (N1572)? valid[2] :
                 (N1574)? valid[3] :
                 (N1576)? valid[4] :
                 (N1578)? valid[5] :
                 (N1580)? valid[6] :
                 (N1582)? valid[7] :
                 (N1584)? valid[8] :
                 (N1586)? valid[9] :
                 (N1588)? valid[10] :
                 (N1590)? valid[11] :
                 (N1592)? valid[12] :
                 (N1594)? valid[13] :
                 (N1596)? valid[14] :
                 (N1598)? valid[15] :
                 (N1600)? valid[16] :
                 (N1602)? valid[17] :
                 (N1604)? valid[18] :
                 (N1606)? valid[19] :
                 (N1608)? valid[20] :
                 (N1610)? valid[21] :
                 (N1612)? valid[22] :
                 (N1614)? valid[23] :
                 (N1616)? valid[24] :
                 (N1618)? valid[25] :
                 (N1620)? valid[26] :
                 (N1622)? valid[27] :
                 (N1624)? valid[28] :
                 (N1626)? valid[29] :
                 (N1628)? valid[30] :
                 (N1630)? valid[31] :
                 (N1632)? valid[32] :
                 (N1634)? valid[33] :
                 (N1636)? valid[34] :
                 (N1638)? valid[35] :
                 (N1640)? valid[36] :
                 (N1642)? valid[37] :
                 (N1644)? valid[38] :
                 (N1646)? valid[39] :
                 (N1648)? valid[40] :
                 (N1650)? valid[41] :
                 (N1652)? valid[42] :
                 (N1654)? valid[43] :
                 (N1656)? valid[44] :
                 (N1658)? valid[45] :
                 (N1660)? valid[46] :
                 (N1662)? valid[47] :
                 (N1664)? valid[48] :
                 (N1666)? valid[49] :
                 (N1668)? valid[50] :
                 (N1670)? valid[51] :
                 (N1672)? valid[52] :
                 (N1674)? valid[53] :
                 (N1676)? valid[54] :
                 (N1678)? valid[55] :
                 (N1680)? valid[56] :
                 (N1682)? valid[57] :
                 (N1684)? valid[58] :
                 (N1686)? valid[59] :
                 (N1688)? valid[60] :
                 (N1690)? valid[61] :
                 (N1692)? valid[62] :
                 (N1694)? valid[63] :
                 (N1696)? valid[64] :
                 (N1698)? valid[65] :
                 (N1700)? valid[66] :
                 (N1702)? valid[67] :
                 (N1704)? valid[68] :
                 (N1706)? valid[69] :
                 (N1708)? valid[70] :
                 (N1710)? valid[71] :
                 (N1712)? valid[72] :
                 (N1714)? valid[73] :
                 (N1716)? valid[74] :
                 (N1718)? valid[75] :
                 (N1720)? valid[76] :
                 (N1722)? valid[77] :
                 (N1724)? valid[78] :
                 (N1726)? valid[79] :
                 (N1728)? valid[80] :
                 (N1730)? valid[81] :
                 (N1732)? valid[82] :
                 (N1734)? valid[83] :
                 (N1736)? valid[84] :
                 (N1738)? valid[85] :
                 (N1740)? valid[86] :
                 (N1742)? valid[87] :
                 (N1744)? valid[88] :
                 (N1746)? valid[89] :
                 (N1748)? valid[90] :
                 (N1750)? valid[91] :
                 (N1752)? valid[92] :
                 (N1754)? valid[93] :
                 (N1756)? valid[94] :
                 (N1758)? valid[95] :
                 (N1760)? valid[96] :
                 (N1762)? valid[97] :
                 (N1764)? valid[98] :
                 (N1766)? valid[99] :
                 (N1768)? valid[100] :
                 (N1770)? valid[101] :
                 (N1772)? valid[102] :
                 (N1774)? valid[103] :
                 (N1776)? valid[104] :
                 (N1778)? valid[105] :
                 (N1780)? valid[106] :
                 (N1782)? valid[107] :
                 (N1784)? valid[108] :
                 (N1786)? valid[109] :
                 (N1788)? valid[110] :
                 (N1790)? valid[111] :
                 (N1792)? valid[112] :
                 (N1794)? valid[113] :
                 (N1796)? valid[114] :
                 (N1798)? valid[115] :
                 (N1800)? valid[116] :
                 (N1802)? valid[117] :
                 (N1804)? valid[118] :
                 (N1806)? valid[119] :
                 (N1808)? valid[120] :
                 (N1810)? valid[121] :
                 (N1812)? valid[122] :
                 (N1814)? valid[123] :
                 (N1816)? valid[124] :
                 (N1818)? valid[125] :
                 (N1820)? valid[126] :
                 (N1822)? valid[127] :
                 (N1824)? valid[128] :
                 (N1826)? valid[129] :
                 (N1828)? valid[130] :
                 (N1830)? valid[131] :
                 (N1832)? valid[132] :
                 (N1834)? valid[133] :
                 (N1836)? valid[134] :
                 (N1838)? valid[135] :
                 (N1840)? valid[136] :
                 (N1842)? valid[137] :
                 (N1844)? valid[138] :
                 (N1846)? valid[139] :
                 (N1848)? valid[140] :
                 (N1850)? valid[141] :
                 (N1852)? valid[142] :
                 (N1854)? valid[143] :
                 (N1856)? valid[144] :
                 (N1858)? valid[145] :
                 (N1860)? valid[146] :
                 (N1862)? valid[147] :
                 (N1864)? valid[148] :
                 (N1866)? valid[149] :
                 (N1868)? valid[150] :
                 (N1870)? valid[151] :
                 (N1872)? valid[152] :
                 (N1874)? valid[153] :
                 (N1876)? valid[154] :
                 (N1878)? valid[155] :
                 (N1880)? valid[156] :
                 (N1882)? valid[157] :
                 (N1884)? valid[158] :
                 (N1886)? valid[159] :
                 (N1888)? valid[160] :
                 (N1890)? valid[161] :
                 (N1892)? valid[162] :
                 (N1894)? valid[163] :
                 (N1896)? valid[164] :
                 (N1898)? valid[165] :
                 (N1900)? valid[166] :
                 (N1902)? valid[167] :
                 (N1904)? valid[168] :
                 (N1906)? valid[169] :
                 (N1908)? valid[170] :
                 (N1910)? valid[171] :
                 (N1912)? valid[172] :
                 (N1914)? valid[173] :
                 (N1916)? valid[174] :
                 (N1918)? valid[175] :
                 (N1920)? valid[176] :
                 (N1922)? valid[177] :
                 (N1924)? valid[178] :
                 (N1926)? valid[179] :
                 (N1928)? valid[180] :
                 (N1930)? valid[181] :
                 (N1932)? valid[182] :
                 (N1934)? valid[183] :
                 (N1936)? valid[184] :
                 (N1938)? valid[185] :
                 (N1940)? valid[186] :
                 (N1942)? valid[187] :
                 (N1944)? valid[188] :
                 (N1946)? valid[189] :
                 (N1948)? valid[190] :
                 (N1950)? valid[191] :
                 (N1952)? valid[192] :
                 (N1954)? valid[193] :
                 (N1956)? valid[194] :
                 (N1958)? valid[195] :
                 (N1960)? valid[196] :
                 (N1962)? valid[197] :
                 (N1964)? valid[198] :
                 (N1966)? valid[199] :
                 (N1968)? valid[200] :
                 (N1970)? valid[201] :
                 (N1972)? valid[202] :
                 (N1974)? valid[203] :
                 (N1976)? valid[204] :
                 (N1978)? valid[205] :
                 (N1980)? valid[206] :
                 (N1982)? valid[207] :
                 (N1984)? valid[208] :
                 (N1986)? valid[209] :
                 (N1988)? valid[210] :
                 (N1990)? valid[211] :
                 (N1992)? valid[212] :
                 (N1994)? valid[213] :
                 (N1996)? valid[214] :
                 (N1998)? valid[215] :
                 (N2000)? valid[216] :
                 (N2002)? valid[217] :
                 (N2004)? valid[218] :
                 (N2006)? valid[219] :
                 (N2008)? valid[220] :
                 (N2010)? valid[221] :
                 (N2012)? valid[222] :
                 (N2014)? valid[223] :
                 (N2016)? valid[224] :
                 (N2018)? valid[225] :
                 (N2020)? valid[226] :
                 (N2022)? valid[227] :
                 (N2024)? valid[228] :
                 (N2026)? valid[229] :
                 (N2028)? valid[230] :
                 (N2030)? valid[231] :
                 (N2032)? valid[232] :
                 (N2034)? valid[233] :
                 (N2036)? valid[234] :
                 (N2038)? valid[235] :
                 (N2040)? valid[236] :
                 (N2042)? valid[237] :
                 (N2044)? valid[238] :
                 (N2046)? valid[239] :
                 (N2048)? valid[240] :
                 (N2050)? valid[241] :
                 (N2052)? valid[242] :
                 (N2054)? valid[243] :
                 (N2056)? valid[244] :
                 (N2058)? valid[245] :
                 (N2060)? valid[246] :
                 (N2062)? valid[247] :
                 (N2064)? valid[248] :
                 (N2066)? valid[249] :
                 (N2068)? valid[250] :
                 (N2070)? valid[251] :
                 (N2072)? valid[252] :
                 (N2074)? valid[253] :
                 (N2076)? valid[254] :
                 (N2078)? valid[255] :
                 (N1569)? valid[256] :
                 (N1571)? valid[257] :
                 (N1573)? valid[258] :
                 (N1575)? valid[259] :
                 (N1577)? valid[260] :
                 (N1579)? valid[261] :
                 (N1581)? valid[262] :
                 (N1583)? valid[263] :
                 (N1585)? valid[264] :
                 (N1587)? valid[265] :
                 (N1589)? valid[266] :
                 (N1591)? valid[267] :
                 (N1593)? valid[268] :
                 (N1595)? valid[269] :
                 (N1597)? valid[270] :
                 (N1599)? valid[271] :
                 (N1601)? valid[272] :
                 (N1603)? valid[273] :
                 (N1605)? valid[274] :
                 (N1607)? valid[275] :
                 (N1609)? valid[276] :
                 (N1611)? valid[277] :
                 (N1613)? valid[278] :
                 (N1615)? valid[279] :
                 (N1617)? valid[280] :
                 (N1619)? valid[281] :
                 (N1621)? valid[282] :
                 (N1623)? valid[283] :
                 (N1625)? valid[284] :
                 (N1627)? valid[285] :
                 (N1629)? valid[286] :
                 (N1631)? valid[287] :
                 (N1633)? valid[288] :
                 (N1635)? valid[289] :
                 (N1637)? valid[290] :
                 (N1639)? valid[291] :
                 (N1641)? valid[292] :
                 (N1643)? valid[293] :
                 (N1645)? valid[294] :
                 (N1647)? valid[295] :
                 (N1649)? valid[296] :
                 (N1651)? valid[297] :
                 (N1653)? valid[298] :
                 (N1655)? valid[299] :
                 (N1657)? valid[300] :
                 (N1659)? valid[301] :
                 (N1661)? valid[302] :
                 (N1663)? valid[303] :
                 (N1665)? valid[304] :
                 (N1667)? valid[305] :
                 (N1669)? valid[306] :
                 (N1671)? valid[307] :
                 (N1673)? valid[308] :
                 (N1675)? valid[309] :
                 (N1677)? valid[310] :
                 (N1679)? valid[311] :
                 (N1681)? valid[312] :
                 (N1683)? valid[313] :
                 (N1685)? valid[314] :
                 (N1687)? valid[315] :
                 (N1689)? valid[316] :
                 (N1691)? valid[317] :
                 (N1693)? valid[318] :
                 (N1695)? valid[319] :
                 (N1697)? valid[320] :
                 (N1699)? valid[321] :
                 (N1701)? valid[322] :
                 (N1703)? valid[323] :
                 (N1705)? valid[324] :
                 (N1707)? valid[325] :
                 (N1709)? valid[326] :
                 (N1711)? valid[327] :
                 (N1713)? valid[328] :
                 (N1715)? valid[329] :
                 (N1717)? valid[330] :
                 (N1719)? valid[331] :
                 (N1721)? valid[332] :
                 (N1723)? valid[333] :
                 (N1725)? valid[334] :
                 (N1727)? valid[335] :
                 (N1729)? valid[336] :
                 (N1731)? valid[337] :
                 (N1733)? valid[338] :
                 (N1735)? valid[339] :
                 (N1737)? valid[340] :
                 (N1739)? valid[341] :
                 (N1741)? valid[342] :
                 (N1743)? valid[343] :
                 (N1745)? valid[344] :
                 (N1747)? valid[345] :
                 (N1749)? valid[346] :
                 (N1751)? valid[347] :
                 (N1753)? valid[348] :
                 (N1755)? valid[349] :
                 (N1757)? valid[350] :
                 (N1759)? valid[351] :
                 (N1761)? valid[352] :
                 (N1763)? valid[353] :
                 (N1765)? valid[354] :
                 (N1767)? valid[355] :
                 (N1769)? valid[356] :
                 (N1771)? valid[357] :
                 (N1773)? valid[358] :
                 (N1775)? valid[359] :
                 (N1777)? valid[360] :
                 (N1779)? valid[361] :
                 (N1781)? valid[362] :
                 (N1783)? valid[363] :
                 (N1785)? valid[364] :
                 (N1787)? valid[365] :
                 (N1789)? valid[366] :
                 (N1791)? valid[367] :
                 (N1793)? valid[368] :
                 (N1795)? valid[369] :
                 (N1797)? valid[370] :
                 (N1799)? valid[371] :
                 (N1801)? valid[372] :
                 (N1803)? valid[373] :
                 (N1805)? valid[374] :
                 (N1807)? valid[375] :
                 (N1809)? valid[376] :
                 (N1811)? valid[377] :
                 (N1813)? valid[378] :
                 (N1815)? valid[379] :
                 (N1817)? valid[380] :
                 (N1819)? valid[381] :
                 (N1821)? valid[382] :
                 (N1823)? valid[383] :
                 (N1825)? valid[384] :
                 (N1827)? valid[385] :
                 (N1829)? valid[386] :
                 (N1831)? valid[387] :
                 (N1833)? valid[388] :
                 (N1835)? valid[389] :
                 (N1837)? valid[390] :
                 (N1839)? valid[391] :
                 (N1841)? valid[392] :
                 (N1843)? valid[393] :
                 (N1845)? valid[394] :
                 (N1847)? valid[395] :
                 (N1849)? valid[396] :
                 (N1851)? valid[397] :
                 (N1853)? valid[398] :
                 (N1855)? valid[399] :
                 (N1857)? valid[400] :
                 (N1859)? valid[401] :
                 (N1861)? valid[402] :
                 (N1863)? valid[403] :
                 (N1865)? valid[404] :
                 (N1867)? valid[405] :
                 (N1869)? valid[406] :
                 (N1871)? valid[407] :
                 (N1873)? valid[408] :
                 (N1875)? valid[409] :
                 (N1877)? valid[410] :
                 (N1879)? valid[411] :
                 (N1881)? valid[412] :
                 (N1883)? valid[413] :
                 (N1885)? valid[414] :
                 (N1887)? valid[415] :
                 (N1889)? valid[416] :
                 (N1891)? valid[417] :
                 (N1893)? valid[418] :
                 (N1895)? valid[419] :
                 (N1897)? valid[420] :
                 (N1899)? valid[421] :
                 (N1901)? valid[422] :
                 (N1903)? valid[423] :
                 (N1905)? valid[424] :
                 (N1907)? valid[425] :
                 (N1909)? valid[426] :
                 (N1911)? valid[427] :
                 (N1913)? valid[428] :
                 (N1915)? valid[429] :
                 (N1917)? valid[430] :
                 (N1919)? valid[431] :
                 (N1921)? valid[432] :
                 (N1923)? valid[433] :
                 (N1925)? valid[434] :
                 (N1927)? valid[435] :
                 (N1929)? valid[436] :
                 (N1931)? valid[437] :
                 (N1933)? valid[438] :
                 (N1935)? valid[439] :
                 (N1937)? valid[440] :
                 (N1939)? valid[441] :
                 (N1941)? valid[442] :
                 (N1943)? valid[443] :
                 (N1945)? valid[444] :
                 (N1947)? valid[445] :
                 (N1949)? valid[446] :
                 (N1951)? valid[447] :
                 (N1953)? valid[448] :
                 (N1955)? valid[449] :
                 (N1957)? valid[450] :
                 (N1959)? valid[451] :
                 (N1961)? valid[452] :
                 (N1963)? valid[453] :
                 (N1965)? valid[454] :
                 (N1967)? valid[455] :
                 (N1969)? valid[456] :
                 (N1971)? valid[457] :
                 (N1973)? valid[458] :
                 (N1975)? valid[459] :
                 (N1977)? valid[460] :
                 (N1979)? valid[461] :
                 (N1981)? valid[462] :
                 (N1983)? valid[463] :
                 (N1985)? valid[464] :
                 (N1987)? valid[465] :
                 (N1989)? valid[466] :
                 (N1991)? valid[467] :
                 (N1993)? valid[468] :
                 (N1995)? valid[469] :
                 (N1997)? valid[470] :
                 (N1999)? valid[471] :
                 (N2001)? valid[472] :
                 (N2003)? valid[473] :
                 (N2005)? valid[474] :
                 (N2007)? valid[475] :
                 (N2009)? valid[476] :
                 (N2011)? valid[477] :
                 (N2013)? valid[478] :
                 (N2015)? valid[479] :
                 (N2017)? valid[480] :
                 (N2019)? valid[481] :
                 (N2021)? valid[482] :
                 (N2023)? valid[483] :
                 (N2025)? valid[484] :
                 (N2027)? valid[485] :
                 (N2029)? valid[486] :
                 (N2031)? valid[487] :
                 (N2033)? valid[488] :
                 (N2035)? valid[489] :
                 (N2037)? valid[490] :
                 (N2039)? valid[491] :
                 (N2041)? valid[492] :
                 (N2043)? valid[493] :
                 (N2045)? valid[494] :
                 (N2047)? valid[495] :
                 (N2049)? valid[496] :
                 (N2051)? valid[497] :
                 (N2053)? valid[498] :
                 (N2055)? valid[499] :
                 (N2057)? valid[500] :
                 (N2059)? valid[501] :
                 (N2061)? valid[502] :
                 (N2063)? valid[503] :
                 (N2065)? valid[504] :
                 (N2067)? valid[505] :
                 (N2069)? valid[506] :
                 (N2071)? valid[507] :
                 (N2073)? valid[508] :
                 (N2075)? valid[509] :
                 (N2077)? valid[510] :
                 (N2079)? valid[511] : 1'b0;

  bsg_mem_1rw_sync_width_p64_els_p512_addr_width_lp9
  btb_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(branch_target_i),
    .addr_i(addr),
    .v_i(n_0_net_),
    .w_i(w_v_i),
    .data_o(branch_target_o)
  );

  assign N2081 = idx_w_i[7] & idx_w_i[8];
  assign N2082 = N0 & idx_w_i[8];
  assign N0 = ~idx_w_i[7];
  assign N2083 = idx_w_i[7] & N1;
  assign N1 = ~idx_w_i[8];
  assign N2084 = N2 & N3;
  assign N2 = ~idx_w_i[7];
  assign N3 = ~idx_w_i[8];
  assign N2085 = idx_w_i[5] & idx_w_i[6];
  assign N2086 = N4 & idx_w_i[6];
  assign N4 = ~idx_w_i[5];
  assign N2087 = idx_w_i[5] & N5;
  assign N5 = ~idx_w_i[6];
  assign N2088 = N6 & N7;
  assign N6 = ~idx_w_i[5];
  assign N7 = ~idx_w_i[6];
  assign N2089 = N2081 & N2085;
  assign N2090 = N2081 & N2086;
  assign N2091 = N2081 & N2087;
  assign N2092 = N2081 & N2088;
  assign N2093 = N2082 & N2085;
  assign N2094 = N2082 & N2086;
  assign N2095 = N2082 & N2087;
  assign N2096 = N2082 & N2088;
  assign N2097 = N2083 & N2085;
  assign N2098 = N2083 & N2086;
  assign N2099 = N2083 & N2087;
  assign N2100 = N2083 & N2088;
  assign N2101 = N2084 & N2085;
  assign N2102 = N2084 & N2086;
  assign N2103 = N2084 & N2087;
  assign N2104 = N2084 & N2088;
  assign N2105 = idx_w_i[3] & idx_w_i[4];
  assign N2106 = N8 & idx_w_i[4];
  assign N8 = ~idx_w_i[3];
  assign N2107 = idx_w_i[3] & N9;
  assign N9 = ~idx_w_i[4];
  assign N2108 = N10 & N11;
  assign N10 = ~idx_w_i[3];
  assign N11 = ~idx_w_i[4];
  assign N2109 = ~idx_w_i[2];
  assign N2110 = idx_w_i[0] & idx_w_i[1];
  assign N2111 = N12 & idx_w_i[1];
  assign N12 = ~idx_w_i[0];
  assign N2112 = idx_w_i[0] & N13;
  assign N13 = ~idx_w_i[1];
  assign N2113 = N14 & N15;
  assign N14 = ~idx_w_i[0];
  assign N15 = ~idx_w_i[1];
  assign N2114 = idx_w_i[2] & N2110;
  assign N2115 = idx_w_i[2] & N2111;
  assign N2116 = idx_w_i[2] & N2112;
  assign N2117 = idx_w_i[2] & N2113;
  assign N2118 = N2109 & N2110;
  assign N2119 = N2109 & N2111;
  assign N2120 = N2109 & N2112;
  assign N2121 = N2109 & N2113;
  assign N2122 = N2105 & N2114;
  assign N2123 = N2105 & N2115;
  assign N2124 = N2105 & N2116;
  assign N2125 = N2105 & N2117;
  assign N2126 = N2105 & N2118;
  assign N2127 = N2105 & N2119;
  assign N2128 = N2105 & N2120;
  assign N2129 = N2105 & N2121;
  assign N2130 = N2106 & N2114;
  assign N2131 = N2106 & N2115;
  assign N2132 = N2106 & N2116;
  assign N2133 = N2106 & N2117;
  assign N2134 = N2106 & N2118;
  assign N2135 = N2106 & N2119;
  assign N2136 = N2106 & N2120;
  assign N2137 = N2106 & N2121;
  assign N2138 = N2107 & N2114;
  assign N2139 = N2107 & N2115;
  assign N2140 = N2107 & N2116;
  assign N2141 = N2107 & N2117;
  assign N2142 = N2107 & N2118;
  assign N2143 = N2107 & N2119;
  assign N2144 = N2107 & N2120;
  assign N2145 = N2107 & N2121;
  assign N2146 = N2108 & N2114;
  assign N2147 = N2108 & N2115;
  assign N2148 = N2108 & N2116;
  assign N2149 = N2108 & N2117;
  assign N2150 = N2108 & N2118;
  assign N2151 = N2108 & N2119;
  assign N2152 = N2108 & N2120;
  assign N2153 = N2108 & N2121;
  assign N534 = N2089 & N2122;
  assign N533 = N2089 & N2123;
  assign N532 = N2089 & N2124;
  assign N531 = N2089 & N2125;
  assign N530 = N2089 & N2126;
  assign N529 = N2089 & N2127;
  assign N528 = N2089 & N2128;
  assign N527 = N2089 & N2129;
  assign N526 = N2089 & N2130;
  assign N525 = N2089 & N2131;
  assign N524 = N2089 & N2132;
  assign N523 = N2089 & N2133;
  assign N522 = N2089 & N2134;
  assign N521 = N2089 & N2135;
  assign N520 = N2089 & N2136;
  assign N519 = N2089 & N2137;
  assign N518 = N2089 & N2138;
  assign N517 = N2089 & N2139;
  assign N516 = N2089 & N2140;
  assign N515 = N2089 & N2141;
  assign N514 = N2089 & N2142;
  assign N513 = N2089 & N2143;
  assign N512 = N2089 & N2144;
  assign N511 = N2089 & N2145;
  assign N510 = N2089 & N2146;
  assign N509 = N2089 & N2147;
  assign N508 = N2089 & N2148;
  assign N507 = N2089 & N2149;
  assign N506 = N2089 & N2150;
  assign N505 = N2089 & N2151;
  assign N504 = N2089 & N2152;
  assign N503 = N2089 & N2153;
  assign N502 = N2090 & N2122;
  assign N501 = N2090 & N2123;
  assign N500 = N2090 & N2124;
  assign N499 = N2090 & N2125;
  assign N498 = N2090 & N2126;
  assign N497 = N2090 & N2127;
  assign N496 = N2090 & N2128;
  assign N495 = N2090 & N2129;
  assign N494 = N2090 & N2130;
  assign N493 = N2090 & N2131;
  assign N492 = N2090 & N2132;
  assign N491 = N2090 & N2133;
  assign N490 = N2090 & N2134;
  assign N489 = N2090 & N2135;
  assign N488 = N2090 & N2136;
  assign N487 = N2090 & N2137;
  assign N486 = N2090 & N2138;
  assign N485 = N2090 & N2139;
  assign N484 = N2090 & N2140;
  assign N483 = N2090 & N2141;
  assign N482 = N2090 & N2142;
  assign N481 = N2090 & N2143;
  assign N480 = N2090 & N2144;
  assign N479 = N2090 & N2145;
  assign N478 = N2090 & N2146;
  assign N477 = N2090 & N2147;
  assign N476 = N2090 & N2148;
  assign N475 = N2090 & N2149;
  assign N474 = N2090 & N2150;
  assign N473 = N2090 & N2151;
  assign N472 = N2090 & N2152;
  assign N471 = N2090 & N2153;
  assign N470 = N2091 & N2122;
  assign N469 = N2091 & N2123;
  assign N468 = N2091 & N2124;
  assign N467 = N2091 & N2125;
  assign N466 = N2091 & N2126;
  assign N465 = N2091 & N2127;
  assign N464 = N2091 & N2128;
  assign N463 = N2091 & N2129;
  assign N462 = N2091 & N2130;
  assign N461 = N2091 & N2131;
  assign N460 = N2091 & N2132;
  assign N459 = N2091 & N2133;
  assign N458 = N2091 & N2134;
  assign N457 = N2091 & N2135;
  assign N456 = N2091 & N2136;
  assign N455 = N2091 & N2137;
  assign N454 = N2091 & N2138;
  assign N453 = N2091 & N2139;
  assign N452 = N2091 & N2140;
  assign N451 = N2091 & N2141;
  assign N450 = N2091 & N2142;
  assign N449 = N2091 & N2143;
  assign N448 = N2091 & N2144;
  assign N447 = N2091 & N2145;
  assign N446 = N2091 & N2146;
  assign N445 = N2091 & N2147;
  assign N444 = N2091 & N2148;
  assign N443 = N2091 & N2149;
  assign N442 = N2091 & N2150;
  assign N441 = N2091 & N2151;
  assign N440 = N2091 & N2152;
  assign N439 = N2091 & N2153;
  assign N438 = N2092 & N2122;
  assign N437 = N2092 & N2123;
  assign N436 = N2092 & N2124;
  assign N435 = N2092 & N2125;
  assign N434 = N2092 & N2126;
  assign N433 = N2092 & N2127;
  assign N432 = N2092 & N2128;
  assign N431 = N2092 & N2129;
  assign N430 = N2092 & N2130;
  assign N429 = N2092 & N2131;
  assign N428 = N2092 & N2132;
  assign N427 = N2092 & N2133;
  assign N426 = N2092 & N2134;
  assign N425 = N2092 & N2135;
  assign N424 = N2092 & N2136;
  assign N423 = N2092 & N2137;
  assign N422 = N2092 & N2138;
  assign N421 = N2092 & N2139;
  assign N420 = N2092 & N2140;
  assign N419 = N2092 & N2141;
  assign N418 = N2092 & N2142;
  assign N417 = N2092 & N2143;
  assign N416 = N2092 & N2144;
  assign N415 = N2092 & N2145;
  assign N414 = N2092 & N2146;
  assign N413 = N2092 & N2147;
  assign N412 = N2092 & N2148;
  assign N411 = N2092 & N2149;
  assign N410 = N2092 & N2150;
  assign N409 = N2092 & N2151;
  assign N408 = N2092 & N2152;
  assign N407 = N2092 & N2153;
  assign N406 = N2093 & N2122;
  assign N405 = N2093 & N2123;
  assign N404 = N2093 & N2124;
  assign N403 = N2093 & N2125;
  assign N402 = N2093 & N2126;
  assign N401 = N2093 & N2127;
  assign N400 = N2093 & N2128;
  assign N399 = N2093 & N2129;
  assign N398 = N2093 & N2130;
  assign N397 = N2093 & N2131;
  assign N396 = N2093 & N2132;
  assign N395 = N2093 & N2133;
  assign N394 = N2093 & N2134;
  assign N393 = N2093 & N2135;
  assign N392 = N2093 & N2136;
  assign N391 = N2093 & N2137;
  assign N390 = N2093 & N2138;
  assign N389 = N2093 & N2139;
  assign N388 = N2093 & N2140;
  assign N387 = N2093 & N2141;
  assign N386 = N2093 & N2142;
  assign N385 = N2093 & N2143;
  assign N384 = N2093 & N2144;
  assign N383 = N2093 & N2145;
  assign N382 = N2093 & N2146;
  assign N381 = N2093 & N2147;
  assign N380 = N2093 & N2148;
  assign N379 = N2093 & N2149;
  assign N378 = N2093 & N2150;
  assign N377 = N2093 & N2151;
  assign N376 = N2093 & N2152;
  assign N375 = N2093 & N2153;
  assign N374 = N2094 & N2122;
  assign N373 = N2094 & N2123;
  assign N372 = N2094 & N2124;
  assign N371 = N2094 & N2125;
  assign N370 = N2094 & N2126;
  assign N369 = N2094 & N2127;
  assign N368 = N2094 & N2128;
  assign N367 = N2094 & N2129;
  assign N366 = N2094 & N2130;
  assign N365 = N2094 & N2131;
  assign N364 = N2094 & N2132;
  assign N363 = N2094 & N2133;
  assign N362 = N2094 & N2134;
  assign N361 = N2094 & N2135;
  assign N360 = N2094 & N2136;
  assign N359 = N2094 & N2137;
  assign N358 = N2094 & N2138;
  assign N357 = N2094 & N2139;
  assign N356 = N2094 & N2140;
  assign N355 = N2094 & N2141;
  assign N354 = N2094 & N2142;
  assign N353 = N2094 & N2143;
  assign N352 = N2094 & N2144;
  assign N351 = N2094 & N2145;
  assign N350 = N2094 & N2146;
  assign N349 = N2094 & N2147;
  assign N348 = N2094 & N2148;
  assign N347 = N2094 & N2149;
  assign N346 = N2094 & N2150;
  assign N345 = N2094 & N2151;
  assign N344 = N2094 & N2152;
  assign N343 = N2094 & N2153;
  assign N342 = N2095 & N2122;
  assign N341 = N2095 & N2123;
  assign N340 = N2095 & N2124;
  assign N339 = N2095 & N2125;
  assign N338 = N2095 & N2126;
  assign N337 = N2095 & N2127;
  assign N336 = N2095 & N2128;
  assign N335 = N2095 & N2129;
  assign N334 = N2095 & N2130;
  assign N333 = N2095 & N2131;
  assign N332 = N2095 & N2132;
  assign N331 = N2095 & N2133;
  assign N330 = N2095 & N2134;
  assign N329 = N2095 & N2135;
  assign N328 = N2095 & N2136;
  assign N327 = N2095 & N2137;
  assign N326 = N2095 & N2138;
  assign N325 = N2095 & N2139;
  assign N324 = N2095 & N2140;
  assign N323 = N2095 & N2141;
  assign N322 = N2095 & N2142;
  assign N321 = N2095 & N2143;
  assign N320 = N2095 & N2144;
  assign N319 = N2095 & N2145;
  assign N318 = N2095 & N2146;
  assign N317 = N2095 & N2147;
  assign N316 = N2095 & N2148;
  assign N315 = N2095 & N2149;
  assign N314 = N2095 & N2150;
  assign N313 = N2095 & N2151;
  assign N312 = N2095 & N2152;
  assign N311 = N2095 & N2153;
  assign N310 = N2096 & N2122;
  assign N309 = N2096 & N2123;
  assign N308 = N2096 & N2124;
  assign N307 = N2096 & N2125;
  assign N306 = N2096 & N2126;
  assign N305 = N2096 & N2127;
  assign N304 = N2096 & N2128;
  assign N303 = N2096 & N2129;
  assign N302 = N2096 & N2130;
  assign N301 = N2096 & N2131;
  assign N300 = N2096 & N2132;
  assign N299 = N2096 & N2133;
  assign N298 = N2096 & N2134;
  assign N297 = N2096 & N2135;
  assign N296 = N2096 & N2136;
  assign N295 = N2096 & N2137;
  assign N294 = N2096 & N2138;
  assign N293 = N2096 & N2139;
  assign N292 = N2096 & N2140;
  assign N291 = N2096 & N2141;
  assign N290 = N2096 & N2142;
  assign N289 = N2096 & N2143;
  assign N288 = N2096 & N2144;
  assign N287 = N2096 & N2145;
  assign N286 = N2096 & N2146;
  assign N285 = N2096 & N2147;
  assign N284 = N2096 & N2148;
  assign N283 = N2096 & N2149;
  assign N282 = N2096 & N2150;
  assign N281 = N2096 & N2151;
  assign N280 = N2096 & N2152;
  assign N279 = N2096 & N2153;
  assign N278 = N2097 & N2122;
  assign N277 = N2097 & N2123;
  assign N276 = N2097 & N2124;
  assign N275 = N2097 & N2125;
  assign N274 = N2097 & N2126;
  assign N273 = N2097 & N2127;
  assign N272 = N2097 & N2128;
  assign N271 = N2097 & N2129;
  assign N270 = N2097 & N2130;
  assign N269 = N2097 & N2131;
  assign N268 = N2097 & N2132;
  assign N267 = N2097 & N2133;
  assign N266 = N2097 & N2134;
  assign N265 = N2097 & N2135;
  assign N264 = N2097 & N2136;
  assign N263 = N2097 & N2137;
  assign N262 = N2097 & N2138;
  assign N261 = N2097 & N2139;
  assign N260 = N2097 & N2140;
  assign N259 = N2097 & N2141;
  assign N258 = N2097 & N2142;
  assign N257 = N2097 & N2143;
  assign N256 = N2097 & N2144;
  assign N255 = N2097 & N2145;
  assign N254 = N2097 & N2146;
  assign N253 = N2097 & N2147;
  assign N252 = N2097 & N2148;
  assign N251 = N2097 & N2149;
  assign N250 = N2097 & N2150;
  assign N249 = N2097 & N2151;
  assign N248 = N2097 & N2152;
  assign N247 = N2097 & N2153;
  assign N246 = N2098 & N2122;
  assign N245 = N2098 & N2123;
  assign N244 = N2098 & N2124;
  assign N243 = N2098 & N2125;
  assign N242 = N2098 & N2126;
  assign N241 = N2098 & N2127;
  assign N240 = N2098 & N2128;
  assign N239 = N2098 & N2129;
  assign N238 = N2098 & N2130;
  assign N237 = N2098 & N2131;
  assign N236 = N2098 & N2132;
  assign N235 = N2098 & N2133;
  assign N234 = N2098 & N2134;
  assign N233 = N2098 & N2135;
  assign N232 = N2098 & N2136;
  assign N231 = N2098 & N2137;
  assign N230 = N2098 & N2138;
  assign N229 = N2098 & N2139;
  assign N228 = N2098 & N2140;
  assign N227 = N2098 & N2141;
  assign N226 = N2098 & N2142;
  assign N225 = N2098 & N2143;
  assign N224 = N2098 & N2144;
  assign N223 = N2098 & N2145;
  assign N222 = N2098 & N2146;
  assign N221 = N2098 & N2147;
  assign N220 = N2098 & N2148;
  assign N219 = N2098 & N2149;
  assign N218 = N2098 & N2150;
  assign N217 = N2098 & N2151;
  assign N216 = N2098 & N2152;
  assign N215 = N2098 & N2153;
  assign N214 = N2099 & N2122;
  assign N213 = N2099 & N2123;
  assign N212 = N2099 & N2124;
  assign N211 = N2099 & N2125;
  assign N210 = N2099 & N2126;
  assign N209 = N2099 & N2127;
  assign N208 = N2099 & N2128;
  assign N207 = N2099 & N2129;
  assign N206 = N2099 & N2130;
  assign N205 = N2099 & N2131;
  assign N204 = N2099 & N2132;
  assign N203 = N2099 & N2133;
  assign N202 = N2099 & N2134;
  assign N201 = N2099 & N2135;
  assign N200 = N2099 & N2136;
  assign N199 = N2099 & N2137;
  assign N198 = N2099 & N2138;
  assign N197 = N2099 & N2139;
  assign N196 = N2099 & N2140;
  assign N195 = N2099 & N2141;
  assign N194 = N2099 & N2142;
  assign N193 = N2099 & N2143;
  assign N192 = N2099 & N2144;
  assign N191 = N2099 & N2145;
  assign N190 = N2099 & N2146;
  assign N189 = N2099 & N2147;
  assign N188 = N2099 & N2148;
  assign N187 = N2099 & N2149;
  assign N186 = N2099 & N2150;
  assign N185 = N2099 & N2151;
  assign N184 = N2099 & N2152;
  assign N183 = N2099 & N2153;
  assign N182 = N2100 & N2122;
  assign N181 = N2100 & N2123;
  assign N180 = N2100 & N2124;
  assign N179 = N2100 & N2125;
  assign N178 = N2100 & N2126;
  assign N177 = N2100 & N2127;
  assign N176 = N2100 & N2128;
  assign N175 = N2100 & N2129;
  assign N174 = N2100 & N2130;
  assign N173 = N2100 & N2131;
  assign N172 = N2100 & N2132;
  assign N171 = N2100 & N2133;
  assign N170 = N2100 & N2134;
  assign N169 = N2100 & N2135;
  assign N168 = N2100 & N2136;
  assign N167 = N2100 & N2137;
  assign N166 = N2100 & N2138;
  assign N165 = N2100 & N2139;
  assign N164 = N2100 & N2140;
  assign N163 = N2100 & N2141;
  assign N162 = N2100 & N2142;
  assign N161 = N2100 & N2143;
  assign N160 = N2100 & N2144;
  assign N159 = N2100 & N2145;
  assign N158 = N2100 & N2146;
  assign N157 = N2100 & N2147;
  assign N156 = N2100 & N2148;
  assign N155 = N2100 & N2149;
  assign N154 = N2100 & N2150;
  assign N153 = N2100 & N2151;
  assign N152 = N2100 & N2152;
  assign N151 = N2100 & N2153;
  assign N150 = N2101 & N2122;
  assign N149 = N2101 & N2123;
  assign N148 = N2101 & N2124;
  assign N147 = N2101 & N2125;
  assign N146 = N2101 & N2126;
  assign N145 = N2101 & N2127;
  assign N144 = N2101 & N2128;
  assign N143 = N2101 & N2129;
  assign N142 = N2101 & N2130;
  assign N141 = N2101 & N2131;
  assign N140 = N2101 & N2132;
  assign N139 = N2101 & N2133;
  assign N138 = N2101 & N2134;
  assign N137 = N2101 & N2135;
  assign N136 = N2101 & N2136;
  assign N135 = N2101 & N2137;
  assign N134 = N2101 & N2138;
  assign N133 = N2101 & N2139;
  assign N132 = N2101 & N2140;
  assign N131 = N2101 & N2141;
  assign N130 = N2101 & N2142;
  assign N129 = N2101 & N2143;
  assign N128 = N2101 & N2144;
  assign N127 = N2101 & N2145;
  assign N126 = N2101 & N2146;
  assign N125 = N2101 & N2147;
  assign N124 = N2101 & N2148;
  assign N123 = N2101 & N2149;
  assign N122 = N2101 & N2150;
  assign N121 = N2101 & N2151;
  assign N120 = N2101 & N2152;
  assign N119 = N2101 & N2153;
  assign N118 = N2102 & N2122;
  assign N117 = N2102 & N2123;
  assign N116 = N2102 & N2124;
  assign N115 = N2102 & N2125;
  assign N114 = N2102 & N2126;
  assign N113 = N2102 & N2127;
  assign N112 = N2102 & N2128;
  assign N111 = N2102 & N2129;
  assign N110 = N2102 & N2130;
  assign N109 = N2102 & N2131;
  assign N108 = N2102 & N2132;
  assign N107 = N2102 & N2133;
  assign N106 = N2102 & N2134;
  assign N105 = N2102 & N2135;
  assign N104 = N2102 & N2136;
  assign N103 = N2102 & N2137;
  assign N102 = N2102 & N2138;
  assign N101 = N2102 & N2139;
  assign N100 = N2102 & N2140;
  assign N99 = N2102 & N2141;
  assign N98 = N2102 & N2142;
  assign N97 = N2102 & N2143;
  assign N96 = N2102 & N2144;
  assign N95 = N2102 & N2145;
  assign N94 = N2102 & N2146;
  assign N93 = N2102 & N2147;
  assign N92 = N2102 & N2148;
  assign N91 = N2102 & N2149;
  assign N90 = N2102 & N2150;
  assign N89 = N2102 & N2151;
  assign N88 = N2102 & N2152;
  assign N87 = N2102 & N2153;
  assign N86 = N2103 & N2122;
  assign N85 = N2103 & N2123;
  assign N84 = N2103 & N2124;
  assign N83 = N2103 & N2125;
  assign N82 = N2103 & N2126;
  assign N81 = N2103 & N2127;
  assign N80 = N2103 & N2128;
  assign N79 = N2103 & N2129;
  assign N78 = N2103 & N2130;
  assign N77 = N2103 & N2131;
  assign N76 = N2103 & N2132;
  assign N75 = N2103 & N2133;
  assign N74 = N2103 & N2134;
  assign N73 = N2103 & N2135;
  assign N72 = N2103 & N2136;
  assign N71 = N2103 & N2137;
  assign N70 = N2103 & N2138;
  assign N69 = N2103 & N2139;
  assign N68 = N2103 & N2140;
  assign N67 = N2103 & N2141;
  assign N66 = N2103 & N2142;
  assign N65 = N2103 & N2143;
  assign N64 = N2103 & N2144;
  assign N63 = N2103 & N2145;
  assign N62 = N2103 & N2146;
  assign N61 = N2103 & N2147;
  assign N60 = N2103 & N2148;
  assign N59 = N2103 & N2149;
  assign N58 = N2103 & N2150;
  assign N57 = N2103 & N2151;
  assign N56 = N2103 & N2152;
  assign N55 = N2103 & N2153;
  assign N54 = N2104 & N2122;
  assign N53 = N2104 & N2123;
  assign N52 = N2104 & N2124;
  assign N51 = N2104 & N2125;
  assign N50 = N2104 & N2126;
  assign N49 = N2104 & N2127;
  assign N48 = N2104 & N2128;
  assign N47 = N2104 & N2129;
  assign N46 = N2104 & N2130;
  assign N45 = N2104 & N2131;
  assign N44 = N2104 & N2132;
  assign N43 = N2104 & N2133;
  assign N42 = N2104 & N2134;
  assign N41 = N2104 & N2135;
  assign N40 = N2104 & N2136;
  assign N39 = N2104 & N2137;
  assign N38 = N2104 & N2138;
  assign N37 = N2104 & N2139;
  assign N36 = N2104 & N2140;
  assign N35 = N2104 & N2141;
  assign N34 = N2104 & N2142;
  assign N33 = N2104 & N2143;
  assign N32 = N2104 & N2144;
  assign N31 = N2104 & N2145;
  assign N30 = N2104 & N2146;
  assign N29 = N2104 & N2147;
  assign N28 = N2104 & N2148;
  assign N27 = N2104 & N2149;
  assign N26 = N2104 & N2150;
  assign N25 = N2104 & N2151;
  assign N24 = N2104 & N2152;
  assign N23 = N2104 & N2153;
  assign { N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N540, N539, N538, N537, N536, N535 } = (N16)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N541)? { N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23 } :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = N19;
  assign addr = (N17)? idx_w_i :
                (N18)? idx_r_i : 1'b0;
  assign N17 = N1050;
  assign N18 = N1049;
  assign N19 = reset_i;
  assign N20 = w_v_i;
  assign N21 = N20 | N19;
  assign N22 = ~N21;
  assign N1048 = ~N19;
  assign N541 = N20 & N1048;
  assign N1049 = ~w_v_i;
  assign N1050 = w_v_i;
  assign N1051 = ~idx_r_i[0];
  assign N1052 = ~idx_r_i[1];
  assign N1053 = N1051 & N1052;
  assign N1054 = N1051 & idx_r_i[1];
  assign N1055 = idx_r_i[0] & N1052;
  assign N1056 = idx_r_i[0] & idx_r_i[1];
  assign N1057 = ~idx_r_i[2];
  assign N1058 = N1053 & N1057;
  assign N1059 = N1053 & idx_r_i[2];
  assign N1060 = N1055 & N1057;
  assign N1061 = N1055 & idx_r_i[2];
  assign N1062 = N1054 & N1057;
  assign N1063 = N1054 & idx_r_i[2];
  assign N1064 = N1056 & N1057;
  assign N1065 = N1056 & idx_r_i[2];
  assign N1066 = ~idx_r_i[3];
  assign N1067 = N1058 & N1066;
  assign N1068 = N1058 & idx_r_i[3];
  assign N1069 = N1060 & N1066;
  assign N1070 = N1060 & idx_r_i[3];
  assign N1071 = N1062 & N1066;
  assign N1072 = N1062 & idx_r_i[3];
  assign N1073 = N1064 & N1066;
  assign N1074 = N1064 & idx_r_i[3];
  assign N1075 = N1059 & N1066;
  assign N1076 = N1059 & idx_r_i[3];
  assign N1077 = N1061 & N1066;
  assign N1078 = N1061 & idx_r_i[3];
  assign N1079 = N1063 & N1066;
  assign N1080 = N1063 & idx_r_i[3];
  assign N1081 = N1065 & N1066;
  assign N1082 = N1065 & idx_r_i[3];
  assign N1083 = ~idx_r_i[4];
  assign N1084 = N1067 & N1083;
  assign N1085 = N1067 & idx_r_i[4];
  assign N1086 = N1069 & N1083;
  assign N1087 = N1069 & idx_r_i[4];
  assign N1088 = N1071 & N1083;
  assign N1089 = N1071 & idx_r_i[4];
  assign N1090 = N1073 & N1083;
  assign N1091 = N1073 & idx_r_i[4];
  assign N1092 = N1075 & N1083;
  assign N1093 = N1075 & idx_r_i[4];
  assign N1094 = N1077 & N1083;
  assign N1095 = N1077 & idx_r_i[4];
  assign N1096 = N1079 & N1083;
  assign N1097 = N1079 & idx_r_i[4];
  assign N1098 = N1081 & N1083;
  assign N1099 = N1081 & idx_r_i[4];
  assign N1100 = N1068 & N1083;
  assign N1101 = N1068 & idx_r_i[4];
  assign N1102 = N1070 & N1083;
  assign N1103 = N1070 & idx_r_i[4];
  assign N1104 = N1072 & N1083;
  assign N1105 = N1072 & idx_r_i[4];
  assign N1106 = N1074 & N1083;
  assign N1107 = N1074 & idx_r_i[4];
  assign N1108 = N1076 & N1083;
  assign N1109 = N1076 & idx_r_i[4];
  assign N1110 = N1078 & N1083;
  assign N1111 = N1078 & idx_r_i[4];
  assign N1112 = N1080 & N1083;
  assign N1113 = N1080 & idx_r_i[4];
  assign N1114 = N1082 & N1083;
  assign N1115 = N1082 & idx_r_i[4];
  assign N1116 = ~idx_r_i[5];
  assign N1117 = N1084 & N1116;
  assign N1118 = N1084 & idx_r_i[5];
  assign N1119 = N1086 & N1116;
  assign N1120 = N1086 & idx_r_i[5];
  assign N1121 = N1088 & N1116;
  assign N1122 = N1088 & idx_r_i[5];
  assign N1123 = N1090 & N1116;
  assign N1124 = N1090 & idx_r_i[5];
  assign N1125 = N1092 & N1116;
  assign N1126 = N1092 & idx_r_i[5];
  assign N1127 = N1094 & N1116;
  assign N1128 = N1094 & idx_r_i[5];
  assign N1129 = N1096 & N1116;
  assign N1130 = N1096 & idx_r_i[5];
  assign N1131 = N1098 & N1116;
  assign N1132 = N1098 & idx_r_i[5];
  assign N1133 = N1100 & N1116;
  assign N1134 = N1100 & idx_r_i[5];
  assign N1135 = N1102 & N1116;
  assign N1136 = N1102 & idx_r_i[5];
  assign N1137 = N1104 & N1116;
  assign N1138 = N1104 & idx_r_i[5];
  assign N1139 = N1106 & N1116;
  assign N1140 = N1106 & idx_r_i[5];
  assign N1141 = N1108 & N1116;
  assign N1142 = N1108 & idx_r_i[5];
  assign N1143 = N1110 & N1116;
  assign N1144 = N1110 & idx_r_i[5];
  assign N1145 = N1112 & N1116;
  assign N1146 = N1112 & idx_r_i[5];
  assign N1147 = N1114 & N1116;
  assign N1148 = N1114 & idx_r_i[5];
  assign N1149 = N1085 & N1116;
  assign N1150 = N1085 & idx_r_i[5];
  assign N1151 = N1087 & N1116;
  assign N1152 = N1087 & idx_r_i[5];
  assign N1153 = N1089 & N1116;
  assign N1154 = N1089 & idx_r_i[5];
  assign N1155 = N1091 & N1116;
  assign N1156 = N1091 & idx_r_i[5];
  assign N1157 = N1093 & N1116;
  assign N1158 = N1093 & idx_r_i[5];
  assign N1159 = N1095 & N1116;
  assign N1160 = N1095 & idx_r_i[5];
  assign N1161 = N1097 & N1116;
  assign N1162 = N1097 & idx_r_i[5];
  assign N1163 = N1099 & N1116;
  assign N1164 = N1099 & idx_r_i[5];
  assign N1165 = N1101 & N1116;
  assign N1166 = N1101 & idx_r_i[5];
  assign N1167 = N1103 & N1116;
  assign N1168 = N1103 & idx_r_i[5];
  assign N1169 = N1105 & N1116;
  assign N1170 = N1105 & idx_r_i[5];
  assign N1171 = N1107 & N1116;
  assign N1172 = N1107 & idx_r_i[5];
  assign N1173 = N1109 & N1116;
  assign N1174 = N1109 & idx_r_i[5];
  assign N1175 = N1111 & N1116;
  assign N1176 = N1111 & idx_r_i[5];
  assign N1177 = N1113 & N1116;
  assign N1178 = N1113 & idx_r_i[5];
  assign N1179 = N1115 & N1116;
  assign N1180 = N1115 & idx_r_i[5];
  assign N1181 = ~idx_r_i[6];
  assign N1182 = N1117 & N1181;
  assign N1183 = N1117 & idx_r_i[6];
  assign N1184 = N1119 & N1181;
  assign N1185 = N1119 & idx_r_i[6];
  assign N1186 = N1121 & N1181;
  assign N1187 = N1121 & idx_r_i[6];
  assign N1188 = N1123 & N1181;
  assign N1189 = N1123 & idx_r_i[6];
  assign N1190 = N1125 & N1181;
  assign N1191 = N1125 & idx_r_i[6];
  assign N1192 = N1127 & N1181;
  assign N1193 = N1127 & idx_r_i[6];
  assign N1194 = N1129 & N1181;
  assign N1195 = N1129 & idx_r_i[6];
  assign N1196 = N1131 & N1181;
  assign N1197 = N1131 & idx_r_i[6];
  assign N1198 = N1133 & N1181;
  assign N1199 = N1133 & idx_r_i[6];
  assign N1200 = N1135 & N1181;
  assign N1201 = N1135 & idx_r_i[6];
  assign N1202 = N1137 & N1181;
  assign N1203 = N1137 & idx_r_i[6];
  assign N1204 = N1139 & N1181;
  assign N1205 = N1139 & idx_r_i[6];
  assign N1206 = N1141 & N1181;
  assign N1207 = N1141 & idx_r_i[6];
  assign N1208 = N1143 & N1181;
  assign N1209 = N1143 & idx_r_i[6];
  assign N1210 = N1145 & N1181;
  assign N1211 = N1145 & idx_r_i[6];
  assign N1212 = N1147 & N1181;
  assign N1213 = N1147 & idx_r_i[6];
  assign N1214 = N1149 & N1181;
  assign N1215 = N1149 & idx_r_i[6];
  assign N1216 = N1151 & N1181;
  assign N1217 = N1151 & idx_r_i[6];
  assign N1218 = N1153 & N1181;
  assign N1219 = N1153 & idx_r_i[6];
  assign N1220 = N1155 & N1181;
  assign N1221 = N1155 & idx_r_i[6];
  assign N1222 = N1157 & N1181;
  assign N1223 = N1157 & idx_r_i[6];
  assign N1224 = N1159 & N1181;
  assign N1225 = N1159 & idx_r_i[6];
  assign N1226 = N1161 & N1181;
  assign N1227 = N1161 & idx_r_i[6];
  assign N1228 = N1163 & N1181;
  assign N1229 = N1163 & idx_r_i[6];
  assign N1230 = N1165 & N1181;
  assign N1231 = N1165 & idx_r_i[6];
  assign N1232 = N1167 & N1181;
  assign N1233 = N1167 & idx_r_i[6];
  assign N1234 = N1169 & N1181;
  assign N1235 = N1169 & idx_r_i[6];
  assign N1236 = N1171 & N1181;
  assign N1237 = N1171 & idx_r_i[6];
  assign N1238 = N1173 & N1181;
  assign N1239 = N1173 & idx_r_i[6];
  assign N1240 = N1175 & N1181;
  assign N1241 = N1175 & idx_r_i[6];
  assign N1242 = N1177 & N1181;
  assign N1243 = N1177 & idx_r_i[6];
  assign N1244 = N1179 & N1181;
  assign N1245 = N1179 & idx_r_i[6];
  assign N1246 = N1118 & N1181;
  assign N1247 = N1118 & idx_r_i[6];
  assign N1248 = N1120 & N1181;
  assign N1249 = N1120 & idx_r_i[6];
  assign N1250 = N1122 & N1181;
  assign N1251 = N1122 & idx_r_i[6];
  assign N1252 = N1124 & N1181;
  assign N1253 = N1124 & idx_r_i[6];
  assign N1254 = N1126 & N1181;
  assign N1255 = N1126 & idx_r_i[6];
  assign N1256 = N1128 & N1181;
  assign N1257 = N1128 & idx_r_i[6];
  assign N1258 = N1130 & N1181;
  assign N1259 = N1130 & idx_r_i[6];
  assign N1260 = N1132 & N1181;
  assign N1261 = N1132 & idx_r_i[6];
  assign N1262 = N1134 & N1181;
  assign N1263 = N1134 & idx_r_i[6];
  assign N1264 = N1136 & N1181;
  assign N1265 = N1136 & idx_r_i[6];
  assign N1266 = N1138 & N1181;
  assign N1267 = N1138 & idx_r_i[6];
  assign N1268 = N1140 & N1181;
  assign N1269 = N1140 & idx_r_i[6];
  assign N1270 = N1142 & N1181;
  assign N1271 = N1142 & idx_r_i[6];
  assign N1272 = N1144 & N1181;
  assign N1273 = N1144 & idx_r_i[6];
  assign N1274 = N1146 & N1181;
  assign N1275 = N1146 & idx_r_i[6];
  assign N1276 = N1148 & N1181;
  assign N1277 = N1148 & idx_r_i[6];
  assign N1278 = N1150 & N1181;
  assign N1279 = N1150 & idx_r_i[6];
  assign N1280 = N1152 & N1181;
  assign N1281 = N1152 & idx_r_i[6];
  assign N1282 = N1154 & N1181;
  assign N1283 = N1154 & idx_r_i[6];
  assign N1284 = N1156 & N1181;
  assign N1285 = N1156 & idx_r_i[6];
  assign N1286 = N1158 & N1181;
  assign N1287 = N1158 & idx_r_i[6];
  assign N1288 = N1160 & N1181;
  assign N1289 = N1160 & idx_r_i[6];
  assign N1290 = N1162 & N1181;
  assign N1291 = N1162 & idx_r_i[6];
  assign N1292 = N1164 & N1181;
  assign N1293 = N1164 & idx_r_i[6];
  assign N1294 = N1166 & N1181;
  assign N1295 = N1166 & idx_r_i[6];
  assign N1296 = N1168 & N1181;
  assign N1297 = N1168 & idx_r_i[6];
  assign N1298 = N1170 & N1181;
  assign N1299 = N1170 & idx_r_i[6];
  assign N1300 = N1172 & N1181;
  assign N1301 = N1172 & idx_r_i[6];
  assign N1302 = N1174 & N1181;
  assign N1303 = N1174 & idx_r_i[6];
  assign N1304 = N1176 & N1181;
  assign N1305 = N1176 & idx_r_i[6];
  assign N1306 = N1178 & N1181;
  assign N1307 = N1178 & idx_r_i[6];
  assign N1308 = N1180 & N1181;
  assign N1309 = N1180 & idx_r_i[6];
  assign N1310 = ~idx_r_i[7];
  assign N1311 = N1182 & N1310;
  assign N1312 = N1182 & idx_r_i[7];
  assign N1313 = N1184 & N1310;
  assign N1314 = N1184 & idx_r_i[7];
  assign N1315 = N1186 & N1310;
  assign N1316 = N1186 & idx_r_i[7];
  assign N1317 = N1188 & N1310;
  assign N1318 = N1188 & idx_r_i[7];
  assign N1319 = N1190 & N1310;
  assign N1320 = N1190 & idx_r_i[7];
  assign N1321 = N1192 & N1310;
  assign N1322 = N1192 & idx_r_i[7];
  assign N1323 = N1194 & N1310;
  assign N1324 = N1194 & idx_r_i[7];
  assign N1325 = N1196 & N1310;
  assign N1326 = N1196 & idx_r_i[7];
  assign N1327 = N1198 & N1310;
  assign N1328 = N1198 & idx_r_i[7];
  assign N1329 = N1200 & N1310;
  assign N1330 = N1200 & idx_r_i[7];
  assign N1331 = N1202 & N1310;
  assign N1332 = N1202 & idx_r_i[7];
  assign N1333 = N1204 & N1310;
  assign N1334 = N1204 & idx_r_i[7];
  assign N1335 = N1206 & N1310;
  assign N1336 = N1206 & idx_r_i[7];
  assign N1337 = N1208 & N1310;
  assign N1338 = N1208 & idx_r_i[7];
  assign N1339 = N1210 & N1310;
  assign N1340 = N1210 & idx_r_i[7];
  assign N1341 = N1212 & N1310;
  assign N1342 = N1212 & idx_r_i[7];
  assign N1343 = N1214 & N1310;
  assign N1344 = N1214 & idx_r_i[7];
  assign N1345 = N1216 & N1310;
  assign N1346 = N1216 & idx_r_i[7];
  assign N1347 = N1218 & N1310;
  assign N1348 = N1218 & idx_r_i[7];
  assign N1349 = N1220 & N1310;
  assign N1350 = N1220 & idx_r_i[7];
  assign N1351 = N1222 & N1310;
  assign N1352 = N1222 & idx_r_i[7];
  assign N1353 = N1224 & N1310;
  assign N1354 = N1224 & idx_r_i[7];
  assign N1355 = N1226 & N1310;
  assign N1356 = N1226 & idx_r_i[7];
  assign N1357 = N1228 & N1310;
  assign N1358 = N1228 & idx_r_i[7];
  assign N1359 = N1230 & N1310;
  assign N1360 = N1230 & idx_r_i[7];
  assign N1361 = N1232 & N1310;
  assign N1362 = N1232 & idx_r_i[7];
  assign N1363 = N1234 & N1310;
  assign N1364 = N1234 & idx_r_i[7];
  assign N1365 = N1236 & N1310;
  assign N1366 = N1236 & idx_r_i[7];
  assign N1367 = N1238 & N1310;
  assign N1368 = N1238 & idx_r_i[7];
  assign N1369 = N1240 & N1310;
  assign N1370 = N1240 & idx_r_i[7];
  assign N1371 = N1242 & N1310;
  assign N1372 = N1242 & idx_r_i[7];
  assign N1373 = N1244 & N1310;
  assign N1374 = N1244 & idx_r_i[7];
  assign N1375 = N1246 & N1310;
  assign N1376 = N1246 & idx_r_i[7];
  assign N1377 = N1248 & N1310;
  assign N1378 = N1248 & idx_r_i[7];
  assign N1379 = N1250 & N1310;
  assign N1380 = N1250 & idx_r_i[7];
  assign N1381 = N1252 & N1310;
  assign N1382 = N1252 & idx_r_i[7];
  assign N1383 = N1254 & N1310;
  assign N1384 = N1254 & idx_r_i[7];
  assign N1385 = N1256 & N1310;
  assign N1386 = N1256 & idx_r_i[7];
  assign N1387 = N1258 & N1310;
  assign N1388 = N1258 & idx_r_i[7];
  assign N1389 = N1260 & N1310;
  assign N1390 = N1260 & idx_r_i[7];
  assign N1391 = N1262 & N1310;
  assign N1392 = N1262 & idx_r_i[7];
  assign N1393 = N1264 & N1310;
  assign N1394 = N1264 & idx_r_i[7];
  assign N1395 = N1266 & N1310;
  assign N1396 = N1266 & idx_r_i[7];
  assign N1397 = N1268 & N1310;
  assign N1398 = N1268 & idx_r_i[7];
  assign N1399 = N1270 & N1310;
  assign N1400 = N1270 & idx_r_i[7];
  assign N1401 = N1272 & N1310;
  assign N1402 = N1272 & idx_r_i[7];
  assign N1403 = N1274 & N1310;
  assign N1404 = N1274 & idx_r_i[7];
  assign N1405 = N1276 & N1310;
  assign N1406 = N1276 & idx_r_i[7];
  assign N1407 = N1278 & N1310;
  assign N1408 = N1278 & idx_r_i[7];
  assign N1409 = N1280 & N1310;
  assign N1410 = N1280 & idx_r_i[7];
  assign N1411 = N1282 & N1310;
  assign N1412 = N1282 & idx_r_i[7];
  assign N1413 = N1284 & N1310;
  assign N1414 = N1284 & idx_r_i[7];
  assign N1415 = N1286 & N1310;
  assign N1416 = N1286 & idx_r_i[7];
  assign N1417 = N1288 & N1310;
  assign N1418 = N1288 & idx_r_i[7];
  assign N1419 = N1290 & N1310;
  assign N1420 = N1290 & idx_r_i[7];
  assign N1421 = N1292 & N1310;
  assign N1422 = N1292 & idx_r_i[7];
  assign N1423 = N1294 & N1310;
  assign N1424 = N1294 & idx_r_i[7];
  assign N1425 = N1296 & N1310;
  assign N1426 = N1296 & idx_r_i[7];
  assign N1427 = N1298 & N1310;
  assign N1428 = N1298 & idx_r_i[7];
  assign N1429 = N1300 & N1310;
  assign N1430 = N1300 & idx_r_i[7];
  assign N1431 = N1302 & N1310;
  assign N1432 = N1302 & idx_r_i[7];
  assign N1433 = N1304 & N1310;
  assign N1434 = N1304 & idx_r_i[7];
  assign N1435 = N1306 & N1310;
  assign N1436 = N1306 & idx_r_i[7];
  assign N1437 = N1308 & N1310;
  assign N1438 = N1308 & idx_r_i[7];
  assign N1439 = N1183 & N1310;
  assign N1440 = N1183 & idx_r_i[7];
  assign N1441 = N1185 & N1310;
  assign N1442 = N1185 & idx_r_i[7];
  assign N1443 = N1187 & N1310;
  assign N1444 = N1187 & idx_r_i[7];
  assign N1445 = N1189 & N1310;
  assign N1446 = N1189 & idx_r_i[7];
  assign N1447 = N1191 & N1310;
  assign N1448 = N1191 & idx_r_i[7];
  assign N1449 = N1193 & N1310;
  assign N1450 = N1193 & idx_r_i[7];
  assign N1451 = N1195 & N1310;
  assign N1452 = N1195 & idx_r_i[7];
  assign N1453 = N1197 & N1310;
  assign N1454 = N1197 & idx_r_i[7];
  assign N1455 = N1199 & N1310;
  assign N1456 = N1199 & idx_r_i[7];
  assign N1457 = N1201 & N1310;
  assign N1458 = N1201 & idx_r_i[7];
  assign N1459 = N1203 & N1310;
  assign N1460 = N1203 & idx_r_i[7];
  assign N1461 = N1205 & N1310;
  assign N1462 = N1205 & idx_r_i[7];
  assign N1463 = N1207 & N1310;
  assign N1464 = N1207 & idx_r_i[7];
  assign N1465 = N1209 & N1310;
  assign N1466 = N1209 & idx_r_i[7];
  assign N1467 = N1211 & N1310;
  assign N1468 = N1211 & idx_r_i[7];
  assign N1469 = N1213 & N1310;
  assign N1470 = N1213 & idx_r_i[7];
  assign N1471 = N1215 & N1310;
  assign N1472 = N1215 & idx_r_i[7];
  assign N1473 = N1217 & N1310;
  assign N1474 = N1217 & idx_r_i[7];
  assign N1475 = N1219 & N1310;
  assign N1476 = N1219 & idx_r_i[7];
  assign N1477 = N1221 & N1310;
  assign N1478 = N1221 & idx_r_i[7];
  assign N1479 = N1223 & N1310;
  assign N1480 = N1223 & idx_r_i[7];
  assign N1481 = N1225 & N1310;
  assign N1482 = N1225 & idx_r_i[7];
  assign N1483 = N1227 & N1310;
  assign N1484 = N1227 & idx_r_i[7];
  assign N1485 = N1229 & N1310;
  assign N1486 = N1229 & idx_r_i[7];
  assign N1487 = N1231 & N1310;
  assign N1488 = N1231 & idx_r_i[7];
  assign N1489 = N1233 & N1310;
  assign N1490 = N1233 & idx_r_i[7];
  assign N1491 = N1235 & N1310;
  assign N1492 = N1235 & idx_r_i[7];
  assign N1493 = N1237 & N1310;
  assign N1494 = N1237 & idx_r_i[7];
  assign N1495 = N1239 & N1310;
  assign N1496 = N1239 & idx_r_i[7];
  assign N1497 = N1241 & N1310;
  assign N1498 = N1241 & idx_r_i[7];
  assign N1499 = N1243 & N1310;
  assign N1500 = N1243 & idx_r_i[7];
  assign N1501 = N1245 & N1310;
  assign N1502 = N1245 & idx_r_i[7];
  assign N1503 = N1247 & N1310;
  assign N1504 = N1247 & idx_r_i[7];
  assign N1505 = N1249 & N1310;
  assign N1506 = N1249 & idx_r_i[7];
  assign N1507 = N1251 & N1310;
  assign N1508 = N1251 & idx_r_i[7];
  assign N1509 = N1253 & N1310;
  assign N1510 = N1253 & idx_r_i[7];
  assign N1511 = N1255 & N1310;
  assign N1512 = N1255 & idx_r_i[7];
  assign N1513 = N1257 & N1310;
  assign N1514 = N1257 & idx_r_i[7];
  assign N1515 = N1259 & N1310;
  assign N1516 = N1259 & idx_r_i[7];
  assign N1517 = N1261 & N1310;
  assign N1518 = N1261 & idx_r_i[7];
  assign N1519 = N1263 & N1310;
  assign N1520 = N1263 & idx_r_i[7];
  assign N1521 = N1265 & N1310;
  assign N1522 = N1265 & idx_r_i[7];
  assign N1523 = N1267 & N1310;
  assign N1524 = N1267 & idx_r_i[7];
  assign N1525 = N1269 & N1310;
  assign N1526 = N1269 & idx_r_i[7];
  assign N1527 = N1271 & N1310;
  assign N1528 = N1271 & idx_r_i[7];
  assign N1529 = N1273 & N1310;
  assign N1530 = N1273 & idx_r_i[7];
  assign N1531 = N1275 & N1310;
  assign N1532 = N1275 & idx_r_i[7];
  assign N1533 = N1277 & N1310;
  assign N1534 = N1277 & idx_r_i[7];
  assign N1535 = N1279 & N1310;
  assign N1536 = N1279 & idx_r_i[7];
  assign N1537 = N1281 & N1310;
  assign N1538 = N1281 & idx_r_i[7];
  assign N1539 = N1283 & N1310;
  assign N1540 = N1283 & idx_r_i[7];
  assign N1541 = N1285 & N1310;
  assign N1542 = N1285 & idx_r_i[7];
  assign N1543 = N1287 & N1310;
  assign N1544 = N1287 & idx_r_i[7];
  assign N1545 = N1289 & N1310;
  assign N1546 = N1289 & idx_r_i[7];
  assign N1547 = N1291 & N1310;
  assign N1548 = N1291 & idx_r_i[7];
  assign N1549 = N1293 & N1310;
  assign N1550 = N1293 & idx_r_i[7];
  assign N1551 = N1295 & N1310;
  assign N1552 = N1295 & idx_r_i[7];
  assign N1553 = N1297 & N1310;
  assign N1554 = N1297 & idx_r_i[7];
  assign N1555 = N1299 & N1310;
  assign N1556 = N1299 & idx_r_i[7];
  assign N1557 = N1301 & N1310;
  assign N1558 = N1301 & idx_r_i[7];
  assign N1559 = N1303 & N1310;
  assign N1560 = N1303 & idx_r_i[7];
  assign N1561 = N1305 & N1310;
  assign N1562 = N1305 & idx_r_i[7];
  assign N1563 = N1307 & N1310;
  assign N1564 = N1307 & idx_r_i[7];
  assign N1565 = N1309 & N1310;
  assign N1566 = N1309 & idx_r_i[7];
  assign N1567 = ~idx_r_i[8];
  assign N1568 = N1311 & N1567;
  assign N1569 = N1311 & idx_r_i[8];
  assign N1570 = N1313 & N1567;
  assign N1571 = N1313 & idx_r_i[8];
  assign N1572 = N1315 & N1567;
  assign N1573 = N1315 & idx_r_i[8];
  assign N1574 = N1317 & N1567;
  assign N1575 = N1317 & idx_r_i[8];
  assign N1576 = N1319 & N1567;
  assign N1577 = N1319 & idx_r_i[8];
  assign N1578 = N1321 & N1567;
  assign N1579 = N1321 & idx_r_i[8];
  assign N1580 = N1323 & N1567;
  assign N1581 = N1323 & idx_r_i[8];
  assign N1582 = N1325 & N1567;
  assign N1583 = N1325 & idx_r_i[8];
  assign N1584 = N1327 & N1567;
  assign N1585 = N1327 & idx_r_i[8];
  assign N1586 = N1329 & N1567;
  assign N1587 = N1329 & idx_r_i[8];
  assign N1588 = N1331 & N1567;
  assign N1589 = N1331 & idx_r_i[8];
  assign N1590 = N1333 & N1567;
  assign N1591 = N1333 & idx_r_i[8];
  assign N1592 = N1335 & N1567;
  assign N1593 = N1335 & idx_r_i[8];
  assign N1594 = N1337 & N1567;
  assign N1595 = N1337 & idx_r_i[8];
  assign N1596 = N1339 & N1567;
  assign N1597 = N1339 & idx_r_i[8];
  assign N1598 = N1341 & N1567;
  assign N1599 = N1341 & idx_r_i[8];
  assign N1600 = N1343 & N1567;
  assign N1601 = N1343 & idx_r_i[8];
  assign N1602 = N1345 & N1567;
  assign N1603 = N1345 & idx_r_i[8];
  assign N1604 = N1347 & N1567;
  assign N1605 = N1347 & idx_r_i[8];
  assign N1606 = N1349 & N1567;
  assign N1607 = N1349 & idx_r_i[8];
  assign N1608 = N1351 & N1567;
  assign N1609 = N1351 & idx_r_i[8];
  assign N1610 = N1353 & N1567;
  assign N1611 = N1353 & idx_r_i[8];
  assign N1612 = N1355 & N1567;
  assign N1613 = N1355 & idx_r_i[8];
  assign N1614 = N1357 & N1567;
  assign N1615 = N1357 & idx_r_i[8];
  assign N1616 = N1359 & N1567;
  assign N1617 = N1359 & idx_r_i[8];
  assign N1618 = N1361 & N1567;
  assign N1619 = N1361 & idx_r_i[8];
  assign N1620 = N1363 & N1567;
  assign N1621 = N1363 & idx_r_i[8];
  assign N1622 = N1365 & N1567;
  assign N1623 = N1365 & idx_r_i[8];
  assign N1624 = N1367 & N1567;
  assign N1625 = N1367 & idx_r_i[8];
  assign N1626 = N1369 & N1567;
  assign N1627 = N1369 & idx_r_i[8];
  assign N1628 = N1371 & N1567;
  assign N1629 = N1371 & idx_r_i[8];
  assign N1630 = N1373 & N1567;
  assign N1631 = N1373 & idx_r_i[8];
  assign N1632 = N1375 & N1567;
  assign N1633 = N1375 & idx_r_i[8];
  assign N1634 = N1377 & N1567;
  assign N1635 = N1377 & idx_r_i[8];
  assign N1636 = N1379 & N1567;
  assign N1637 = N1379 & idx_r_i[8];
  assign N1638 = N1381 & N1567;
  assign N1639 = N1381 & idx_r_i[8];
  assign N1640 = N1383 & N1567;
  assign N1641 = N1383 & idx_r_i[8];
  assign N1642 = N1385 & N1567;
  assign N1643 = N1385 & idx_r_i[8];
  assign N1644 = N1387 & N1567;
  assign N1645 = N1387 & idx_r_i[8];
  assign N1646 = N1389 & N1567;
  assign N1647 = N1389 & idx_r_i[8];
  assign N1648 = N1391 & N1567;
  assign N1649 = N1391 & idx_r_i[8];
  assign N1650 = N1393 & N1567;
  assign N1651 = N1393 & idx_r_i[8];
  assign N1652 = N1395 & N1567;
  assign N1653 = N1395 & idx_r_i[8];
  assign N1654 = N1397 & N1567;
  assign N1655 = N1397 & idx_r_i[8];
  assign N1656 = N1399 & N1567;
  assign N1657 = N1399 & idx_r_i[8];
  assign N1658 = N1401 & N1567;
  assign N1659 = N1401 & idx_r_i[8];
  assign N1660 = N1403 & N1567;
  assign N1661 = N1403 & idx_r_i[8];
  assign N1662 = N1405 & N1567;
  assign N1663 = N1405 & idx_r_i[8];
  assign N1664 = N1407 & N1567;
  assign N1665 = N1407 & idx_r_i[8];
  assign N1666 = N1409 & N1567;
  assign N1667 = N1409 & idx_r_i[8];
  assign N1668 = N1411 & N1567;
  assign N1669 = N1411 & idx_r_i[8];
  assign N1670 = N1413 & N1567;
  assign N1671 = N1413 & idx_r_i[8];
  assign N1672 = N1415 & N1567;
  assign N1673 = N1415 & idx_r_i[8];
  assign N1674 = N1417 & N1567;
  assign N1675 = N1417 & idx_r_i[8];
  assign N1676 = N1419 & N1567;
  assign N1677 = N1419 & idx_r_i[8];
  assign N1678 = N1421 & N1567;
  assign N1679 = N1421 & idx_r_i[8];
  assign N1680 = N1423 & N1567;
  assign N1681 = N1423 & idx_r_i[8];
  assign N1682 = N1425 & N1567;
  assign N1683 = N1425 & idx_r_i[8];
  assign N1684 = N1427 & N1567;
  assign N1685 = N1427 & idx_r_i[8];
  assign N1686 = N1429 & N1567;
  assign N1687 = N1429 & idx_r_i[8];
  assign N1688 = N1431 & N1567;
  assign N1689 = N1431 & idx_r_i[8];
  assign N1690 = N1433 & N1567;
  assign N1691 = N1433 & idx_r_i[8];
  assign N1692 = N1435 & N1567;
  assign N1693 = N1435 & idx_r_i[8];
  assign N1694 = N1437 & N1567;
  assign N1695 = N1437 & idx_r_i[8];
  assign N1696 = N1439 & N1567;
  assign N1697 = N1439 & idx_r_i[8];
  assign N1698 = N1441 & N1567;
  assign N1699 = N1441 & idx_r_i[8];
  assign N1700 = N1443 & N1567;
  assign N1701 = N1443 & idx_r_i[8];
  assign N1702 = N1445 & N1567;
  assign N1703 = N1445 & idx_r_i[8];
  assign N1704 = N1447 & N1567;
  assign N1705 = N1447 & idx_r_i[8];
  assign N1706 = N1449 & N1567;
  assign N1707 = N1449 & idx_r_i[8];
  assign N1708 = N1451 & N1567;
  assign N1709 = N1451 & idx_r_i[8];
  assign N1710 = N1453 & N1567;
  assign N1711 = N1453 & idx_r_i[8];
  assign N1712 = N1455 & N1567;
  assign N1713 = N1455 & idx_r_i[8];
  assign N1714 = N1457 & N1567;
  assign N1715 = N1457 & idx_r_i[8];
  assign N1716 = N1459 & N1567;
  assign N1717 = N1459 & idx_r_i[8];
  assign N1718 = N1461 & N1567;
  assign N1719 = N1461 & idx_r_i[8];
  assign N1720 = N1463 & N1567;
  assign N1721 = N1463 & idx_r_i[8];
  assign N1722 = N1465 & N1567;
  assign N1723 = N1465 & idx_r_i[8];
  assign N1724 = N1467 & N1567;
  assign N1725 = N1467 & idx_r_i[8];
  assign N1726 = N1469 & N1567;
  assign N1727 = N1469 & idx_r_i[8];
  assign N1728 = N1471 & N1567;
  assign N1729 = N1471 & idx_r_i[8];
  assign N1730 = N1473 & N1567;
  assign N1731 = N1473 & idx_r_i[8];
  assign N1732 = N1475 & N1567;
  assign N1733 = N1475 & idx_r_i[8];
  assign N1734 = N1477 & N1567;
  assign N1735 = N1477 & idx_r_i[8];
  assign N1736 = N1479 & N1567;
  assign N1737 = N1479 & idx_r_i[8];
  assign N1738 = N1481 & N1567;
  assign N1739 = N1481 & idx_r_i[8];
  assign N1740 = N1483 & N1567;
  assign N1741 = N1483 & idx_r_i[8];
  assign N1742 = N1485 & N1567;
  assign N1743 = N1485 & idx_r_i[8];
  assign N1744 = N1487 & N1567;
  assign N1745 = N1487 & idx_r_i[8];
  assign N1746 = N1489 & N1567;
  assign N1747 = N1489 & idx_r_i[8];
  assign N1748 = N1491 & N1567;
  assign N1749 = N1491 & idx_r_i[8];
  assign N1750 = N1493 & N1567;
  assign N1751 = N1493 & idx_r_i[8];
  assign N1752 = N1495 & N1567;
  assign N1753 = N1495 & idx_r_i[8];
  assign N1754 = N1497 & N1567;
  assign N1755 = N1497 & idx_r_i[8];
  assign N1756 = N1499 & N1567;
  assign N1757 = N1499 & idx_r_i[8];
  assign N1758 = N1501 & N1567;
  assign N1759 = N1501 & idx_r_i[8];
  assign N1760 = N1503 & N1567;
  assign N1761 = N1503 & idx_r_i[8];
  assign N1762 = N1505 & N1567;
  assign N1763 = N1505 & idx_r_i[8];
  assign N1764 = N1507 & N1567;
  assign N1765 = N1507 & idx_r_i[8];
  assign N1766 = N1509 & N1567;
  assign N1767 = N1509 & idx_r_i[8];
  assign N1768 = N1511 & N1567;
  assign N1769 = N1511 & idx_r_i[8];
  assign N1770 = N1513 & N1567;
  assign N1771 = N1513 & idx_r_i[8];
  assign N1772 = N1515 & N1567;
  assign N1773 = N1515 & idx_r_i[8];
  assign N1774 = N1517 & N1567;
  assign N1775 = N1517 & idx_r_i[8];
  assign N1776 = N1519 & N1567;
  assign N1777 = N1519 & idx_r_i[8];
  assign N1778 = N1521 & N1567;
  assign N1779 = N1521 & idx_r_i[8];
  assign N1780 = N1523 & N1567;
  assign N1781 = N1523 & idx_r_i[8];
  assign N1782 = N1525 & N1567;
  assign N1783 = N1525 & idx_r_i[8];
  assign N1784 = N1527 & N1567;
  assign N1785 = N1527 & idx_r_i[8];
  assign N1786 = N1529 & N1567;
  assign N1787 = N1529 & idx_r_i[8];
  assign N1788 = N1531 & N1567;
  assign N1789 = N1531 & idx_r_i[8];
  assign N1790 = N1533 & N1567;
  assign N1791 = N1533 & idx_r_i[8];
  assign N1792 = N1535 & N1567;
  assign N1793 = N1535 & idx_r_i[8];
  assign N1794 = N1537 & N1567;
  assign N1795 = N1537 & idx_r_i[8];
  assign N1796 = N1539 & N1567;
  assign N1797 = N1539 & idx_r_i[8];
  assign N1798 = N1541 & N1567;
  assign N1799 = N1541 & idx_r_i[8];
  assign N1800 = N1543 & N1567;
  assign N1801 = N1543 & idx_r_i[8];
  assign N1802 = N1545 & N1567;
  assign N1803 = N1545 & idx_r_i[8];
  assign N1804 = N1547 & N1567;
  assign N1805 = N1547 & idx_r_i[8];
  assign N1806 = N1549 & N1567;
  assign N1807 = N1549 & idx_r_i[8];
  assign N1808 = N1551 & N1567;
  assign N1809 = N1551 & idx_r_i[8];
  assign N1810 = N1553 & N1567;
  assign N1811 = N1553 & idx_r_i[8];
  assign N1812 = N1555 & N1567;
  assign N1813 = N1555 & idx_r_i[8];
  assign N1814 = N1557 & N1567;
  assign N1815 = N1557 & idx_r_i[8];
  assign N1816 = N1559 & N1567;
  assign N1817 = N1559 & idx_r_i[8];
  assign N1818 = N1561 & N1567;
  assign N1819 = N1561 & idx_r_i[8];
  assign N1820 = N1563 & N1567;
  assign N1821 = N1563 & idx_r_i[8];
  assign N1822 = N1565 & N1567;
  assign N1823 = N1565 & idx_r_i[8];
  assign N1824 = N1312 & N1567;
  assign N1825 = N1312 & idx_r_i[8];
  assign N1826 = N1314 & N1567;
  assign N1827 = N1314 & idx_r_i[8];
  assign N1828 = N1316 & N1567;
  assign N1829 = N1316 & idx_r_i[8];
  assign N1830 = N1318 & N1567;
  assign N1831 = N1318 & idx_r_i[8];
  assign N1832 = N1320 & N1567;
  assign N1833 = N1320 & idx_r_i[8];
  assign N1834 = N1322 & N1567;
  assign N1835 = N1322 & idx_r_i[8];
  assign N1836 = N1324 & N1567;
  assign N1837 = N1324 & idx_r_i[8];
  assign N1838 = N1326 & N1567;
  assign N1839 = N1326 & idx_r_i[8];
  assign N1840 = N1328 & N1567;
  assign N1841 = N1328 & idx_r_i[8];
  assign N1842 = N1330 & N1567;
  assign N1843 = N1330 & idx_r_i[8];
  assign N1844 = N1332 & N1567;
  assign N1845 = N1332 & idx_r_i[8];
  assign N1846 = N1334 & N1567;
  assign N1847 = N1334 & idx_r_i[8];
  assign N1848 = N1336 & N1567;
  assign N1849 = N1336 & idx_r_i[8];
  assign N1850 = N1338 & N1567;
  assign N1851 = N1338 & idx_r_i[8];
  assign N1852 = N1340 & N1567;
  assign N1853 = N1340 & idx_r_i[8];
  assign N1854 = N1342 & N1567;
  assign N1855 = N1342 & idx_r_i[8];
  assign N1856 = N1344 & N1567;
  assign N1857 = N1344 & idx_r_i[8];
  assign N1858 = N1346 & N1567;
  assign N1859 = N1346 & idx_r_i[8];
  assign N1860 = N1348 & N1567;
  assign N1861 = N1348 & idx_r_i[8];
  assign N1862 = N1350 & N1567;
  assign N1863 = N1350 & idx_r_i[8];
  assign N1864 = N1352 & N1567;
  assign N1865 = N1352 & idx_r_i[8];
  assign N1866 = N1354 & N1567;
  assign N1867 = N1354 & idx_r_i[8];
  assign N1868 = N1356 & N1567;
  assign N1869 = N1356 & idx_r_i[8];
  assign N1870 = N1358 & N1567;
  assign N1871 = N1358 & idx_r_i[8];
  assign N1872 = N1360 & N1567;
  assign N1873 = N1360 & idx_r_i[8];
  assign N1874 = N1362 & N1567;
  assign N1875 = N1362 & idx_r_i[8];
  assign N1876 = N1364 & N1567;
  assign N1877 = N1364 & idx_r_i[8];
  assign N1878 = N1366 & N1567;
  assign N1879 = N1366 & idx_r_i[8];
  assign N1880 = N1368 & N1567;
  assign N1881 = N1368 & idx_r_i[8];
  assign N1882 = N1370 & N1567;
  assign N1883 = N1370 & idx_r_i[8];
  assign N1884 = N1372 & N1567;
  assign N1885 = N1372 & idx_r_i[8];
  assign N1886 = N1374 & N1567;
  assign N1887 = N1374 & idx_r_i[8];
  assign N1888 = N1376 & N1567;
  assign N1889 = N1376 & idx_r_i[8];
  assign N1890 = N1378 & N1567;
  assign N1891 = N1378 & idx_r_i[8];
  assign N1892 = N1380 & N1567;
  assign N1893 = N1380 & idx_r_i[8];
  assign N1894 = N1382 & N1567;
  assign N1895 = N1382 & idx_r_i[8];
  assign N1896 = N1384 & N1567;
  assign N1897 = N1384 & idx_r_i[8];
  assign N1898 = N1386 & N1567;
  assign N1899 = N1386 & idx_r_i[8];
  assign N1900 = N1388 & N1567;
  assign N1901 = N1388 & idx_r_i[8];
  assign N1902 = N1390 & N1567;
  assign N1903 = N1390 & idx_r_i[8];
  assign N1904 = N1392 & N1567;
  assign N1905 = N1392 & idx_r_i[8];
  assign N1906 = N1394 & N1567;
  assign N1907 = N1394 & idx_r_i[8];
  assign N1908 = N1396 & N1567;
  assign N1909 = N1396 & idx_r_i[8];
  assign N1910 = N1398 & N1567;
  assign N1911 = N1398 & idx_r_i[8];
  assign N1912 = N1400 & N1567;
  assign N1913 = N1400 & idx_r_i[8];
  assign N1914 = N1402 & N1567;
  assign N1915 = N1402 & idx_r_i[8];
  assign N1916 = N1404 & N1567;
  assign N1917 = N1404 & idx_r_i[8];
  assign N1918 = N1406 & N1567;
  assign N1919 = N1406 & idx_r_i[8];
  assign N1920 = N1408 & N1567;
  assign N1921 = N1408 & idx_r_i[8];
  assign N1922 = N1410 & N1567;
  assign N1923 = N1410 & idx_r_i[8];
  assign N1924 = N1412 & N1567;
  assign N1925 = N1412 & idx_r_i[8];
  assign N1926 = N1414 & N1567;
  assign N1927 = N1414 & idx_r_i[8];
  assign N1928 = N1416 & N1567;
  assign N1929 = N1416 & idx_r_i[8];
  assign N1930 = N1418 & N1567;
  assign N1931 = N1418 & idx_r_i[8];
  assign N1932 = N1420 & N1567;
  assign N1933 = N1420 & idx_r_i[8];
  assign N1934 = N1422 & N1567;
  assign N1935 = N1422 & idx_r_i[8];
  assign N1936 = N1424 & N1567;
  assign N1937 = N1424 & idx_r_i[8];
  assign N1938 = N1426 & N1567;
  assign N1939 = N1426 & idx_r_i[8];
  assign N1940 = N1428 & N1567;
  assign N1941 = N1428 & idx_r_i[8];
  assign N1942 = N1430 & N1567;
  assign N1943 = N1430 & idx_r_i[8];
  assign N1944 = N1432 & N1567;
  assign N1945 = N1432 & idx_r_i[8];
  assign N1946 = N1434 & N1567;
  assign N1947 = N1434 & idx_r_i[8];
  assign N1948 = N1436 & N1567;
  assign N1949 = N1436 & idx_r_i[8];
  assign N1950 = N1438 & N1567;
  assign N1951 = N1438 & idx_r_i[8];
  assign N1952 = N1440 & N1567;
  assign N1953 = N1440 & idx_r_i[8];
  assign N1954 = N1442 & N1567;
  assign N1955 = N1442 & idx_r_i[8];
  assign N1956 = N1444 & N1567;
  assign N1957 = N1444 & idx_r_i[8];
  assign N1958 = N1446 & N1567;
  assign N1959 = N1446 & idx_r_i[8];
  assign N1960 = N1448 & N1567;
  assign N1961 = N1448 & idx_r_i[8];
  assign N1962 = N1450 & N1567;
  assign N1963 = N1450 & idx_r_i[8];
  assign N1964 = N1452 & N1567;
  assign N1965 = N1452 & idx_r_i[8];
  assign N1966 = N1454 & N1567;
  assign N1967 = N1454 & idx_r_i[8];
  assign N1968 = N1456 & N1567;
  assign N1969 = N1456 & idx_r_i[8];
  assign N1970 = N1458 & N1567;
  assign N1971 = N1458 & idx_r_i[8];
  assign N1972 = N1460 & N1567;
  assign N1973 = N1460 & idx_r_i[8];
  assign N1974 = N1462 & N1567;
  assign N1975 = N1462 & idx_r_i[8];
  assign N1976 = N1464 & N1567;
  assign N1977 = N1464 & idx_r_i[8];
  assign N1978 = N1466 & N1567;
  assign N1979 = N1466 & idx_r_i[8];
  assign N1980 = N1468 & N1567;
  assign N1981 = N1468 & idx_r_i[8];
  assign N1982 = N1470 & N1567;
  assign N1983 = N1470 & idx_r_i[8];
  assign N1984 = N1472 & N1567;
  assign N1985 = N1472 & idx_r_i[8];
  assign N1986 = N1474 & N1567;
  assign N1987 = N1474 & idx_r_i[8];
  assign N1988 = N1476 & N1567;
  assign N1989 = N1476 & idx_r_i[8];
  assign N1990 = N1478 & N1567;
  assign N1991 = N1478 & idx_r_i[8];
  assign N1992 = N1480 & N1567;
  assign N1993 = N1480 & idx_r_i[8];
  assign N1994 = N1482 & N1567;
  assign N1995 = N1482 & idx_r_i[8];
  assign N1996 = N1484 & N1567;
  assign N1997 = N1484 & idx_r_i[8];
  assign N1998 = N1486 & N1567;
  assign N1999 = N1486 & idx_r_i[8];
  assign N2000 = N1488 & N1567;
  assign N2001 = N1488 & idx_r_i[8];
  assign N2002 = N1490 & N1567;
  assign N2003 = N1490 & idx_r_i[8];
  assign N2004 = N1492 & N1567;
  assign N2005 = N1492 & idx_r_i[8];
  assign N2006 = N1494 & N1567;
  assign N2007 = N1494 & idx_r_i[8];
  assign N2008 = N1496 & N1567;
  assign N2009 = N1496 & idx_r_i[8];
  assign N2010 = N1498 & N1567;
  assign N2011 = N1498 & idx_r_i[8];
  assign N2012 = N1500 & N1567;
  assign N2013 = N1500 & idx_r_i[8];
  assign N2014 = N1502 & N1567;
  assign N2015 = N1502 & idx_r_i[8];
  assign N2016 = N1504 & N1567;
  assign N2017 = N1504 & idx_r_i[8];
  assign N2018 = N1506 & N1567;
  assign N2019 = N1506 & idx_r_i[8];
  assign N2020 = N1508 & N1567;
  assign N2021 = N1508 & idx_r_i[8];
  assign N2022 = N1510 & N1567;
  assign N2023 = N1510 & idx_r_i[8];
  assign N2024 = N1512 & N1567;
  assign N2025 = N1512 & idx_r_i[8];
  assign N2026 = N1514 & N1567;
  assign N2027 = N1514 & idx_r_i[8];
  assign N2028 = N1516 & N1567;
  assign N2029 = N1516 & idx_r_i[8];
  assign N2030 = N1518 & N1567;
  assign N2031 = N1518 & idx_r_i[8];
  assign N2032 = N1520 & N1567;
  assign N2033 = N1520 & idx_r_i[8];
  assign N2034 = N1522 & N1567;
  assign N2035 = N1522 & idx_r_i[8];
  assign N2036 = N1524 & N1567;
  assign N2037 = N1524 & idx_r_i[8];
  assign N2038 = N1526 & N1567;
  assign N2039 = N1526 & idx_r_i[8];
  assign N2040 = N1528 & N1567;
  assign N2041 = N1528 & idx_r_i[8];
  assign N2042 = N1530 & N1567;
  assign N2043 = N1530 & idx_r_i[8];
  assign N2044 = N1532 & N1567;
  assign N2045 = N1532 & idx_r_i[8];
  assign N2046 = N1534 & N1567;
  assign N2047 = N1534 & idx_r_i[8];
  assign N2048 = N1536 & N1567;
  assign N2049 = N1536 & idx_r_i[8];
  assign N2050 = N1538 & N1567;
  assign N2051 = N1538 & idx_r_i[8];
  assign N2052 = N1540 & N1567;
  assign N2053 = N1540 & idx_r_i[8];
  assign N2054 = N1542 & N1567;
  assign N2055 = N1542 & idx_r_i[8];
  assign N2056 = N1544 & N1567;
  assign N2057 = N1544 & idx_r_i[8];
  assign N2058 = N1546 & N1567;
  assign N2059 = N1546 & idx_r_i[8];
  assign N2060 = N1548 & N1567;
  assign N2061 = N1548 & idx_r_i[8];
  assign N2062 = N1550 & N1567;
  assign N2063 = N1550 & idx_r_i[8];
  assign N2064 = N1552 & N1567;
  assign N2065 = N1552 & idx_r_i[8];
  assign N2066 = N1554 & N1567;
  assign N2067 = N1554 & idx_r_i[8];
  assign N2068 = N1556 & N1567;
  assign N2069 = N1556 & idx_r_i[8];
  assign N2070 = N1558 & N1567;
  assign N2071 = N1558 & idx_r_i[8];
  assign N2072 = N1560 & N1567;
  assign N2073 = N1560 & idx_r_i[8];
  assign N2074 = N1562 & N1567;
  assign N2075 = N1562 & idx_r_i[8];
  assign N2076 = N1564 & N1567;
  assign N2077 = N1564 & idx_r_i[8];
  assign N2078 = N1566 & N1567;
  assign N2079 = N1566 & idx_r_i[8];
  assign n_0_net_ = w_v_i | r_v_i;

  always @(posedge clk_i) begin
    if(N1047) begin
      { valid[511:511] } <= { N541 };
    end
    if(N1046) begin
      { valid[510:510] } <= { N541 };
    end
    if(N1045) begin
      { valid[509:509] } <= { N541 };
    end
    if(N1044) begin
      { valid[508:508] } <= { N541 };
    end
    if(N1043) begin
      { valid[507:507] } <= { N541 };
    end
    if(N1042) begin
      { valid[506:506] } <= { N541 };
    end
    if(N1041) begin
      { valid[505:505] } <= { N541 };
    end
    if(N1040) begin
      { valid[504:504] } <= { N541 };
    end
    if(N1039) begin
      { valid[503:503] } <= { N541 };
    end
    if(N1038) begin
      { valid[502:502] } <= { N541 };
    end
    if(N1037) begin
      { valid[501:501] } <= { N541 };
    end
    if(N1036) begin
      { valid[500:500] } <= { N541 };
    end
    if(N1035) begin
      { valid[499:499] } <= { N541 };
    end
    if(N1034) begin
      { valid[498:498] } <= { N541 };
    end
    if(N1033) begin
      { valid[497:497] } <= { N541 };
    end
    if(N1032) begin
      { valid[496:496] } <= { N541 };
    end
    if(N1031) begin
      { valid[495:495] } <= { N541 };
    end
    if(N1030) begin
      { valid[494:494] } <= { N541 };
    end
    if(N1029) begin
      { valid[493:493] } <= { N541 };
    end
    if(N1028) begin
      { valid[492:492] } <= { N541 };
    end
    if(N1027) begin
      { valid[491:491] } <= { N541 };
    end
    if(N1026) begin
      { valid[490:490] } <= { N541 };
    end
    if(N1025) begin
      { valid[489:489] } <= { N541 };
    end
    if(N1024) begin
      { valid[488:488] } <= { N541 };
    end
    if(N1023) begin
      { valid[487:487] } <= { N541 };
    end
    if(N1022) begin
      { valid[486:486] } <= { N541 };
    end
    if(N1021) begin
      { valid[485:485] } <= { N541 };
    end
    if(N1020) begin
      { valid[484:484] } <= { N541 };
    end
    if(N1019) begin
      { valid[483:483] } <= { N541 };
    end
    if(N1018) begin
      { valid[482:482] } <= { N541 };
    end
    if(N1017) begin
      { valid[481:481] } <= { N541 };
    end
    if(N1016) begin
      { valid[480:480] } <= { N541 };
    end
    if(N1015) begin
      { valid[479:479] } <= { N541 };
    end
    if(N1014) begin
      { valid[478:478] } <= { N541 };
    end
    if(N1013) begin
      { valid[477:477] } <= { N541 };
    end
    if(N1012) begin
      { valid[476:476] } <= { N541 };
    end
    if(N1011) begin
      { valid[475:475] } <= { N541 };
    end
    if(N1010) begin
      { valid[474:474] } <= { N541 };
    end
    if(N1009) begin
      { valid[473:473] } <= { N541 };
    end
    if(N1008) begin
      { valid[472:472] } <= { N541 };
    end
    if(N1007) begin
      { valid[471:471] } <= { N541 };
    end
    if(N1006) begin
      { valid[470:470] } <= { N541 };
    end
    if(N1005) begin
      { valid[469:469] } <= { N541 };
    end
    if(N1004) begin
      { valid[468:468] } <= { N541 };
    end
    if(N1003) begin
      { valid[467:467] } <= { N541 };
    end
    if(N1002) begin
      { valid[466:466] } <= { N541 };
    end
    if(N1001) begin
      { valid[465:465] } <= { N541 };
    end
    if(N1000) begin
      { valid[464:464] } <= { N541 };
    end
    if(N999) begin
      { valid[463:463] } <= { N541 };
    end
    if(N998) begin
      { valid[462:462] } <= { N541 };
    end
    if(N997) begin
      { valid[461:461] } <= { N541 };
    end
    if(N996) begin
      { valid[460:460] } <= { N541 };
    end
    if(N995) begin
      { valid[459:459] } <= { N541 };
    end
    if(N994) begin
      { valid[458:458] } <= { N541 };
    end
    if(N993) begin
      { valid[457:457] } <= { N541 };
    end
    if(N992) begin
      { valid[456:456] } <= { N541 };
    end
    if(N991) begin
      { valid[455:455] } <= { N541 };
    end
    if(N990) begin
      { valid[454:454] } <= { N541 };
    end
    if(N989) begin
      { valid[453:453] } <= { N541 };
    end
    if(N988) begin
      { valid[452:452] } <= { N541 };
    end
    if(N987) begin
      { valid[451:451] } <= { N541 };
    end
    if(N986) begin
      { valid[450:450] } <= { N541 };
    end
    if(N985) begin
      { valid[449:449] } <= { N541 };
    end
    if(N984) begin
      { valid[448:448] } <= { N541 };
    end
    if(N983) begin
      { valid[447:447] } <= { N541 };
    end
    if(N982) begin
      { valid[446:446] } <= { N541 };
    end
    if(N981) begin
      { valid[445:445] } <= { N541 };
    end
    if(N980) begin
      { valid[444:444] } <= { N541 };
    end
    if(N979) begin
      { valid[443:443] } <= { N541 };
    end
    if(N978) begin
      { valid[442:442] } <= { N541 };
    end
    if(N977) begin
      { valid[441:441] } <= { N541 };
    end
    if(N976) begin
      { valid[440:440] } <= { N541 };
    end
    if(N975) begin
      { valid[439:439] } <= { N541 };
    end
    if(N974) begin
      { valid[438:438] } <= { N541 };
    end
    if(N973) begin
      { valid[437:437] } <= { N541 };
    end
    if(N972) begin
      { valid[436:436] } <= { N541 };
    end
    if(N971) begin
      { valid[435:435] } <= { N541 };
    end
    if(N970) begin
      { valid[434:434] } <= { N541 };
    end
    if(N969) begin
      { valid[433:433] } <= { N541 };
    end
    if(N968) begin
      { valid[432:432] } <= { N541 };
    end
    if(N967) begin
      { valid[431:431] } <= { N541 };
    end
    if(N966) begin
      { valid[430:430] } <= { N541 };
    end
    if(N965) begin
      { valid[429:429] } <= { N541 };
    end
    if(N964) begin
      { valid[428:428] } <= { N541 };
    end
    if(N963) begin
      { valid[427:427] } <= { N541 };
    end
    if(N962) begin
      { valid[426:426] } <= { N541 };
    end
    if(N961) begin
      { valid[425:425] } <= { N541 };
    end
    if(N960) begin
      { valid[424:424] } <= { N541 };
    end
    if(N959) begin
      { valid[423:423] } <= { N541 };
    end
    if(N958) begin
      { valid[422:422] } <= { N541 };
    end
    if(N957) begin
      { valid[421:421] } <= { N541 };
    end
    if(N956) begin
      { valid[420:420] } <= { N541 };
    end
    if(N955) begin
      { valid[419:419] } <= { N541 };
    end
    if(N954) begin
      { valid[418:418] } <= { N541 };
    end
    if(N953) begin
      { valid[417:417] } <= { N541 };
    end
    if(N952) begin
      { valid[416:416] } <= { N541 };
    end
    if(N951) begin
      { valid[415:415] } <= { N541 };
    end
    if(N950) begin
      { valid[414:414] } <= { N541 };
    end
    if(N949) begin
      { valid[413:413] } <= { N541 };
    end
    if(N948) begin
      { valid[412:412] } <= { N541 };
    end
    if(N947) begin
      { valid[411:411] } <= { N541 };
    end
    if(N946) begin
      { valid[410:410] } <= { N541 };
    end
    if(N945) begin
      { valid[409:409] } <= { N541 };
    end
    if(N944) begin
      { valid[408:408] } <= { N541 };
    end
    if(N943) begin
      { valid[407:407] } <= { N541 };
    end
    if(N942) begin
      { valid[406:406] } <= { N541 };
    end
    if(N941) begin
      { valid[405:405] } <= { N541 };
    end
    if(N940) begin
      { valid[404:404] } <= { N541 };
    end
    if(N939) begin
      { valid[403:403] } <= { N541 };
    end
    if(N938) begin
      { valid[402:402] } <= { N541 };
    end
    if(N937) begin
      { valid[401:401] } <= { N541 };
    end
    if(N936) begin
      { valid[400:400] } <= { N541 };
    end
    if(N935) begin
      { valid[399:399] } <= { N541 };
    end
    if(N934) begin
      { valid[398:398] } <= { N541 };
    end
    if(N933) begin
      { valid[397:397] } <= { N541 };
    end
    if(N932) begin
      { valid[396:396] } <= { N541 };
    end
    if(N931) begin
      { valid[395:395] } <= { N541 };
    end
    if(N930) begin
      { valid[394:394] } <= { N541 };
    end
    if(N929) begin
      { valid[393:393] } <= { N541 };
    end
    if(N928) begin
      { valid[392:392] } <= { N541 };
    end
    if(N927) begin
      { valid[391:391] } <= { N541 };
    end
    if(N926) begin
      { valid[390:390] } <= { N541 };
    end
    if(N925) begin
      { valid[389:389] } <= { N541 };
    end
    if(N924) begin
      { valid[388:388] } <= { N541 };
    end
    if(N923) begin
      { valid[387:387] } <= { N541 };
    end
    if(N922) begin
      { valid[386:386] } <= { N541 };
    end
    if(N921) begin
      { valid[385:385] } <= { N541 };
    end
    if(N920) begin
      { valid[384:384] } <= { N541 };
    end
    if(N919) begin
      { valid[383:383] } <= { N541 };
    end
    if(N918) begin
      { valid[382:382] } <= { N541 };
    end
    if(N917) begin
      { valid[381:381] } <= { N541 };
    end
    if(N916) begin
      { valid[380:380] } <= { N541 };
    end
    if(N915) begin
      { valid[379:379] } <= { N541 };
    end
    if(N914) begin
      { valid[378:378] } <= { N541 };
    end
    if(N913) begin
      { valid[377:377] } <= { N541 };
    end
    if(N912) begin
      { valid[376:376] } <= { N541 };
    end
    if(N911) begin
      { valid[375:375] } <= { N541 };
    end
    if(N910) begin
      { valid[374:374] } <= { N541 };
    end
    if(N909) begin
      { valid[373:373] } <= { N541 };
    end
    if(N908) begin
      { valid[372:372] } <= { N541 };
    end
    if(N907) begin
      { valid[371:371] } <= { N541 };
    end
    if(N906) begin
      { valid[370:370] } <= { N541 };
    end
    if(N905) begin
      { valid[369:369] } <= { N541 };
    end
    if(N904) begin
      { valid[368:368] } <= { N541 };
    end
    if(N903) begin
      { valid[367:367] } <= { N541 };
    end
    if(N902) begin
      { valid[366:366] } <= { N541 };
    end
    if(N901) begin
      { valid[365:365] } <= { N541 };
    end
    if(N900) begin
      { valid[364:364] } <= { N541 };
    end
    if(N899) begin
      { valid[363:363] } <= { N541 };
    end
    if(N898) begin
      { valid[362:362] } <= { N541 };
    end
    if(N897) begin
      { valid[361:361] } <= { N541 };
    end
    if(N896) begin
      { valid[360:360] } <= { N541 };
    end
    if(N895) begin
      { valid[359:359] } <= { N541 };
    end
    if(N894) begin
      { valid[358:358] } <= { N541 };
    end
    if(N893) begin
      { valid[357:357] } <= { N541 };
    end
    if(N892) begin
      { valid[356:356] } <= { N541 };
    end
    if(N891) begin
      { valid[355:355] } <= { N541 };
    end
    if(N890) begin
      { valid[354:354] } <= { N541 };
    end
    if(N889) begin
      { valid[353:353] } <= { N541 };
    end
    if(N888) begin
      { valid[352:352] } <= { N541 };
    end
    if(N887) begin
      { valid[351:351] } <= { N541 };
    end
    if(N886) begin
      { valid[350:350] } <= { N541 };
    end
    if(N885) begin
      { valid[349:349] } <= { N541 };
    end
    if(N884) begin
      { valid[348:348] } <= { N541 };
    end
    if(N883) begin
      { valid[347:347] } <= { N541 };
    end
    if(N882) begin
      { valid[346:346] } <= { N541 };
    end
    if(N881) begin
      { valid[345:345] } <= { N541 };
    end
    if(N880) begin
      { valid[344:344] } <= { N541 };
    end
    if(N879) begin
      { valid[343:343] } <= { N541 };
    end
    if(N878) begin
      { valid[342:342] } <= { N541 };
    end
    if(N877) begin
      { valid[341:341] } <= { N541 };
    end
    if(N876) begin
      { valid[340:340] } <= { N541 };
    end
    if(N875) begin
      { valid[339:339] } <= { N541 };
    end
    if(N874) begin
      { valid[338:338] } <= { N541 };
    end
    if(N873) begin
      { valid[337:337] } <= { N541 };
    end
    if(N872) begin
      { valid[336:336] } <= { N541 };
    end
    if(N871) begin
      { valid[335:335] } <= { N541 };
    end
    if(N870) begin
      { valid[334:334] } <= { N541 };
    end
    if(N869) begin
      { valid[333:333] } <= { N541 };
    end
    if(N868) begin
      { valid[332:332] } <= { N541 };
    end
    if(N867) begin
      { valid[331:331] } <= { N541 };
    end
    if(N866) begin
      { valid[330:330] } <= { N541 };
    end
    if(N865) begin
      { valid[329:329] } <= { N541 };
    end
    if(N864) begin
      { valid[328:328] } <= { N541 };
    end
    if(N863) begin
      { valid[327:327] } <= { N541 };
    end
    if(N862) begin
      { valid[326:326] } <= { N541 };
    end
    if(N861) begin
      { valid[325:325] } <= { N541 };
    end
    if(N860) begin
      { valid[324:324] } <= { N541 };
    end
    if(N859) begin
      { valid[323:323] } <= { N541 };
    end
    if(N858) begin
      { valid[322:322] } <= { N541 };
    end
    if(N857) begin
      { valid[321:321] } <= { N541 };
    end
    if(N856) begin
      { valid[320:320] } <= { N541 };
    end
    if(N855) begin
      { valid[319:319] } <= { N541 };
    end
    if(N854) begin
      { valid[318:318] } <= { N541 };
    end
    if(N853) begin
      { valid[317:317] } <= { N541 };
    end
    if(N852) begin
      { valid[316:316] } <= { N541 };
    end
    if(N851) begin
      { valid[315:315] } <= { N541 };
    end
    if(N850) begin
      { valid[314:314] } <= { N541 };
    end
    if(N849) begin
      { valid[313:313] } <= { N541 };
    end
    if(N848) begin
      { valid[312:312] } <= { N541 };
    end
    if(N847) begin
      { valid[311:311] } <= { N541 };
    end
    if(N846) begin
      { valid[310:310] } <= { N541 };
    end
    if(N845) begin
      { valid[309:309] } <= { N541 };
    end
    if(N844) begin
      { valid[308:308] } <= { N541 };
    end
    if(N843) begin
      { valid[307:307] } <= { N541 };
    end
    if(N842) begin
      { valid[306:306] } <= { N541 };
    end
    if(N841) begin
      { valid[305:305] } <= { N541 };
    end
    if(N840) begin
      { valid[304:304] } <= { N541 };
    end
    if(N839) begin
      { valid[303:303] } <= { N541 };
    end
    if(N838) begin
      { valid[302:302] } <= { N541 };
    end
    if(N837) begin
      { valid[301:301] } <= { N541 };
    end
    if(N836) begin
      { valid[300:300] } <= { N541 };
    end
    if(N835) begin
      { valid[299:299] } <= { N541 };
    end
    if(N834) begin
      { valid[298:298] } <= { N541 };
    end
    if(N833) begin
      { valid[297:297] } <= { N541 };
    end
    if(N832) begin
      { valid[296:296] } <= { N541 };
    end
    if(N831) begin
      { valid[295:295] } <= { N541 };
    end
    if(N830) begin
      { valid[294:294] } <= { N541 };
    end
    if(N829) begin
      { valid[293:293] } <= { N541 };
    end
    if(N828) begin
      { valid[292:292] } <= { N541 };
    end
    if(N827) begin
      { valid[291:291] } <= { N541 };
    end
    if(N826) begin
      { valid[290:290] } <= { N541 };
    end
    if(N825) begin
      { valid[289:289] } <= { N541 };
    end
    if(N824) begin
      { valid[288:288] } <= { N541 };
    end
    if(N823) begin
      { valid[287:287] } <= { N541 };
    end
    if(N822) begin
      { valid[286:286] } <= { N541 };
    end
    if(N821) begin
      { valid[285:285] } <= { N541 };
    end
    if(N820) begin
      { valid[284:284] } <= { N541 };
    end
    if(N819) begin
      { valid[283:283] } <= { N541 };
    end
    if(N818) begin
      { valid[282:282] } <= { N541 };
    end
    if(N817) begin
      { valid[281:281] } <= { N541 };
    end
    if(N816) begin
      { valid[280:280] } <= { N541 };
    end
    if(N815) begin
      { valid[279:279] } <= { N541 };
    end
    if(N814) begin
      { valid[278:278] } <= { N541 };
    end
    if(N813) begin
      { valid[277:277] } <= { N541 };
    end
    if(N812) begin
      { valid[276:276] } <= { N541 };
    end
    if(N811) begin
      { valid[275:275] } <= { N541 };
    end
    if(N810) begin
      { valid[274:274] } <= { N541 };
    end
    if(N809) begin
      { valid[273:273] } <= { N541 };
    end
    if(N808) begin
      { valid[272:272] } <= { N541 };
    end
    if(N807) begin
      { valid[271:271] } <= { N541 };
    end
    if(N806) begin
      { valid[270:270] } <= { N541 };
    end
    if(N805) begin
      { valid[269:269] } <= { N541 };
    end
    if(N804) begin
      { valid[268:268] } <= { N541 };
    end
    if(N803) begin
      { valid[267:267] } <= { N541 };
    end
    if(N802) begin
      { valid[266:266] } <= { N541 };
    end
    if(N801) begin
      { valid[265:265] } <= { N541 };
    end
    if(N800) begin
      { valid[264:264] } <= { N541 };
    end
    if(N799) begin
      { valid[263:263] } <= { N541 };
    end
    if(N798) begin
      { valid[262:262] } <= { N541 };
    end
    if(N797) begin
      { valid[261:261] } <= { N541 };
    end
    if(N796) begin
      { valid[260:260] } <= { N541 };
    end
    if(N795) begin
      { valid[259:259] } <= { N541 };
    end
    if(N794) begin
      { valid[258:258] } <= { N541 };
    end
    if(N793) begin
      { valid[257:257] } <= { N541 };
    end
    if(N792) begin
      { valid[256:256] } <= { N541 };
    end
    if(N791) begin
      { valid[255:255] } <= { N541 };
    end
    if(N790) begin
      { valid[254:254] } <= { N541 };
    end
    if(N789) begin
      { valid[253:253] } <= { N541 };
    end
    if(N788) begin
      { valid[252:252] } <= { N541 };
    end
    if(N787) begin
      { valid[251:251] } <= { N541 };
    end
    if(N786) begin
      { valid[250:250] } <= { N541 };
    end
    if(N785) begin
      { valid[249:249] } <= { N541 };
    end
    if(N784) begin
      { valid[248:248] } <= { N541 };
    end
    if(N783) begin
      { valid[247:247] } <= { N541 };
    end
    if(N782) begin
      { valid[246:246] } <= { N541 };
    end
    if(N781) begin
      { valid[245:245] } <= { N541 };
    end
    if(N780) begin
      { valid[244:244] } <= { N541 };
    end
    if(N779) begin
      { valid[243:243] } <= { N541 };
    end
    if(N778) begin
      { valid[242:242] } <= { N541 };
    end
    if(N777) begin
      { valid[241:241] } <= { N541 };
    end
    if(N776) begin
      { valid[240:240] } <= { N541 };
    end
    if(N775) begin
      { valid[239:239] } <= { N541 };
    end
    if(N774) begin
      { valid[238:238] } <= { N541 };
    end
    if(N773) begin
      { valid[237:237] } <= { N541 };
    end
    if(N772) begin
      { valid[236:236] } <= { N541 };
    end
    if(N771) begin
      { valid[235:235] } <= { N541 };
    end
    if(N770) begin
      { valid[234:234] } <= { N541 };
    end
    if(N769) begin
      { valid[233:233] } <= { N541 };
    end
    if(N768) begin
      { valid[232:232] } <= { N541 };
    end
    if(N767) begin
      { valid[231:231] } <= { N541 };
    end
    if(N766) begin
      { valid[230:230] } <= { N541 };
    end
    if(N765) begin
      { valid[229:229] } <= { N541 };
    end
    if(N764) begin
      { valid[228:228] } <= { N541 };
    end
    if(N763) begin
      { valid[227:227] } <= { N541 };
    end
    if(N762) begin
      { valid[226:226] } <= { N541 };
    end
    if(N761) begin
      { valid[225:225] } <= { N541 };
    end
    if(N760) begin
      { valid[224:224] } <= { N541 };
    end
    if(N759) begin
      { valid[223:223] } <= { N541 };
    end
    if(N758) begin
      { valid[222:222] } <= { N541 };
    end
    if(N757) begin
      { valid[221:221] } <= { N541 };
    end
    if(N756) begin
      { valid[220:220] } <= { N541 };
    end
    if(N755) begin
      { valid[219:219] } <= { N541 };
    end
    if(N754) begin
      { valid[218:218] } <= { N541 };
    end
    if(N753) begin
      { valid[217:217] } <= { N541 };
    end
    if(N752) begin
      { valid[216:216] } <= { N541 };
    end
    if(N751) begin
      { valid[215:215] } <= { N541 };
    end
    if(N750) begin
      { valid[214:214] } <= { N541 };
    end
    if(N749) begin
      { valid[213:213] } <= { N541 };
    end
    if(N748) begin
      { valid[212:212] } <= { N541 };
    end
    if(N747) begin
      { valid[211:211] } <= { N541 };
    end
    if(N746) begin
      { valid[210:210] } <= { N541 };
    end
    if(N745) begin
      { valid[209:209] } <= { N541 };
    end
    if(N744) begin
      { valid[208:208] } <= { N541 };
    end
    if(N743) begin
      { valid[207:207] } <= { N541 };
    end
    if(N742) begin
      { valid[206:206] } <= { N541 };
    end
    if(N741) begin
      { valid[205:205] } <= { N541 };
    end
    if(N740) begin
      { valid[204:204] } <= { N541 };
    end
    if(N739) begin
      { valid[203:203] } <= { N541 };
    end
    if(N738) begin
      { valid[202:202] } <= { N541 };
    end
    if(N737) begin
      { valid[201:201] } <= { N541 };
    end
    if(N736) begin
      { valid[200:200] } <= { N541 };
    end
    if(N735) begin
      { valid[199:199] } <= { N541 };
    end
    if(N734) begin
      { valid[198:198] } <= { N541 };
    end
    if(N733) begin
      { valid[197:197] } <= { N541 };
    end
    if(N732) begin
      { valid[196:196] } <= { N541 };
    end
    if(N731) begin
      { valid[195:195] } <= { N541 };
    end
    if(N730) begin
      { valid[194:194] } <= { N541 };
    end
    if(N729) begin
      { valid[193:193] } <= { N541 };
    end
    if(N728) begin
      { valid[192:192] } <= { N541 };
    end
    if(N727) begin
      { valid[191:191] } <= { N541 };
    end
    if(N726) begin
      { valid[190:190] } <= { N541 };
    end
    if(N725) begin
      { valid[189:189] } <= { N541 };
    end
    if(N724) begin
      { valid[188:188] } <= { N541 };
    end
    if(N723) begin
      { valid[187:187] } <= { N541 };
    end
    if(N722) begin
      { valid[186:186] } <= { N541 };
    end
    if(N721) begin
      { valid[185:185] } <= { N541 };
    end
    if(N720) begin
      { valid[184:184] } <= { N541 };
    end
    if(N719) begin
      { valid[183:183] } <= { N541 };
    end
    if(N718) begin
      { valid[182:182] } <= { N541 };
    end
    if(N717) begin
      { valid[181:181] } <= { N541 };
    end
    if(N716) begin
      { valid[180:180] } <= { N541 };
    end
    if(N715) begin
      { valid[179:179] } <= { N541 };
    end
    if(N714) begin
      { valid[178:178] } <= { N541 };
    end
    if(N713) begin
      { valid[177:177] } <= { N541 };
    end
    if(N712) begin
      { valid[176:176] } <= { N541 };
    end
    if(N711) begin
      { valid[175:175] } <= { N541 };
    end
    if(N710) begin
      { valid[174:174] } <= { N541 };
    end
    if(N709) begin
      { valid[173:173] } <= { N541 };
    end
    if(N708) begin
      { valid[172:172] } <= { N541 };
    end
    if(N707) begin
      { valid[171:171] } <= { N541 };
    end
    if(N706) begin
      { valid[170:170] } <= { N541 };
    end
    if(N705) begin
      { valid[169:169] } <= { N541 };
    end
    if(N704) begin
      { valid[168:168] } <= { N541 };
    end
    if(N703) begin
      { valid[167:167] } <= { N541 };
    end
    if(N702) begin
      { valid[166:166] } <= { N541 };
    end
    if(N701) begin
      { valid[165:165] } <= { N541 };
    end
    if(N700) begin
      { valid[164:164] } <= { N541 };
    end
    if(N699) begin
      { valid[163:163] } <= { N541 };
    end
    if(N698) begin
      { valid[162:162] } <= { N541 };
    end
    if(N697) begin
      { valid[161:161] } <= { N541 };
    end
    if(N696) begin
      { valid[160:160] } <= { N541 };
    end
    if(N695) begin
      { valid[159:159] } <= { N541 };
    end
    if(N694) begin
      { valid[158:158] } <= { N541 };
    end
    if(N693) begin
      { valid[157:157] } <= { N541 };
    end
    if(N692) begin
      { valid[156:156] } <= { N541 };
    end
    if(N691) begin
      { valid[155:155] } <= { N541 };
    end
    if(N690) begin
      { valid[154:154] } <= { N541 };
    end
    if(N689) begin
      { valid[153:153] } <= { N541 };
    end
    if(N688) begin
      { valid[152:152] } <= { N541 };
    end
    if(N687) begin
      { valid[151:151] } <= { N541 };
    end
    if(N686) begin
      { valid[150:150] } <= { N541 };
    end
    if(N685) begin
      { valid[149:149] } <= { N541 };
    end
    if(N684) begin
      { valid[148:148] } <= { N541 };
    end
    if(N683) begin
      { valid[147:147] } <= { N541 };
    end
    if(N682) begin
      { valid[146:146] } <= { N541 };
    end
    if(N681) begin
      { valid[145:145] } <= { N541 };
    end
    if(N680) begin
      { valid[144:144] } <= { N541 };
    end
    if(N679) begin
      { valid[143:143] } <= { N541 };
    end
    if(N678) begin
      { valid[142:142] } <= { N541 };
    end
    if(N677) begin
      { valid[141:141] } <= { N541 };
    end
    if(N676) begin
      { valid[140:140] } <= { N541 };
    end
    if(N675) begin
      { valid[139:139] } <= { N541 };
    end
    if(N674) begin
      { valid[138:138] } <= { N541 };
    end
    if(N673) begin
      { valid[137:137] } <= { N541 };
    end
    if(N672) begin
      { valid[136:136] } <= { N541 };
    end
    if(N671) begin
      { valid[135:135] } <= { N541 };
    end
    if(N670) begin
      { valid[134:134] } <= { N541 };
    end
    if(N669) begin
      { valid[133:133] } <= { N541 };
    end
    if(N668) begin
      { valid[132:132] } <= { N541 };
    end
    if(N667) begin
      { valid[131:131] } <= { N541 };
    end
    if(N666) begin
      { valid[130:130] } <= { N541 };
    end
    if(N665) begin
      { valid[129:129] } <= { N541 };
    end
    if(N664) begin
      { valid[128:128] } <= { N541 };
    end
    if(N663) begin
      { valid[127:127] } <= { N541 };
    end
    if(N662) begin
      { valid[126:126] } <= { N541 };
    end
    if(N661) begin
      { valid[125:125] } <= { N541 };
    end
    if(N660) begin
      { valid[124:124] } <= { N541 };
    end
    if(N659) begin
      { valid[123:123] } <= { N541 };
    end
    if(N658) begin
      { valid[122:122] } <= { N541 };
    end
    if(N657) begin
      { valid[121:121] } <= { N541 };
    end
    if(N656) begin
      { valid[120:120] } <= { N541 };
    end
    if(N655) begin
      { valid[119:119] } <= { N541 };
    end
    if(N654) begin
      { valid[118:118] } <= { N541 };
    end
    if(N653) begin
      { valid[117:117] } <= { N541 };
    end
    if(N652) begin
      { valid[116:116] } <= { N541 };
    end
    if(N651) begin
      { valid[115:115] } <= { N541 };
    end
    if(N650) begin
      { valid[114:114] } <= { N541 };
    end
    if(N649) begin
      { valid[113:113] } <= { N541 };
    end
    if(N648) begin
      { valid[112:112] } <= { N541 };
    end
    if(N647) begin
      { valid[111:111] } <= { N541 };
    end
    if(N646) begin
      { valid[110:110] } <= { N541 };
    end
    if(N645) begin
      { valid[109:109] } <= { N541 };
    end
    if(N644) begin
      { valid[108:108] } <= { N541 };
    end
    if(N643) begin
      { valid[107:107] } <= { N541 };
    end
    if(N642) begin
      { valid[106:106] } <= { N541 };
    end
    if(N641) begin
      { valid[105:105] } <= { N541 };
    end
    if(N640) begin
      { valid[104:104] } <= { N541 };
    end
    if(N639) begin
      { valid[103:103] } <= { N541 };
    end
    if(N638) begin
      { valid[102:102] } <= { N541 };
    end
    if(N637) begin
      { valid[101:101] } <= { N541 };
    end
    if(N636) begin
      { valid[100:100] } <= { N541 };
    end
    if(N635) begin
      { valid[99:99] } <= { N541 };
    end
    if(N634) begin
      { valid[98:98] } <= { N541 };
    end
    if(N633) begin
      { valid[97:97] } <= { N541 };
    end
    if(N632) begin
      { valid[96:96] } <= { N541 };
    end
    if(N631) begin
      { valid[95:95] } <= { N541 };
    end
    if(N630) begin
      { valid[94:94] } <= { N541 };
    end
    if(N629) begin
      { valid[93:93] } <= { N541 };
    end
    if(N628) begin
      { valid[92:92] } <= { N541 };
    end
    if(N627) begin
      { valid[91:91] } <= { N541 };
    end
    if(N626) begin
      { valid[90:90] } <= { N541 };
    end
    if(N625) begin
      { valid[89:89] } <= { N541 };
    end
    if(N624) begin
      { valid[88:88] } <= { N541 };
    end
    if(N623) begin
      { valid[87:87] } <= { N541 };
    end
    if(N622) begin
      { valid[86:86] } <= { N541 };
    end
    if(N621) begin
      { valid[85:85] } <= { N541 };
    end
    if(N620) begin
      { valid[84:84] } <= { N541 };
    end
    if(N619) begin
      { valid[83:83] } <= { N541 };
    end
    if(N618) begin
      { valid[82:82] } <= { N541 };
    end
    if(N617) begin
      { valid[81:81] } <= { N541 };
    end
    if(N616) begin
      { valid[80:80] } <= { N541 };
    end
    if(N615) begin
      { valid[79:79] } <= { N541 };
    end
    if(N614) begin
      { valid[78:78] } <= { N541 };
    end
    if(N613) begin
      { valid[77:77] } <= { N541 };
    end
    if(N612) begin
      { valid[76:76] } <= { N541 };
    end
    if(N611) begin
      { valid[75:75] } <= { N541 };
    end
    if(N610) begin
      { valid[74:74] } <= { N541 };
    end
    if(N609) begin
      { valid[73:73] } <= { N541 };
    end
    if(N608) begin
      { valid[72:72] } <= { N541 };
    end
    if(N607) begin
      { valid[71:71] } <= { N541 };
    end
    if(N606) begin
      { valid[70:70] } <= { N541 };
    end
    if(N605) begin
      { valid[69:69] } <= { N541 };
    end
    if(N604) begin
      { valid[68:68] } <= { N541 };
    end
    if(N603) begin
      { valid[67:67] } <= { N541 };
    end
    if(N602) begin
      { valid[66:66] } <= { N541 };
    end
    if(N601) begin
      { valid[65:65] } <= { N541 };
    end
    if(N600) begin
      { valid[64:64] } <= { N541 };
    end
    if(N599) begin
      { valid[63:63] } <= { N541 };
    end
    if(N598) begin
      { valid[62:62] } <= { N541 };
    end
    if(N597) begin
      { valid[61:61] } <= { N541 };
    end
    if(N596) begin
      { valid[60:60] } <= { N541 };
    end
    if(N595) begin
      { valid[59:59] } <= { N541 };
    end
    if(N594) begin
      { valid[58:58] } <= { N541 };
    end
    if(N593) begin
      { valid[57:57] } <= { N541 };
    end
    if(N592) begin
      { valid[56:56] } <= { N541 };
    end
    if(N591) begin
      { valid[55:55] } <= { N541 };
    end
    if(N590) begin
      { valid[54:54] } <= { N541 };
    end
    if(N589) begin
      { valid[53:53] } <= { N541 };
    end
    if(N588) begin
      { valid[52:52] } <= { N541 };
    end
    if(N587) begin
      { valid[51:51] } <= { N541 };
    end
    if(N586) begin
      { valid[50:50] } <= { N541 };
    end
    if(N585) begin
      { valid[49:49] } <= { N541 };
    end
    if(N584) begin
      { valid[48:48] } <= { N541 };
    end
    if(N583) begin
      { valid[47:47] } <= { N541 };
    end
    if(N582) begin
      { valid[46:46] } <= { N541 };
    end
    if(N581) begin
      { valid[45:45] } <= { N541 };
    end
    if(N580) begin
      { valid[44:44] } <= { N541 };
    end
    if(N579) begin
      { valid[43:43] } <= { N541 };
    end
    if(N578) begin
      { valid[42:42] } <= { N541 };
    end
    if(N577) begin
      { valid[41:41] } <= { N541 };
    end
    if(N576) begin
      { valid[40:40] } <= { N541 };
    end
    if(N575) begin
      { valid[39:39] } <= { N541 };
    end
    if(N574) begin
      { valid[38:38] } <= { N541 };
    end
    if(N573) begin
      { valid[37:37] } <= { N541 };
    end
    if(N572) begin
      { valid[36:36] } <= { N541 };
    end
    if(N571) begin
      { valid[35:35] } <= { N541 };
    end
    if(N570) begin
      { valid[34:34] } <= { N541 };
    end
    if(N569) begin
      { valid[33:33] } <= { N541 };
    end
    if(N568) begin
      { valid[32:32] } <= { N541 };
    end
    if(N567) begin
      { valid[31:31] } <= { N541 };
    end
    if(N566) begin
      { valid[30:30] } <= { N541 };
    end
    if(N565) begin
      { valid[29:29] } <= { N541 };
    end
    if(N564) begin
      { valid[28:28] } <= { N541 };
    end
    if(N563) begin
      { valid[27:27] } <= { N541 };
    end
    if(N562) begin
      { valid[26:26] } <= { N541 };
    end
    if(N561) begin
      { valid[25:25] } <= { N541 };
    end
    if(N560) begin
      { valid[24:24] } <= { N541 };
    end
    if(N559) begin
      { valid[23:23] } <= { N541 };
    end
    if(N558) begin
      { valid[22:22] } <= { N541 };
    end
    if(N557) begin
      { valid[21:21] } <= { N541 };
    end
    if(N556) begin
      { valid[20:20] } <= { N541 };
    end
    if(N555) begin
      { valid[19:19] } <= { N541 };
    end
    if(N554) begin
      { valid[18:18] } <= { N541 };
    end
    if(N553) begin
      { valid[17:17] } <= { N541 };
    end
    if(N552) begin
      { valid[16:16] } <= { N541 };
    end
    if(N551) begin
      { valid[15:15] } <= { N541 };
    end
    if(N550) begin
      { valid[14:14] } <= { N541 };
    end
    if(N549) begin
      { valid[13:13] } <= { N541 };
    end
    if(N548) begin
      { valid[12:12] } <= { N541 };
    end
    if(N547) begin
      { valid[11:11] } <= { N541 };
    end
    if(N546) begin
      { valid[10:10] } <= { N541 };
    end
    if(N545) begin
      { valid[9:9] } <= { N541 };
    end
    if(N544) begin
      { valid[8:8] } <= { N541 };
    end
    if(N543) begin
      { valid[7:7] } <= { N541 };
    end
    if(N542) begin
      { valid[6:6] } <= { N541 };
    end
    if(N540) begin
      { valid[5:5] } <= { N541 };
    end
    if(N539) begin
      { valid[4:4] } <= { N541 };
    end
    if(N538) begin
      { valid[3:3] } <= { N541 };
    end
    if(N537) begin
      { valid[2:2] } <= { N541 };
    end
    if(N536) begin
      { valid[1:1] } <= { N541 };
    end
    if(N535) begin
      { valid[0:0] } <= { N541 };
    end
    if(1'b1) begin
      read_valid_o <= N2080;
    end
  end


endmodule



module bp_fe_branch_predictor_eaddr_width_p64_btb_indx_width_p9_bht_indx_width_p5_ras_addr_width_p22
(
  clk_i,
  reset_i,
  attaboy_i,
  r_v_i,
  btb_r_v_i,
  w_v_i,
  pc_queue_i,
  pc_cmd_i,
  pc_fwd_i,
  branch_metadata_fwd_i,
  predict_o,
  pc_o,
  branch_metadata_fwd_o
);

  input [63:0] pc_queue_i;
  input [63:0] pc_cmd_i;
  input [63:0] pc_fwd_i;
  input [35:0] branch_metadata_fwd_i;
  output [63:0] pc_o;
  output [35:0] branch_metadata_fwd_o;
  input clk_i;
  input reset_i;
  input attaboy_i;
  input r_v_i;
  input btb_r_v_i;
  input w_v_i;
  output predict_o;
  wire [63:0] pc_o;
  wire [35:0] branch_metadata_fwd_o;
  wire predict_o,predict,read_valid;
  assign branch_metadata_fwd_o[0] = 1'b0;
  assign branch_metadata_fwd_o[1] = 1'b0;
  assign branch_metadata_fwd_o[2] = 1'b0;
  assign branch_metadata_fwd_o[3] = 1'b0;
  assign branch_metadata_fwd_o[4] = 1'b0;
  assign branch_metadata_fwd_o[5] = 1'b0;
  assign branch_metadata_fwd_o[6] = 1'b0;
  assign branch_metadata_fwd_o[7] = 1'b0;
  assign branch_metadata_fwd_o[8] = 1'b0;
  assign branch_metadata_fwd_o[9] = 1'b0;
  assign branch_metadata_fwd_o[10] = 1'b0;
  assign branch_metadata_fwd_o[11] = 1'b0;
  assign branch_metadata_fwd_o[12] = 1'b0;
  assign branch_metadata_fwd_o[13] = 1'b0;
  assign branch_metadata_fwd_o[14] = 1'b0;
  assign branch_metadata_fwd_o[15] = 1'b0;
  assign branch_metadata_fwd_o[16] = 1'b0;
  assign branch_metadata_fwd_o[17] = 1'b0;
  assign branch_metadata_fwd_o[18] = 1'b0;
  assign branch_metadata_fwd_o[19] = 1'b0;
  assign branch_metadata_fwd_o[20] = 1'b0;
  assign branch_metadata_fwd_o[21] = 1'b0;
  assign branch_metadata_fwd_o[35] = pc_fwd_i[8];
  assign branch_metadata_fwd_o[34] = pc_fwd_i[7];
  assign branch_metadata_fwd_o[33] = pc_fwd_i[6];
  assign branch_metadata_fwd_o[32] = pc_fwd_i[5];
  assign branch_metadata_fwd_o[26] = pc_fwd_i[4];
  assign branch_metadata_fwd_o[31] = pc_fwd_i[4];
  assign branch_metadata_fwd_o[25] = pc_fwd_i[3];
  assign branch_metadata_fwd_o[30] = pc_fwd_i[3];
  assign branch_metadata_fwd_o[24] = pc_fwd_i[2];
  assign branch_metadata_fwd_o[29] = pc_fwd_i[2];
  assign branch_metadata_fwd_o[23] = pc_fwd_i[1];
  assign branch_metadata_fwd_o[28] = pc_fwd_i[1];
  assign branch_metadata_fwd_o[22] = pc_fwd_i[0];
  assign branch_metadata_fwd_o[27] = pc_fwd_i[0];

  bp_fe_bht_bht_indx_width_p5
  bht_1
  (
    .clk_i(clk_i),
    .en_i(1'b1),
    .reset_i(reset_i),
    .idx_r_i(pc_fwd_i[4:0]),
    .idx_w_i(branch_metadata_fwd_i[26:22]),
    .r_v_i(r_v_i),
    .w_v_i(w_v_i),
    .correct_i(attaboy_i),
    .predict_o(predict)
  );


  bp_fe_btb_bp_fe_pc_gen_btb_idx_width_lp9_eaddr_width_p64
  btb_1
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .idx_w_i(branch_metadata_fwd_i[35:27]),
    .idx_r_i(pc_queue_i[8:0]),
    .r_v_i(btb_r_v_i),
    .w_v_i(w_v_i),
    .branch_target_i(pc_cmd_i),
    .branch_target_o(pc_o),
    .read_valid_o(read_valid)
  );

  assign predict_o = predict & read_valid;

endmodule



module bp_fe_pc_gen_39_22_64_9_5_22_32_10_80000124_1
(
  clk_i,
  reset_i,
  v_i,
  pc_gen_icache_o,
  pc_gen_icache_v_o,
  pc_gen_icache_ready_i,
  icache_pc_gen_i,
  icache_pc_gen_v_i,
  icache_pc_gen_ready_o,
  icache_miss_i,
  pc_gen_itlb_o,
  pc_gen_itlb_v_o,
  pc_gen_itlb_ready_i,
  pc_gen_fe_o,
  pc_gen_fe_v_o,
  pc_gen_fe_ready_i,
  fe_pc_gen_i,
  fe_pc_gen_v_i,
  fe_pc_gen_ready_o
);

  output [63:0] pc_gen_icache_o;
  input [95:0] icache_pc_gen_i;
  output [63:0] pc_gen_itlb_o;
  output [202:0] pc_gen_fe_o;
  input [101:0] fe_pc_gen_i;
  input clk_i;
  input reset_i;
  input v_i;
  input pc_gen_icache_ready_i;
  input icache_pc_gen_v_i;
  input icache_miss_i;
  input pc_gen_itlb_ready_i;
  input pc_gen_fe_ready_i;
  input fe_pc_gen_v_i;
  output pc_gen_icache_v_o;
  output icache_pc_gen_ready_o;
  output pc_gen_itlb_v_o;
  output pc_gen_fe_v_o;
  output fe_pc_gen_ready_o;
  wire [63:0] pc_gen_itlb_o,next_pc,btb_target;
  wire [202:0] pc_gen_fe_o;
  wire pc_gen_icache_v_o,icache_pc_gen_ready_o,pc_gen_itlb_v_o,pc_gen_fe_v_o,
  fe_pc_gen_ready_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,misalignment,N12,
  pc_gen_exception_exception_code__1_,pc_gen_fetch_branch_metadata_fwd__35_,
  pc_gen_fetch_branch_metadata_fwd__34_,pc_gen_fetch_branch_metadata_fwd__33_,
  pc_gen_fetch_branch_metadata_fwd__32_,pc_gen_fetch_branch_metadata_fwd__31_,
  pc_gen_fetch_branch_metadata_fwd__30_,pc_gen_fetch_branch_metadata_fwd__29_,
  pc_gen_fetch_branch_metadata_fwd__28_,pc_gen_fetch_branch_metadata_fwd__27_,pc_gen_fetch_branch_metadata_fwd__26_,
  pc_gen_fetch_branch_metadata_fwd__25_,pc_gen_fetch_branch_metadata_fwd__24_,
  pc_gen_fetch_branch_metadata_fwd__23_,pc_gen_fetch_branch_metadata_fwd__22_,
  pc_gen_fetch_branch_metadata_fwd__21_,pc_gen_fetch_branch_metadata_fwd__20_,
  pc_gen_fetch_branch_metadata_fwd__19_,pc_gen_fetch_branch_metadata_fwd__18_,
  pc_gen_fetch_branch_metadata_fwd__17_,pc_gen_fetch_branch_metadata_fwd__16_,
  pc_gen_fetch_branch_metadata_fwd__15_,pc_gen_fetch_branch_metadata_fwd__14_,
  pc_gen_fetch_branch_metadata_fwd__13_,pc_gen_fetch_branch_metadata_fwd__12_,
  pc_gen_fetch_branch_metadata_fwd__11_,pc_gen_fetch_branch_metadata_fwd__10_,
  pc_gen_fetch_branch_metadata_fwd__9_,pc_gen_fetch_branch_metadata_fwd__8_,pc_gen_fetch_branch_metadata_fwd__7_,
  pc_gen_fetch_branch_metadata_fwd__6_,pc_gen_fetch_branch_metadata_fwd__5_,
  pc_gen_fetch_branch_metadata_fwd__4_,pc_gen_fetch_branch_metadata_fwd__3_,
  pc_gen_fetch_branch_metadata_fwd__2_,pc_gen_fetch_branch_metadata_fwd__1_,
  pc_gen_fetch_branch_metadata_fwd__0_,N13,N14,N15,N16,N17,predict,scan_instr_is_compressed_,
  scan_instr_instr_scan_class__3_,scan_instr_instr_scan_class__2_,
  scan_instr_instr_scan_class__1_,scan_instr_instr_scan_class__0_,scan_instr_imm__63_,scan_instr_imm__62_,
  scan_instr_imm__61_,scan_instr_imm__60_,scan_instr_imm__59_,scan_instr_imm__58_,
  scan_instr_imm__57_,scan_instr_imm__56_,scan_instr_imm__55_,scan_instr_imm__54_,
  scan_instr_imm__53_,scan_instr_imm__52_,scan_instr_imm__51_,scan_instr_imm__50_,
  scan_instr_imm__49_,scan_instr_imm__48_,scan_instr_imm__47_,scan_instr_imm__46_,
  scan_instr_imm__45_,scan_instr_imm__44_,scan_instr_imm__43_,scan_instr_imm__42_,
  scan_instr_imm__41_,scan_instr_imm__40_,scan_instr_imm__39_,scan_instr_imm__38_,
  scan_instr_imm__37_,scan_instr_imm__36_,scan_instr_imm__35_,scan_instr_imm__34_,
  scan_instr_imm__33_,scan_instr_imm__32_,scan_instr_imm__31_,scan_instr_imm__30_,
  scan_instr_imm__29_,scan_instr_imm__28_,scan_instr_imm__27_,scan_instr_imm__26_,
  scan_instr_imm__25_,scan_instr_imm__24_,scan_instr_imm__23_,scan_instr_imm__22_,
  scan_instr_imm__21_,scan_instr_imm__20_,scan_instr_imm__19_,scan_instr_imm__18_,
  scan_instr_imm__17_,scan_instr_imm__16_,scan_instr_imm__15_,scan_instr_imm__14_,
  scan_instr_imm__13_,scan_instr_imm__12_,scan_instr_imm__11_,scan_instr_imm__10_,
  scan_instr_imm__9_,scan_instr_imm__8_,scan_instr_imm__7_,scan_instr_imm__6_,
  scan_instr_imm__5_,scan_instr_imm__4_,scan_instr_imm__3_,scan_instr_imm__2_,
  scan_instr_imm__1_,scan_instr_imm__0_,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,
  N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,
  N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,
  N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,
  N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,
  N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,
  N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,
  N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,
  N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,
  N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,
  N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,
  N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,
  N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,
  N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,
  N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,
  N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,
  N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,
  N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,
  N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,
  N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,
  N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,
  N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,
  N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,
  N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,
  N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,
  N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,
  N444,stalled_pc_redirect_n,N445,N446,N447,bht_r_v_branch_jalr_inst,N448,N449,N450,
  N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,
  N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,
  N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,
  N499,N500,N501,N502,N503,N504;
  reg btb_r_v_i,stalled_pc_redirect;
  reg [63:0] pc_gen_icache_o,last_pc,icache_miss_pc,pc_redirect;
  assign pc_gen_fe_o[0] = 1'b0;
  assign pc_gen_itlb_v_o = 1'b0;
  assign icache_pc_gen_ready_o = 1'b0;
  assign pc_gen_itlb_o[63] = pc_gen_icache_o[63];
  assign pc_gen_itlb_o[62] = pc_gen_icache_o[62];
  assign pc_gen_itlb_o[61] = pc_gen_icache_o[61];
  assign pc_gen_itlb_o[60] = pc_gen_icache_o[60];
  assign pc_gen_itlb_o[59] = pc_gen_icache_o[59];
  assign pc_gen_itlb_o[58] = pc_gen_icache_o[58];
  assign pc_gen_itlb_o[57] = pc_gen_icache_o[57];
  assign pc_gen_itlb_o[56] = pc_gen_icache_o[56];
  assign pc_gen_itlb_o[55] = pc_gen_icache_o[55];
  assign pc_gen_itlb_o[54] = pc_gen_icache_o[54];
  assign pc_gen_itlb_o[53] = pc_gen_icache_o[53];
  assign pc_gen_itlb_o[52] = pc_gen_icache_o[52];
  assign pc_gen_itlb_o[51] = pc_gen_icache_o[51];
  assign pc_gen_itlb_o[50] = pc_gen_icache_o[50];
  assign pc_gen_itlb_o[49] = pc_gen_icache_o[49];
  assign pc_gen_itlb_o[48] = pc_gen_icache_o[48];
  assign pc_gen_itlb_o[47] = pc_gen_icache_o[47];
  assign pc_gen_itlb_o[46] = pc_gen_icache_o[46];
  assign pc_gen_itlb_o[45] = pc_gen_icache_o[45];
  assign pc_gen_itlb_o[44] = pc_gen_icache_o[44];
  assign pc_gen_itlb_o[43] = pc_gen_icache_o[43];
  assign pc_gen_itlb_o[42] = pc_gen_icache_o[42];
  assign pc_gen_itlb_o[41] = pc_gen_icache_o[41];
  assign pc_gen_itlb_o[40] = pc_gen_icache_o[40];
  assign pc_gen_itlb_o[39] = pc_gen_icache_o[39];
  assign pc_gen_itlb_o[38] = pc_gen_icache_o[38];
  assign pc_gen_itlb_o[37] = pc_gen_icache_o[37];
  assign pc_gen_itlb_o[36] = pc_gen_icache_o[36];
  assign pc_gen_itlb_o[35] = pc_gen_icache_o[35];
  assign pc_gen_itlb_o[34] = pc_gen_icache_o[34];
  assign pc_gen_itlb_o[33] = pc_gen_icache_o[33];
  assign pc_gen_itlb_o[32] = pc_gen_icache_o[32];
  assign pc_gen_itlb_o[31] = pc_gen_icache_o[31];
  assign pc_gen_itlb_o[30] = pc_gen_icache_o[30];
  assign pc_gen_itlb_o[29] = pc_gen_icache_o[29];
  assign pc_gen_itlb_o[28] = pc_gen_icache_o[28];
  assign pc_gen_itlb_o[27] = pc_gen_icache_o[27];
  assign pc_gen_itlb_o[26] = pc_gen_icache_o[26];
  assign pc_gen_itlb_o[25] = pc_gen_icache_o[25];
  assign pc_gen_itlb_o[24] = pc_gen_icache_o[24];
  assign pc_gen_itlb_o[23] = pc_gen_icache_o[23];
  assign pc_gen_itlb_o[22] = pc_gen_icache_o[22];
  assign pc_gen_itlb_o[21] = pc_gen_icache_o[21];
  assign pc_gen_itlb_o[20] = pc_gen_icache_o[20];
  assign pc_gen_itlb_o[19] = pc_gen_icache_o[19];
  assign pc_gen_itlb_o[18] = pc_gen_icache_o[18];
  assign pc_gen_itlb_o[17] = pc_gen_icache_o[17];
  assign pc_gen_itlb_o[16] = pc_gen_icache_o[16];
  assign pc_gen_itlb_o[15] = pc_gen_icache_o[15];
  assign pc_gen_itlb_o[14] = pc_gen_icache_o[14];
  assign pc_gen_itlb_o[13] = pc_gen_icache_o[13];
  assign pc_gen_itlb_o[12] = pc_gen_icache_o[12];
  assign pc_gen_itlb_o[11] = pc_gen_icache_o[11];
  assign pc_gen_itlb_o[10] = pc_gen_icache_o[10];
  assign pc_gen_itlb_o[9] = pc_gen_icache_o[9];
  assign pc_gen_itlb_o[8] = pc_gen_icache_o[8];
  assign pc_gen_itlb_o[7] = pc_gen_icache_o[7];
  assign pc_gen_itlb_o[6] = pc_gen_icache_o[6];
  assign pc_gen_itlb_o[5] = pc_gen_icache_o[5];
  assign pc_gen_itlb_o[4] = pc_gen_icache_o[4];
  assign pc_gen_itlb_o[3] = pc_gen_icache_o[3];
  assign pc_gen_itlb_o[2] = pc_gen_icache_o[2];
  assign pc_gen_itlb_o[1] = pc_gen_icache_o[1];
  assign pc_gen_itlb_o[0] = pc_gen_icache_o[0];
  assign N443 = icache_pc_gen_i[63:0] != pc_redirect;
  assign N444 = icache_pc_gen_i[63:0] == pc_redirect;

  instr_scan_eaddr_width_p64_instr_width_p32
  instr_scan_1
  (
    .instr_i(icache_pc_gen_i[95:64]),
    .scan_o({ scan_instr_is_compressed_, scan_instr_instr_scan_class__3_, scan_instr_instr_scan_class__2_, scan_instr_instr_scan_class__1_, scan_instr_instr_scan_class__0_, scan_instr_imm__63_, scan_instr_imm__62_, scan_instr_imm__61_, scan_instr_imm__60_, scan_instr_imm__59_, scan_instr_imm__58_, scan_instr_imm__57_, scan_instr_imm__56_, scan_instr_imm__55_, scan_instr_imm__54_, scan_instr_imm__53_, scan_instr_imm__52_, scan_instr_imm__51_, scan_instr_imm__50_, scan_instr_imm__49_, scan_instr_imm__48_, scan_instr_imm__47_, scan_instr_imm__46_, scan_instr_imm__45_, scan_instr_imm__44_, scan_instr_imm__43_, scan_instr_imm__42_, scan_instr_imm__41_, scan_instr_imm__40_, scan_instr_imm__39_, scan_instr_imm__38_, scan_instr_imm__37_, scan_instr_imm__36_, scan_instr_imm__35_, scan_instr_imm__34_, scan_instr_imm__33_, scan_instr_imm__32_, scan_instr_imm__31_, scan_instr_imm__30_, scan_instr_imm__29_, scan_instr_imm__28_, scan_instr_imm__27_, scan_instr_imm__26_, scan_instr_imm__25_, scan_instr_imm__24_, scan_instr_imm__23_, scan_instr_imm__22_, scan_instr_imm__21_, scan_instr_imm__20_, scan_instr_imm__19_, scan_instr_imm__18_, scan_instr_imm__17_, scan_instr_imm__16_, scan_instr_imm__15_, scan_instr_imm__14_, scan_instr_imm__13_, scan_instr_imm__12_, scan_instr_imm__11_, scan_instr_imm__10_, scan_instr_imm__9_, scan_instr_imm__8_, scan_instr_imm__7_, scan_instr_imm__6_, scan_instr_imm__5_, scan_instr_imm__4_, scan_instr_imm__3_, scan_instr_imm__2_, scan_instr_imm__1_, scan_instr_imm__0_ })
  );


  bp_fe_branch_predictor_eaddr_width_p64_btb_indx_width_p9_bht_indx_width_p5_ras_addr_width_p22
  genblk1_branch_prediction_1
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .attaboy_i(fe_pc_gen_i[0]),
    .r_v_i(bht_r_v_branch_jalr_inst),
    .btb_r_v_i(btb_r_v_i),
    .w_v_i(fe_pc_gen_v_i),
    .pc_queue_i(last_pc),
    .pc_cmd_i(fe_pc_gen_i[101:38]),
    .pc_fwd_i(icache_pc_gen_i[63:0]),
    .branch_metadata_fwd_i(fe_pc_gen_i[37:2]),
    .predict_o(predict),
    .pc_o(btb_target),
    .branch_metadata_fwd_o({ pc_gen_fetch_branch_metadata_fwd__35_, pc_gen_fetch_branch_metadata_fwd__34_, pc_gen_fetch_branch_metadata_fwd__33_, pc_gen_fetch_branch_metadata_fwd__32_, pc_gen_fetch_branch_metadata_fwd__31_, pc_gen_fetch_branch_metadata_fwd__30_, pc_gen_fetch_branch_metadata_fwd__29_, pc_gen_fetch_branch_metadata_fwd__28_, pc_gen_fetch_branch_metadata_fwd__27_, pc_gen_fetch_branch_metadata_fwd__26_, pc_gen_fetch_branch_metadata_fwd__25_, pc_gen_fetch_branch_metadata_fwd__24_, pc_gen_fetch_branch_metadata_fwd__23_, pc_gen_fetch_branch_metadata_fwd__22_, pc_gen_fetch_branch_metadata_fwd__21_, pc_gen_fetch_branch_metadata_fwd__20_, pc_gen_fetch_branch_metadata_fwd__19_, pc_gen_fetch_branch_metadata_fwd__18_, pc_gen_fetch_branch_metadata_fwd__17_, pc_gen_fetch_branch_metadata_fwd__16_, pc_gen_fetch_branch_metadata_fwd__15_, pc_gen_fetch_branch_metadata_fwd__14_, pc_gen_fetch_branch_metadata_fwd__13_, pc_gen_fetch_branch_metadata_fwd__12_, pc_gen_fetch_branch_metadata_fwd__11_, pc_gen_fetch_branch_metadata_fwd__10_, pc_gen_fetch_branch_metadata_fwd__9_, pc_gen_fetch_branch_metadata_fwd__8_, pc_gen_fetch_branch_metadata_fwd__7_, pc_gen_fetch_branch_metadata_fwd__6_, pc_gen_fetch_branch_metadata_fwd__5_, pc_gen_fetch_branch_metadata_fwd__4_, pc_gen_fetch_branch_metadata_fwd__3_, pc_gen_fetch_branch_metadata_fwd__2_, pc_gen_fetch_branch_metadata_fwd__1_, pc_gen_fetch_branch_metadata_fwd__0_ })
  );

  assign N448 = ~scan_instr_instr_scan_class__0_;
  assign N449 = scan_instr_instr_scan_class__2_ | scan_instr_instr_scan_class__3_;
  assign N450 = scan_instr_instr_scan_class__1_ | N449;
  assign N451 = N448 | N450;
  assign N452 = ~N451;
  assign N453 = scan_instr_instr_scan_class__2_ | scan_instr_instr_scan_class__3_;
  assign N454 = scan_instr_instr_scan_class__1_ | N453;
  assign N455 = scan_instr_instr_scan_class__0_ | N454;
  assign N456 = ~N455;
  assign N457 = ~pc_gen_fe_o[202];
  assign N458 = N9 | N8;
  assign N459 = N10 | N458;
  assign N460 = N11 | N459;
  assign N461 = ~N460;
  assign N462 = ~N9;
  assign N463 = N462 | N8;
  assign N464 = N10 | N463;
  assign N465 = N11 | N464;
  assign N466 = ~N465;
  assign N467 = ~N8;
  assign N468 = N9 | N467;
  assign N469 = N10 | N468;
  assign N470 = N11 | N469;
  assign N471 = ~N470;
  assign N472 = N462 | N467;
  assign N473 = N10 | N472;
  assign N474 = N11 | N473;
  assign N475 = ~N474;
  assign N476 = ~scan_instr_instr_scan_class__1_;
  assign N477 = scan_instr_instr_scan_class__2_ | scan_instr_instr_scan_class__3_;
  assign N478 = N476 | N477;
  assign N479 = scan_instr_instr_scan_class__0_ | N478;
  assign N480 = ~N479;
  assign N481 = scan_instr_instr_scan_class__2_ | scan_instr_instr_scan_class__3_;
  assign N482 = scan_instr_instr_scan_class__1_ | N481;
  assign N483 = scan_instr_instr_scan_class__0_ | N482;
  assign N484 = ~N483;
  assign N485 = scan_instr_instr_scan_class__2_ | scan_instr_instr_scan_class__3_;
  assign N486 = scan_instr_instr_scan_class__1_ | N485;
  assign N487 = N448 | N486;
  assign N488 = ~N487;
  assign { N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156 } = pc_gen_icache_o + { 1'b1, 1'b0, 1'b0 };
  assign { N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27 } = icache_pc_gen_i[63:0] + { scan_instr_imm__63_, scan_instr_imm__62_, scan_instr_imm__61_, scan_instr_imm__60_, scan_instr_imm__59_, scan_instr_imm__58_, scan_instr_imm__57_, scan_instr_imm__56_, scan_instr_imm__55_, scan_instr_imm__54_, scan_instr_imm__53_, scan_instr_imm__52_, scan_instr_imm__51_, scan_instr_imm__50_, scan_instr_imm__49_, scan_instr_imm__48_, scan_instr_imm__47_, scan_instr_imm__46_, scan_instr_imm__45_, scan_instr_imm__44_, scan_instr_imm__43_, scan_instr_imm__42_, scan_instr_imm__41_, scan_instr_imm__40_, scan_instr_imm__39_, scan_instr_imm__38_, scan_instr_imm__37_, scan_instr_imm__36_, scan_instr_imm__35_, scan_instr_imm__34_, scan_instr_imm__33_, scan_instr_imm__32_, scan_instr_imm__31_, scan_instr_imm__30_, scan_instr_imm__29_, scan_instr_imm__28_, scan_instr_imm__27_, scan_instr_imm__26_, scan_instr_imm__25_, scan_instr_imm__24_, scan_instr_imm__23_, scan_instr_imm__22_, scan_instr_imm__21_, scan_instr_imm__20_, scan_instr_imm__19_, scan_instr_imm__18_, scan_instr_imm__17_, scan_instr_imm__16_, scan_instr_imm__15_, scan_instr_imm__14_, scan_instr_imm__13_, scan_instr_imm__12_, scan_instr_imm__11_, scan_instr_imm__10_, scan_instr_imm__9_, scan_instr_imm__8_, scan_instr_imm__7_, scan_instr_imm__6_, scan_instr_imm__5_, scan_instr_imm__4_, scan_instr_imm__3_, scan_instr_imm__2_, scan_instr_imm__1_, scan_instr_imm__0_ };
  assign { N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92 } = icache_pc_gen_i[63:0] + { scan_instr_imm__63_, scan_instr_imm__62_, scan_instr_imm__61_, scan_instr_imm__60_, scan_instr_imm__59_, scan_instr_imm__58_, scan_instr_imm__57_, scan_instr_imm__56_, scan_instr_imm__55_, scan_instr_imm__54_, scan_instr_imm__53_, scan_instr_imm__52_, scan_instr_imm__51_, scan_instr_imm__50_, scan_instr_imm__49_, scan_instr_imm__48_, scan_instr_imm__47_, scan_instr_imm__46_, scan_instr_imm__45_, scan_instr_imm__44_, scan_instr_imm__43_, scan_instr_imm__42_, scan_instr_imm__41_, scan_instr_imm__40_, scan_instr_imm__39_, scan_instr_imm__38_, scan_instr_imm__37_, scan_instr_imm__36_, scan_instr_imm__35_, scan_instr_imm__34_, scan_instr_imm__33_, scan_instr_imm__32_, scan_instr_imm__31_, scan_instr_imm__30_, scan_instr_imm__29_, scan_instr_imm__28_, scan_instr_imm__27_, scan_instr_imm__26_, scan_instr_imm__25_, scan_instr_imm__24_, scan_instr_imm__23_, scan_instr_imm__22_, scan_instr_imm__21_, scan_instr_imm__20_, scan_instr_imm__19_, scan_instr_imm__18_, scan_instr_imm__17_, scan_instr_imm__16_, scan_instr_imm__15_, scan_instr_imm__14_, scan_instr_imm__13_, scan_instr_imm__12_, scan_instr_imm__11_, scan_instr_imm__10_, scan_instr_imm__9_, scan_instr_imm__8_, scan_instr_imm__7_, scan_instr_imm__6_, scan_instr_imm__5_, scan_instr_imm__4_, scan_instr_imm__3_, scan_instr_imm__2_, scan_instr_imm__1_, scan_instr_imm__0_ };
  assign pc_gen_fe_o[132:1] = (N0)? { icache_pc_gen_i[63:0], icache_pc_gen_i[95:64], pc_gen_fetch_branch_metadata_fwd__35_, pc_gen_fetch_branch_metadata_fwd__34_, pc_gen_fetch_branch_metadata_fwd__33_, pc_gen_fetch_branch_metadata_fwd__32_, pc_gen_fetch_branch_metadata_fwd__31_, pc_gen_fetch_branch_metadata_fwd__30_, pc_gen_fetch_branch_metadata_fwd__29_, pc_gen_fetch_branch_metadata_fwd__28_, pc_gen_fetch_branch_metadata_fwd__27_, pc_gen_fetch_branch_metadata_fwd__26_, pc_gen_fetch_branch_metadata_fwd__25_, pc_gen_fetch_branch_metadata_fwd__24_, pc_gen_fetch_branch_metadata_fwd__23_, pc_gen_fetch_branch_metadata_fwd__22_, pc_gen_fetch_branch_metadata_fwd__21_, pc_gen_fetch_branch_metadata_fwd__20_, pc_gen_fetch_branch_metadata_fwd__19_, pc_gen_fetch_branch_metadata_fwd__18_, pc_gen_fetch_branch_metadata_fwd__17_, pc_gen_fetch_branch_metadata_fwd__16_, pc_gen_fetch_branch_metadata_fwd__15_, pc_gen_fetch_branch_metadata_fwd__14_, pc_gen_fetch_branch_metadata_fwd__13_, pc_gen_fetch_branch_metadata_fwd__12_, pc_gen_fetch_branch_metadata_fwd__11_, pc_gen_fetch_branch_metadata_fwd__10_, pc_gen_fetch_branch_metadata_fwd__9_, pc_gen_fetch_branch_metadata_fwd__8_, pc_gen_fetch_branch_metadata_fwd__7_, pc_gen_fetch_branch_metadata_fwd__6_, pc_gen_fetch_branch_metadata_fwd__5_, pc_gen_fetch_branch_metadata_fwd__4_, pc_gen_fetch_branch_metadata_fwd__3_, pc_gen_fetch_branch_metadata_fwd__2_, pc_gen_fetch_branch_metadata_fwd__1_, pc_gen_fetch_branch_metadata_fwd__0_ } :
                              (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, pc_gen_exception_exception_code__1_, pc_gen_exception_exception_code__1_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N457;
  assign N1 = pc_gen_fe_o[202];
  assign pc_gen_fe_v_o = (N2)? 1'b0 :
                         (N3)? N15 : 1'b0;
  assign N2 = N14;
  assign N3 = N13;
  assign fe_pc_gen_ready_o = (N2)? 1'b0 :
                             (N3)? fe_pc_gen_v_i : 1'b0;
  assign pc_gen_icache_v_o = (N2)? 1'b0 :
                             (N3)? N16 : 1'b0;
  assign next_pc = (N4)? icache_miss_pc :
                   (N221)? fe_pc_gen_i[101:38] :
                   (N224)? btb_target :
                   (N227)? { N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27 } :
                   (N230)? { N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92 } :
                   (N25)? { N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156 } : 1'b0;
  assign N4 = icache_miss_i;
  assign { N241, N239 } = (N5)? { 1'b1, 1'b1 } :
                          (N435)? { 1'b1, 1'b1 } :
                          (N438)? { 1'b1, 1'b1 } :
                          (N441)? { 1'b1, 1'b1 } :
                          (N238)? { 1'b0, 1'b0 } : 1'b0;
  assign N5 = N234;
  assign { N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N240 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } :
                                                                                                                                                                                                                                                                                                                                                                                                              (N435)? pc_redirect :
                                                                                                                                                                                                                                                                                                                                                                                                              (N438)? next_pc :
                                                                                                                                                                                                                                                                                                                                                                                                              (N441)? icache_miss_pc : 1'b0;
  assign { N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                                                                                                                                                                                                                                                                              (N435)? pc_gen_icache_o :
                                                                                                                                                                                                                                                                                                                                                                                                              (N438)? pc_gen_icache_o :
                                                                                                                                                                                                                                                                                                                                                                                                              (N441)? pc_gen_icache_o : 1'b0;
  assign { N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                                                                                                                                                                                                                                                                              (N435)? last_pc :
                                                                                                                                                                                                                                                                                                                                                                                                              (N438)? last_pc :
                                                                                                                                                                                                                                                                                                                                                                                                              (N441)? last_pc : 1'b0;
  assign N433 = (N5)? 1'b0 :
                (N435)? pc_gen_icache_v_o :
                (N438)? pc_gen_icache_v_o :
                (N441)? pc_gen_icache_v_o : 1'b0;
  assign N447 = (N6)? 1'b0 :
                (N7)? stalled_pc_redirect_n : 1'b0;
  assign N6 = N446;
  assign N7 = N445;
  assign N8 = ~fe_pc_gen_i[41];
  assign N9 = ~fe_pc_gen_i[40];
  assign N10 = ~fe_pc_gen_i[39];
  assign N11 = ~fe_pc_gen_i[38];
  assign misalignment = N492 & N475;
  assign N492 = N491 & N471;
  assign N491 = N490 & N466;
  assign N490 = N489 & N461;
  assign N489 = fe_pc_gen_v_i & fe_pc_gen_i[1];
  assign pc_gen_fe_o[202] = misalignment;
  assign N12 = ~misalignment;
  assign pc_gen_exception_exception_code__1_ = N12;
  assign N13 = ~reset_i;
  assign N14 = reset_i;
  assign N15 = N493 & N494;
  assign N493 = pc_gen_fe_ready_i & icache_pc_gen_v_i;
  assign N494 = ~icache_miss_i;
  assign N16 = pc_gen_fe_ready_i & N494;
  assign N17 = fe_pc_gen_i[1] & fe_pc_gen_v_i;
  assign N18 = N495 & N488;
  assign N495 = predict & icache_pc_gen_v_i;
  assign N19 = N496 & N484;
  assign N496 = predict & icache_pc_gen_v_i;
  assign N20 = icache_pc_gen_v_i & N480;
  assign N21 = N17 | icache_miss_i;
  assign N22 = N18 | N21;
  assign N23 = N19 | N22;
  assign N24 = N20 | N23;
  assign N25 = ~N24;
  assign N26 = N227;
  assign N91 = N230;
  assign N220 = ~icache_miss_i;
  assign N221 = N17 & N220;
  assign N222 = ~N17;
  assign N223 = N220 & N222;
  assign N224 = N18 & N223;
  assign N225 = ~N18;
  assign N226 = N223 & N225;
  assign N227 = N19 & N226;
  assign N228 = ~N19;
  assign N229 = N226 & N228;
  assign N230 = N20 & N229;
  assign N231 = stalled_pc_redirect & icache_miss_i;
  assign N232 = pc_gen_icache_ready_i & pc_gen_fe_ready_i;
  assign N233 = icache_miss_i & N497;
  assign N497 = ~pc_gen_icache_ready_i;
  assign N234 = reset_i;
  assign N235 = N231 | N234;
  assign N236 = N232 | N235;
  assign N237 = N233 | N236;
  assign N238 = ~N237;
  assign N434 = ~N234;
  assign N435 = N231 & N434;
  assign N436 = ~N231;
  assign N437 = N434 & N436;
  assign N438 = N232 & N437;
  assign N439 = ~N232;
  assign N440 = N437 & N439;
  assign N441 = N233 & N440;
  assign N442 = fe_pc_gen_v_i & fe_pc_gen_i[1];
  assign stalled_pc_redirect_n = N500 | N503;
  assign N500 = N498 | N499;
  assign N498 = fe_pc_gen_v_i & fe_pc_gen_i[1];
  assign N499 = stalled_pc_redirect & N443;
  assign N503 = N501 & N502;
  assign N501 = stalled_pc_redirect & N444;
  assign N502 = ~pc_gen_fe_v_o;
  assign N445 = ~reset_i;
  assign N446 = reset_i;
  assign bht_r_v_branch_jalr_inst = icache_pc_gen_v_i & N504;
  assign N504 = N452 | N456;

  always @(posedge clk_i) begin
    if(N239) begin
      btb_r_v_i <= N433;
      { pc_gen_icache_o[0:0] } <= { N240 };
      { last_pc[63:30] } <= { N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335 };
      { icache_miss_pc[63:0] } <= { N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369 };
    end
    if(N241) begin
      { pc_gen_icache_o[63:1] } <= { N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242 };
      { last_pc[29:0] } <= { N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305 };
    end
    if(N442) begin
      { pc_redirect[63:0] } <= { fe_pc_gen_i[101:38] };
    end
    if(1'b1) begin
      stalled_pc_redirect <= N447;
    end
  end


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p96_els_p64
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [95:0] data_i;
  input [5:0] addr_i;
  input [95:0] w_mask_i;
  output [95:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [95:0] data_o;

  hard_mem_1rw_bit_mask_d64_w96_wrapper
  macro_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  addr_i,
  data_i,
  write_mask_i,
  data_o
);

  input [8:0] addr_i;
  input [63:0] data_i;
  input [7:0] write_mask_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [63:0] data_o;

  hard_mem_1rw_byte_mask_d512_w64_wrapper
  macro_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .w_i(w_i),
    .addr_i(addr_i),
    .data_i(data_i),
    .write_mask_i(write_mask_i),
    .data_o(data_o)
  );


endmodule



module bsg_scan_width_p8_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [7:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__7_,t_1__6_,
  t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__7_ = i[0] | 1'b0;
  assign t_1__6_ = i[1] | i[0];
  assign t_1__5_ = i[2] | i[1];
  assign t_1__4_ = i[3] | i[2];
  assign t_1__3_ = i[4] | i[3];
  assign t_1__2_ = i[5] | i[4];
  assign t_1__1_ = i[6] | i[5];
  assign t_1__0_ = i[7] | i[6];
  assign t_2__7_ = t_1__7_ | 1'b0;
  assign t_2__6_ = t_1__6_ | 1'b0;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign o[0] = t_2__7_ | 1'b0;
  assign o[1] = t_2__6_ | 1'b0;
  assign o[2] = t_2__5_ | 1'b0;
  assign o[3] = t_2__4_ | 1'b0;
  assign o[4] = t_2__3_ | t_2__7_;
  assign o[5] = t_2__2_ | t_2__6_;
  assign o[6] = t_2__1_ | t_2__5_;
  assign o[7] = t_2__0_ | t_2__4_;

endmodule



module bsg_priority_encode_one_hot_out_width_p8_lo_to_hi_p1
(
  i,
  o
);

  input [7:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire N0,N1,N2,N3,N4,N5,N6;
  wire [7:1] scan_lo;

  bsg_scan_width_p8_or_p1_lo_to_hi_p1
  scan
  (
    .i(i),
    .o({ scan_lo, o[0:0] })
  );

  assign o[7] = scan_lo[7] & N0;
  assign N0 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N1;
  assign N1 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N2;
  assign N2 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N3;
  assign N3 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N4;
  assign N4 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N5;
  assign N5 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N6;
  assign N6 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p1
(
  i,
  addr_o,
  v_o
);

  input [0:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign v_o = i[0];
  assign addr_o[0] = 1'b0;

endmodule



module bsg_encode_one_hot_width_p2
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o,aligned_vs;
  wire v_o;
  wire [1:0] aligned_addrs;

  bsg_encode_one_hot_width_p1
  aligned_left
  (
    .i(i[0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p1
  aligned_right
  (
    .i(i[1]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[0])
  );

  assign v_o = addr_o[0] | aligned_vs[0];

endmodule



module bsg_encode_one_hot_width_p4
(
  i,
  addr_o,
  v_o
);

  input [3:0] i;
  output [1:0] addr_o;
  output v_o;
  wire [1:0] addr_o,aligned_addrs;
  wire v_o;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p2
  aligned_left
  (
    .i(i[1:0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p2
  aligned_right
  (
    .i(i[3:2]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[1])
  );

  assign v_o = addr_o[1] | aligned_vs[0];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[1];

endmodule



module bsg_encode_one_hot_width_p8_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [3:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p4
  aligned_left
  (
    .i(i[3:0]),
    .addr_o(aligned_addrs[1:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p4
  aligned_right
  (
    .i(i[7:4]),
    .addr_o(aligned_addrs[3:2]),
    .v_o(addr_o[2])
  );

  assign v_o = addr_o[2] | aligned_vs[0];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[3];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[2];

endmodule



module bsg_priority_encode_width_p8_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [7:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p8_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo)
  );


  bsg_encode_one_hot_width_p8_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o),
    .v_o(v_o)
  );


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p7_els_p64
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [6:0] data_i;
  input [5:0] addr_i;
  input [6:0] w_mask_i;
  output [6:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [6:0] data_o;

  hard_mem_1rw_bit_mask_d64_w7_wrapper
  macro_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_scan_7_1_1
(
  i,
  o
);

  input [6:0] i;
  output [6:0] o;
  wire [6:0] o;
  wire t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__6_,t_1__5_,t_1__4_,
  t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__6_ = i[0] | 1'b0;
  assign t_1__5_ = i[1] | i[0];
  assign t_1__4_ = i[2] | i[1];
  assign t_1__3_ = i[3] | i[2];
  assign t_1__2_ = i[4] | i[3];
  assign t_1__1_ = i[5] | i[4];
  assign t_1__0_ = i[6] | i[5];
  assign t_2__6_ = t_1__6_ | 1'b0;
  assign t_2__5_ = t_1__5_ | 1'b0;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign o[0] = t_2__6_ | 1'b0;
  assign o[1] = t_2__5_ | 1'b0;
  assign o[2] = t_2__4_ | 1'b0;
  assign o[3] = t_2__3_ | 1'b0;
  assign o[4] = t_2__2_ | t_2__6_;
  assign o[5] = t_2__1_ | t_2__5_;
  assign o[6] = t_2__0_ | t_2__4_;

endmodule



module bsg_priority_encode_one_hot_out_7_1
(
  i,
  o
);

  input [6:0] i;
  output [6:0] o;
  wire [6:0] o;
  wire N0,N1,N2,N3,N4,N5;
  wire [6:1] scan_lo;

  bsg_scan_7_1_1
  scan
  (
    .i(i),
    .o({ scan_lo, o[0:0] })
  );

  assign o[6] = scan_lo[6] & N0;
  assign N0 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N1;
  assign N1 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N2;
  assign N2 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N3;
  assign N3 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N4;
  assign N4 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N5;
  assign N5 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p8
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [3:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p4
  aligned_left
  (
    .i(i[3:0]),
    .addr_o(aligned_addrs[1:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p4
  aligned_right
  (
    .i(i[7:4]),
    .addr_o(aligned_addrs[3:2]),
    .v_o(addr_o[2])
  );

  assign v_o = addr_o[2] | aligned_vs[0];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[3];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[2];

endmodule



module bsg_encode_one_hot_7_1
(
  i,
  addr_o,
  v_o
);

  input [6:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;

  bsg_encode_one_hot_width_p8
  unaligned_align
  (
    .i({ 1'b0, i }),
    .addr_o(addr_o),
    .v_o(v_o)
  );


endmodule



module bsg_priority_encode_7_1
(
  i,
  addr_o,
  v_o
);

  input [6:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [6:0] enc_lo;

  bsg_priority_encode_one_hot_out_7_1
  a
  (
    .i(i),
    .o(enc_lo)
  );


  bsg_encode_one_hot_7_1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o),
    .v_o(v_o)
  );


endmodule



module bsg_lru_pseudo_tree_encode_ways_p8
(
  lru_i,
  way_id_o
);

  input [6:0] lru_i;
  output [2:0] way_id_o;
  wire [2:0] way_id_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,pe_o_2__2_,pe_o_2__1_,pe_o_2__0_,
  pe_o_1__2_,pe_o_1__1_,pe_o_1__0_,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,
  pe_i_2__6_,pe_i_2__5_,pe_i_2__4_,pe_i_2__3_,pe_i_2__2_,pe_i_2__1_,pe_i_2__0_,pe_i_1__6_,
  pe_i_1__5_,pe_i_1__4_,pe_i_1__3_,pe_i_1__2_,pe_i_1__1_,pe_i_1__0_,N44,N45,N46,
  N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
  N67;
  wire [6:1] mask;

  bsg_priority_encode_7_1
  rof2_1__fi3_pe
  (
    .i({ pe_i_1__6_, pe_i_1__5_, pe_i_1__4_, pe_i_1__3_, pe_i_1__2_, pe_i_1__1_, pe_i_1__0_ }),
    .addr_o({ pe_o_1__2_, pe_o_1__1_, pe_o_1__0_ })
  );

  assign { N64, N63, N62, N61, N60, N59, N58 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << { pe_o_1__2_, pe_o_1__1_, pe_o_1__0_ };

  bsg_priority_encode_7_1
  rof2_2__fi3_pe
  (
    .i({ pe_i_2__6_, pe_i_2__5_, pe_i_2__4_, pe_i_2__3_, pe_i_2__2_, pe_i_2__1_, pe_i_2__0_ }),
    .addr_o({ pe_o_2__2_, pe_o_2__1_, pe_o_2__0_ })
  );

  assign N44 = N0 & N1 & N2;
  assign N0 = ~pe_o_1__2_;
  assign N1 = ~pe_o_1__0_;
  assign N2 = ~pe_o_1__1_;
  assign N45 = pe_o_1__2_ & N3 & N4;
  assign N3 = ~pe_o_1__0_;
  assign N4 = ~pe_o_1__1_;
  assign N46 = N5 & pe_o_1__0_ & N6;
  assign N5 = ~pe_o_1__2_;
  assign N6 = ~pe_o_1__1_;
  assign N48 = N7 & N8 & pe_o_1__1_;
  assign N7 = ~pe_o_1__2_;
  assign N8 = ~pe_o_1__0_;
  assign N50 = pe_o_1__0_ & pe_o_1__1_;
  assign N47 = pe_o_1__2_ & pe_o_1__0_;
  assign N49 = pe_o_1__2_ & pe_o_1__1_;
  assign N51 = N9 & N10 & N11;
  assign N9 = ~pe_o_2__2_;
  assign N10 = ~pe_o_2__0_;
  assign N11 = ~pe_o_2__1_;
  assign N52 = pe_o_2__2_ & N12 & N13;
  assign N12 = ~pe_o_2__0_;
  assign N13 = ~pe_o_2__1_;
  assign N53 = N14 & pe_o_2__0_ & N15;
  assign N14 = ~pe_o_2__2_;
  assign N15 = ~pe_o_2__1_;
  assign N55 = N16 & N17 & pe_o_2__1_;
  assign N16 = ~pe_o_2__2_;
  assign N17 = ~pe_o_2__0_;
  assign N57 = pe_o_2__0_ & pe_o_2__1_;
  assign N54 = pe_o_2__2_ & pe_o_2__0_;
  assign N56 = pe_o_2__2_ & pe_o_2__1_;
  assign way_id_o[1] = (N18)? lru_i[0] :
                       (N19)? lru_i[1] :
                       (N20)? lru_i[2] :
                       (N21)? lru_i[3] :
                       (N22)? lru_i[4] :
                       (N23)? lru_i[5] :
                       (N24)? lru_i[6] : 1'b0;
  assign N18 = N44;
  assign N19 = N46;
  assign N20 = N48;
  assign N21 = N50;
  assign N22 = N45;
  assign N23 = N47;
  assign N24 = N49;
  assign way_id_o[0] = (N25)? lru_i[0] :
                       (N26)? lru_i[1] :
                       (N27)? lru_i[2] :
                       (N28)? lru_i[3] :
                       (N29)? lru_i[4] :
                       (N30)? lru_i[5] :
                       (N31)? lru_i[6] : 1'b0;
  assign N25 = N51;
  assign N26 = N53;
  assign N27 = N55;
  assign N28 = N57;
  assign N29 = N52;
  assign N30 = N54;
  assign N31 = N56;
  assign way_id_o[2] = (N37)? lru_i[0] :
                       (N39)? lru_i[1] :
                       (N41)? lru_i[2] :
                       (N43)? lru_i[3] :
                       (N38)? lru_i[4] :
                       (N40)? lru_i[5] :
                       (N42)? lru_i[6] : 1'b0;
  assign mask[1] = 1'b1 & N65;
  assign N65 = ~lru_i[0];
  assign mask[2] = 1'b1 & lru_i[0];
  assign mask[3] = mask[1] & N66;
  assign N66 = ~lru_i[1];
  assign mask[4] = mask[1] & lru_i[1];
  assign mask[5] = mask[2] & N67;
  assign N67 = ~lru_i[2];
  assign mask[6] = mask[2] & lru_i[2];
  assign N32 = N36 & N36;
  assign N33 = N36 & 1'b0;
  assign N34 = 1'b0 & N36;
  assign N35 = 1'b0 & 1'b0;
  assign N36 = ~1'b0;
  assign N37 = N32 & N36;
  assign N38 = N32 & 1'b0;
  assign N39 = N34 & N36;
  assign N40 = N34 & 1'b0;
  assign N41 = N33 & N36;
  assign N42 = N33 & 1'b0;
  assign N43 = N35 & N36;
  assign pe_i_1__6_ = mask[6] ^ 1'b0;
  assign pe_i_1__5_ = mask[5] ^ 1'b0;
  assign pe_i_1__4_ = mask[4] ^ 1'b0;
  assign pe_i_1__3_ = mask[3] ^ 1'b0;
  assign pe_i_1__2_ = mask[2] ^ 1'b0;
  assign pe_i_1__1_ = mask[1] ^ 1'b0;
  assign pe_i_1__0_ = 1'b1 ^ 1'b1;
  assign pe_i_2__6_ = pe_i_1__6_ ^ N64;
  assign pe_i_2__5_ = pe_i_1__5_ ^ N63;
  assign pe_i_2__4_ = pe_i_1__4_ ^ N62;
  assign pe_i_2__3_ = pe_i_1__3_ ^ N61;
  assign pe_i_2__2_ = pe_i_1__2_ ^ N60;
  assign pe_i_2__1_ = pe_i_1__1_ ^ N59;
  assign pe_i_2__0_ = pe_i_1__0_ ^ N58;

endmodule



module bp_fe_lce_req_data_width_p64_paddr_width_p22_num_cce_p1_num_lce_p2_sets_p64_ways_p8
(
  clk_i,
  reset_i,
  id_i,
  miss_i,
  miss_addr_i,
  lru_way_i,
  cache_miss_o,
  miss_addr_o,
  tr_data_received_i,
  cce_data_received_i,
  set_tag_received_i,
  set_tag_wakeup_received_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_yumi_i
);

  input [0:0] id_i;
  input [21:0] miss_addr_i;
  input [2:0] lru_way_i;
  output [21:0] miss_addr_o;
  output [96:0] lce_req_o;
  output [25:0] lce_resp_o;
  input clk_i;
  input reset_i;
  input miss_i;
  input tr_data_received_i;
  input cce_data_received_i;
  input set_tag_received_i;
  input set_tag_wakeup_received_i;
  input lce_req_ready_i;
  input lce_resp_yumi_i;
  output cache_miss_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  wire [96:0] lce_req_o;
  wire cache_miss_o,lce_req_v_o,lce_resp_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,
  tr_data_received_n,cce_data_received_n,set_tag_received_n,tr_data_received,
  cce_data_received,set_tag_received,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,
  N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,
  N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,
  N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,
  N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100;
  wire [2:0] state_n;
  reg [25:0] lce_resp_o;
  reg [2:0] lru_way_r,state_r;
  reg lru_flopped_r,tr_data_received_r,cce_data_received_r,set_tag_received_r;
  reg [21:0] miss_addr_o;
  assign lce_resp_o[23] = 1'b1;
  assign lce_req_o[29] = 1'b1;
  assign lce_req_o[0] = 1'b0;
  assign lce_req_o[1] = 1'b0;
  assign lce_req_o[2] = 1'b0;
  assign lce_req_o[3] = 1'b0;
  assign lce_req_o[30] = 1'b0;
  assign lce_req_o[33] = 1'b0;
  assign lce_req_o[34] = 1'b0;
  assign lce_req_o[35] = 1'b0;
  assign lce_req_o[36] = 1'b0;
  assign lce_req_o[37] = 1'b0;
  assign lce_req_o[38] = 1'b0;
  assign lce_req_o[39] = 1'b0;
  assign lce_req_o[40] = 1'b0;
  assign lce_req_o[41] = 1'b0;
  assign lce_req_o[42] = 1'b0;
  assign lce_req_o[43] = 1'b0;
  assign lce_req_o[44] = 1'b0;
  assign lce_req_o[45] = 1'b0;
  assign lce_req_o[46] = 1'b0;
  assign lce_req_o[47] = 1'b0;
  assign lce_req_o[48] = 1'b0;
  assign lce_req_o[49] = 1'b0;
  assign lce_req_o[50] = 1'b0;
  assign lce_req_o[51] = 1'b0;
  assign lce_req_o[52] = 1'b0;
  assign lce_req_o[53] = 1'b0;
  assign lce_req_o[54] = 1'b0;
  assign lce_req_o[55] = 1'b0;
  assign lce_req_o[56] = 1'b0;
  assign lce_req_o[57] = 1'b0;
  assign lce_req_o[58] = 1'b0;
  assign lce_req_o[59] = 1'b0;
  assign lce_req_o[60] = 1'b0;
  assign lce_req_o[61] = 1'b0;
  assign lce_req_o[62] = 1'b0;
  assign lce_req_o[63] = 1'b0;
  assign lce_req_o[64] = 1'b0;
  assign lce_req_o[65] = 1'b0;
  assign lce_req_o[66] = 1'b0;
  assign lce_req_o[67] = 1'b0;
  assign lce_req_o[68] = 1'b0;
  assign lce_req_o[69] = 1'b0;
  assign lce_req_o[70] = 1'b0;
  assign lce_req_o[71] = 1'b0;
  assign lce_req_o[72] = 1'b0;
  assign lce_req_o[73] = 1'b0;
  assign lce_req_o[74] = 1'b0;
  assign lce_req_o[75] = 1'b0;
  assign lce_req_o[76] = 1'b0;
  assign lce_req_o[77] = 1'b0;
  assign lce_req_o[78] = 1'b0;
  assign lce_req_o[79] = 1'b0;
  assign lce_req_o[80] = 1'b0;
  assign lce_req_o[81] = 1'b0;
  assign lce_req_o[82] = 1'b0;
  assign lce_req_o[83] = 1'b0;
  assign lce_req_o[84] = 1'b0;
  assign lce_req_o[85] = 1'b0;
  assign lce_req_o[86] = 1'b0;
  assign lce_req_o[87] = 1'b0;
  assign lce_req_o[88] = 1'b0;
  assign lce_req_o[89] = 1'b0;
  assign lce_req_o[90] = 1'b0;
  assign lce_req_o[91] = 1'b0;
  assign lce_req_o[92] = 1'b0;
  assign lce_req_o[93] = 1'b0;
  assign lce_req_o[94] = 1'b0;
  assign lce_req_o[95] = 1'b0;
  assign lce_req_o[96] = 1'b0;
  assign lce_resp_o[21] = miss_addr_o[21];
  assign lce_req_o[28] = miss_addr_o[21];
  assign lce_resp_o[20] = miss_addr_o[20];
  assign lce_req_o[27] = miss_addr_o[20];
  assign lce_resp_o[19] = miss_addr_o[19];
  assign lce_req_o[26] = miss_addr_o[19];
  assign lce_resp_o[18] = miss_addr_o[18];
  assign lce_req_o[25] = miss_addr_o[18];
  assign lce_resp_o[17] = miss_addr_o[17];
  assign lce_req_o[24] = miss_addr_o[17];
  assign lce_resp_o[16] = miss_addr_o[16];
  assign lce_req_o[23] = miss_addr_o[16];
  assign lce_resp_o[15] = miss_addr_o[15];
  assign lce_req_o[22] = miss_addr_o[15];
  assign lce_resp_o[14] = miss_addr_o[14];
  assign lce_req_o[21] = miss_addr_o[14];
  assign lce_resp_o[13] = miss_addr_o[13];
  assign lce_req_o[20] = miss_addr_o[13];
  assign lce_resp_o[12] = miss_addr_o[12];
  assign lce_req_o[19] = miss_addr_o[12];
  assign lce_resp_o[11] = miss_addr_o[11];
  assign lce_req_o[18] = miss_addr_o[11];
  assign lce_resp_o[10] = miss_addr_o[10];
  assign lce_req_o[17] = miss_addr_o[10];
  assign lce_resp_o[9] = miss_addr_o[9];
  assign lce_req_o[16] = miss_addr_o[9];
  assign lce_resp_o[8] = miss_addr_o[8];
  assign lce_req_o[15] = miss_addr_o[8];
  assign lce_resp_o[7] = miss_addr_o[7];
  assign lce_req_o[14] = miss_addr_o[7];
  assign lce_resp_o[6] = miss_addr_o[6];
  assign lce_req_o[13] = miss_addr_o[6];
  assign lce_resp_o[5] = miss_addr_o[5];
  assign lce_req_o[12] = miss_addr_o[5];
  assign lce_resp_o[4] = miss_addr_o[4];
  assign lce_req_o[11] = miss_addr_o[4];
  assign lce_resp_o[3] = miss_addr_o[3];
  assign lce_req_o[10] = miss_addr_o[3];
  assign lce_resp_o[2] = miss_addr_o[2];
  assign lce_req_o[9] = miss_addr_o[2];
  assign lce_resp_o[1] = miss_addr_o[1];
  assign lce_req_o[8] = miss_addr_o[1];
  assign lce_resp_o[0] = miss_addr_o[0];
  assign lce_req_o[7] = miss_addr_o[0];
  assign lce_resp_o[24] = id_i[0];
  assign lce_req_o[31] = id_i[0];
  assign lce_req_o[32] = lce_resp_o[25];
  assign N16 = N13 & N14;
  assign N17 = N16 & N15;
  assign N18 = state_r[2] | state_r[1];
  assign N19 = N18 | N15;
  assign N21 = N13 | state_r[1];
  assign N22 = N21 | state_r[0];
  assign N24 = state_r[2] | N14;
  assign N25 = N24 | state_r[0];
  assign N27 = state_r[2] | N14;
  assign N28 = N27 | N15;
  assign N30 = state_r[2] & state_r[0];
  assign N31 = state_r[2] & state_r[1];
  assign lce_req_o[6:4] = (N0)? lru_way_r :
                          (N1)? lru_way_i : 1'b0;
  assign N0 = lru_flopped_r;
  assign N1 = N12;
  assign { N44, N43, N42 } = (N2)? { 1'b0, 1'b1, 1'b0 } :
                             (N52)? { 1'b0, 1'b1, 1'b1 } :
                             (N41)? { 1'b1, 1'b0, 1'b0 } : 1'b0;
  assign N2 = tr_data_received;
  assign { N47, N46, N45 } = (N3)? { 1'b0, 1'b0, 1'b0 } :
                             (N50)? { N44, N43, N42 } :
                             (N39)? { 1'b1, 1'b0, 1'b0 } : 1'b0;
  assign N3 = set_tag_wakeup_received_i;
  assign cache_miss_o = (N4)? miss_i :
                        (N5)? 1'b1 :
                        (N6)? 1'b1 :
                        (N7)? 1'b1 :
                        (N8)? 1'b1 :
                        (N9)? 1'b0 : 1'b0;
  assign N4 = N17;
  assign N5 = N20;
  assign N6 = N23;
  assign N7 = N26;
  assign N8 = N29;
  assign N9 = N32;
  assign state_n = (N4)? { 1'b0, 1'b0, 1'b1 } :
                   (N5)? { lce_req_ready_i, 1'b0, N34 } :
                   (N6)? { N47, N46, N45 } :
                   (N7)? { 1'b0, N48, 1'b0 } :
                   (N8)? { 1'b0, N48, N48 } :
                   (N9)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tr_data_received_n = (N4)? 1'b0 :
                              (N6)? 1'b1 : 1'b0;
  assign cce_data_received_n = (N4)? 1'b0 :
                               (N6)? 1'b1 : 1'b0;
  assign set_tag_received_n = (N4)? 1'b0 :
                              (N6)? 1'b1 : 1'b0;
  assign lce_req_v_o = (N4)? 1'b0 :
                       (N5)? 1'b1 :
                       (N6)? 1'b0 :
                       (N7)? 1'b0 :
                       (N8)? 1'b0 :
                       (N9)? 1'b0 : 1'b0;
  assign lce_resp_v_o = (N4)? 1'b0 :
                        (N5)? 1'b0 :
                        (N6)? 1'b0 :
                        (N7)? 1'b1 :
                        (N8)? 1'b1 :
                        (N9)? 1'b0 : 1'b0;
  assign lce_resp_o[22] = (N4)? 1'b0 :
                          (N5)? 1'b0 :
                          (N6)? 1'b0 :
                          (N7)? 1'b1 :
                          (N8)? 1'b1 :
                          (N9)? 1'b0 : 1'b0;
  assign { N56, N55, N54 } = (N10)? { 1'b0, 1'b0, 1'b0 } :
                             (N11)? state_n : 1'b0;
  assign N10 = reset_i;
  assign N11 = N53;
  assign N57 = (N10)? 1'b0 :
               (N11)? tr_data_received_n : 1'b0;
  assign N58 = (N10)? 1'b0 :
               (N11)? cce_data_received_n : 1'b0;
  assign N59 = (N10)? 1'b0 :
               (N11)? set_tag_received_n : 1'b0;
  assign tr_data_received = tr_data_received_r | tr_data_received_i;
  assign cce_data_received = cce_data_received_r | cce_data_received_i;
  assign set_tag_received = set_tag_received_r | set_tag_received_i;
  assign N12 = ~lru_flopped_r;
  assign N13 = ~state_r[2];
  assign N14 = ~state_r[1];
  assign N15 = ~state_r[0];
  assign N20 = ~N19;
  assign N23 = ~N22;
  assign N26 = ~N25;
  assign N29 = ~N28;
  assign N32 = N30 | N31;
  assign N33 = ~miss_i;
  assign N34 = ~lce_req_ready_i;
  assign N35 = ~tr_data_received_i;
  assign N36 = ~cce_data_received_i;
  assign N37 = ~set_tag_received_i;
  assign N38 = set_tag_received | set_tag_wakeup_received_i;
  assign N39 = ~N38;
  assign N40 = cce_data_received | tr_data_received;
  assign N41 = ~N40;
  assign N48 = ~lce_resp_yumi_i;
  assign N49 = ~set_tag_wakeup_received_i;
  assign N50 = set_tag_received & N49;
  assign N51 = ~tr_data_received;
  assign N52 = cce_data_received & N51;
  assign N53 = ~reset_i;
  assign N60 = N17 & N53;
  assign N61 = N20 & N53;
  assign N62 = lru_flopped_r & N61;
  assign N63 = N60 | N62;
  assign N64 = N23 & N53;
  assign N65 = N63 | N64;
  assign N66 = N26 & N53;
  assign N67 = N65 | N66;
  assign N68 = N29 & N53;
  assign N69 = N67 | N68;
  assign N70 = N32 & N53;
  assign N71 = N69 | N70;
  assign N72 = ~N71;
  assign N73 = N53 & N72;
  assign N74 = N33 & N60;
  assign N75 = ~N74;
  assign N76 = N74 | N61;
  assign N77 = N35 & N64;
  assign N78 = N76 | N77;
  assign N79 = N78 | N66;
  assign N80 = N79 | N68;
  assign N81 = N80 | N70;
  assign N82 = ~N81;
  assign N83 = N36 & N64;
  assign N84 = N76 | N83;
  assign N85 = N84 | N66;
  assign N86 = N85 | N68;
  assign N87 = N86 | N70;
  assign N88 = ~N87;
  assign N89 = N37 & N64;
  assign N90 = N76 | N89;
  assign N91 = N90 | N66;
  assign N92 = N91 | N68;
  assign N93 = N92 | N70;
  assign N94 = ~N93;
  assign N95 = N76 | N64;
  assign N96 = N95 | N66;
  assign N97 = N96 | N68;
  assign N98 = N97 | N70;
  assign N99 = ~N98;
  assign N100 = N53 & N99;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { lce_resp_o[25:25] } <= { 1'b0 };
    end
    if(N73) begin
      { lru_way_r[2:0] } <= { lru_way_i[2:0] };
    end
    if(N75) begin
      { state_r[2:0] } <= { N56, N55, N54 };
    end
    if(reset_i) begin
      lru_flopped_r <= 1'b0;
    end
    if(N82) begin
      tr_data_received_r <= N57;
    end
    if(N88) begin
      cce_data_received_r <= N58;
    end
    if(N94) begin
      set_tag_received_r <= N59;
    end
    if(N100) begin
      { miss_addr_o[21:0] } <= { miss_addr_i[21:0] };
    end
  end


endmodule



module bp_fe_lce_cmd_data_width_p64_paddr_width_p22_lce_data_width_p512_sets_p64_ways_p8_num_cce_p1_num_lce_p2
(
  clk_i,
  reset_i,
  id_i,
  lce_ready_o,
  set_tag_received_o,
  set_tag_wakeup_received_o,
  data_mem_data_i,
  data_mem_pkt_o,
  data_mem_pkt_v_o,
  data_mem_pkt_yumi_i,
  tag_mem_pkt_o,
  tag_mem_pkt_v_o,
  tag_mem_pkt_yumi_i,
  metadata_mem_pkt_v_o,
  metadata_mem_pkt_o,
  metadata_mem_pkt_yumi_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_yumi_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_yumi_o,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i
);

  input [0:0] id_i;
  input [511:0] data_mem_data_i;
  output [521:0] data_mem_pkt_o;
  output [22:0] tag_mem_pkt_o;
  output [9:0] metadata_mem_pkt_o;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  input [35:0] lce_cmd_i;
  output [517:0] lce_data_cmd_o;
  input clk_i;
  input reset_i;
  input data_mem_pkt_yumi_i;
  input tag_mem_pkt_yumi_i;
  input metadata_mem_pkt_yumi_i;
  input lce_resp_yumi_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_ready_i;
  output lce_ready_o;
  output set_tag_received_o;
  output set_tag_wakeup_received_o;
  output data_mem_pkt_v_o;
  output tag_mem_pkt_v_o;
  output metadata_mem_pkt_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_yumi_o;
  output lce_data_cmd_v_o;
  wire [521:0] data_mem_pkt_o;
  wire [22:0] tag_mem_pkt_o;
  wire [9:0] metadata_mem_pkt_o;
  wire [25:0] lce_resp_o;
  wire [536:0] lce_data_resp_o;
  wire [517:0] lce_data_cmd_o;
  wire lce_ready_o,set_tag_received_o,set_tag_wakeup_received_o,data_mem_pkt_v_o,
  tag_mem_pkt_v_o,metadata_mem_pkt_v_o,lce_resp_v_o,lce_data_resp_v_o,lce_cmd_yumi_o,
  lce_data_cmd_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,
  N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,
  N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,
  N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,
  N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,
  N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
  N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,
  N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,
  N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,
  N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,
  N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,
  N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,
  N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
  N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,
  N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,
  N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,
  N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,
  N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,
  N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,
  N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,
  N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,
  N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,
  N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,
  N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,
  N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,
  N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,
  N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,
  N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,
  N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,
  N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,
  N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,
  N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,
  N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,
  N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,
  N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,
  N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,
  N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,
  N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,
  N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,
  N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,
  N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,
  N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,
  N803,N804,N805,N806,N807,N808,N809,N811,N812,N813,N814,N815,N816,N817,N818,N819,
  N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832;
  wire [1:0] state_n;
  reg [511:0] data_r;
  reg [1:0] state_r;
  reg [0:0] syn_ack_cnt_r;
  reg flag_data_buffered_r,flag_invalidate_r;
  assign metadata_mem_pkt_o[0] = 1'b0;
  assign metadata_mem_pkt_o[1] = 1'b0;
  assign metadata_mem_pkt_o[2] = 1'b0;
  assign metadata_mem_pkt_o[3] = 1'b0;
  assign data_mem_pkt_o[0] = 1'b0;
  assign data_mem_pkt_o[1] = 1'b0;
  assign data_mem_pkt_o[2] = 1'b0;
  assign data_mem_pkt_o[3] = 1'b0;
  assign data_mem_pkt_o[4] = 1'b0;
  assign data_mem_pkt_o[5] = 1'b0;
  assign data_mem_pkt_o[6] = 1'b0;
  assign data_mem_pkt_o[7] = 1'b0;
  assign data_mem_pkt_o[8] = 1'b0;
  assign data_mem_pkt_o[9] = 1'b0;
  assign data_mem_pkt_o[10] = 1'b0;
  assign data_mem_pkt_o[11] = 1'b0;
  assign data_mem_pkt_o[12] = 1'b0;
  assign data_mem_pkt_o[13] = 1'b0;
  assign data_mem_pkt_o[14] = 1'b0;
  assign data_mem_pkt_o[15] = 1'b0;
  assign data_mem_pkt_o[16] = 1'b0;
  assign data_mem_pkt_o[17] = 1'b0;
  assign data_mem_pkt_o[18] = 1'b0;
  assign data_mem_pkt_o[19] = 1'b0;
  assign data_mem_pkt_o[20] = 1'b0;
  assign data_mem_pkt_o[21] = 1'b0;
  assign data_mem_pkt_o[22] = 1'b0;
  assign data_mem_pkt_o[23] = 1'b0;
  assign data_mem_pkt_o[24] = 1'b0;
  assign data_mem_pkt_o[25] = 1'b0;
  assign data_mem_pkt_o[26] = 1'b0;
  assign data_mem_pkt_o[27] = 1'b0;
  assign data_mem_pkt_o[28] = 1'b0;
  assign data_mem_pkt_o[29] = 1'b0;
  assign data_mem_pkt_o[30] = 1'b0;
  assign data_mem_pkt_o[31] = 1'b0;
  assign data_mem_pkt_o[32] = 1'b0;
  assign data_mem_pkt_o[33] = 1'b0;
  assign data_mem_pkt_o[34] = 1'b0;
  assign data_mem_pkt_o[35] = 1'b0;
  assign data_mem_pkt_o[36] = 1'b0;
  assign data_mem_pkt_o[37] = 1'b0;
  assign data_mem_pkt_o[38] = 1'b0;
  assign data_mem_pkt_o[39] = 1'b0;
  assign data_mem_pkt_o[40] = 1'b0;
  assign data_mem_pkt_o[41] = 1'b0;
  assign data_mem_pkt_o[42] = 1'b0;
  assign data_mem_pkt_o[43] = 1'b0;
  assign data_mem_pkt_o[44] = 1'b0;
  assign data_mem_pkt_o[45] = 1'b0;
  assign data_mem_pkt_o[46] = 1'b0;
  assign data_mem_pkt_o[47] = 1'b0;
  assign data_mem_pkt_o[48] = 1'b0;
  assign data_mem_pkt_o[49] = 1'b0;
  assign data_mem_pkt_o[50] = 1'b0;
  assign data_mem_pkt_o[51] = 1'b0;
  assign data_mem_pkt_o[52] = 1'b0;
  assign data_mem_pkt_o[53] = 1'b0;
  assign data_mem_pkt_o[54] = 1'b0;
  assign data_mem_pkt_o[55] = 1'b0;
  assign data_mem_pkt_o[56] = 1'b0;
  assign data_mem_pkt_o[57] = 1'b0;
  assign data_mem_pkt_o[58] = 1'b0;
  assign data_mem_pkt_o[59] = 1'b0;
  assign data_mem_pkt_o[60] = 1'b0;
  assign data_mem_pkt_o[61] = 1'b0;
  assign data_mem_pkt_o[62] = 1'b0;
  assign data_mem_pkt_o[63] = 1'b0;
  assign data_mem_pkt_o[64] = 1'b0;
  assign data_mem_pkt_o[65] = 1'b0;
  assign data_mem_pkt_o[66] = 1'b0;
  assign data_mem_pkt_o[67] = 1'b0;
  assign data_mem_pkt_o[68] = 1'b0;
  assign data_mem_pkt_o[69] = 1'b0;
  assign data_mem_pkt_o[70] = 1'b0;
  assign data_mem_pkt_o[71] = 1'b0;
  assign data_mem_pkt_o[72] = 1'b0;
  assign data_mem_pkt_o[73] = 1'b0;
  assign data_mem_pkt_o[74] = 1'b0;
  assign data_mem_pkt_o[75] = 1'b0;
  assign data_mem_pkt_o[76] = 1'b0;
  assign data_mem_pkt_o[77] = 1'b0;
  assign data_mem_pkt_o[78] = 1'b0;
  assign data_mem_pkt_o[79] = 1'b0;
  assign data_mem_pkt_o[80] = 1'b0;
  assign data_mem_pkt_o[81] = 1'b0;
  assign data_mem_pkt_o[82] = 1'b0;
  assign data_mem_pkt_o[83] = 1'b0;
  assign data_mem_pkt_o[84] = 1'b0;
  assign data_mem_pkt_o[85] = 1'b0;
  assign data_mem_pkt_o[86] = 1'b0;
  assign data_mem_pkt_o[87] = 1'b0;
  assign data_mem_pkt_o[88] = 1'b0;
  assign data_mem_pkt_o[89] = 1'b0;
  assign data_mem_pkt_o[90] = 1'b0;
  assign data_mem_pkt_o[91] = 1'b0;
  assign data_mem_pkt_o[92] = 1'b0;
  assign data_mem_pkt_o[93] = 1'b0;
  assign data_mem_pkt_o[94] = 1'b0;
  assign data_mem_pkt_o[95] = 1'b0;
  assign data_mem_pkt_o[96] = 1'b0;
  assign data_mem_pkt_o[97] = 1'b0;
  assign data_mem_pkt_o[98] = 1'b0;
  assign data_mem_pkt_o[99] = 1'b0;
  assign data_mem_pkt_o[100] = 1'b0;
  assign data_mem_pkt_o[101] = 1'b0;
  assign data_mem_pkt_o[102] = 1'b0;
  assign data_mem_pkt_o[103] = 1'b0;
  assign data_mem_pkt_o[104] = 1'b0;
  assign data_mem_pkt_o[105] = 1'b0;
  assign data_mem_pkt_o[106] = 1'b0;
  assign data_mem_pkt_o[107] = 1'b0;
  assign data_mem_pkt_o[108] = 1'b0;
  assign data_mem_pkt_o[109] = 1'b0;
  assign data_mem_pkt_o[110] = 1'b0;
  assign data_mem_pkt_o[111] = 1'b0;
  assign data_mem_pkt_o[112] = 1'b0;
  assign data_mem_pkt_o[113] = 1'b0;
  assign data_mem_pkt_o[114] = 1'b0;
  assign data_mem_pkt_o[115] = 1'b0;
  assign data_mem_pkt_o[116] = 1'b0;
  assign data_mem_pkt_o[117] = 1'b0;
  assign data_mem_pkt_o[118] = 1'b0;
  assign data_mem_pkt_o[119] = 1'b0;
  assign data_mem_pkt_o[120] = 1'b0;
  assign data_mem_pkt_o[121] = 1'b0;
  assign data_mem_pkt_o[122] = 1'b0;
  assign data_mem_pkt_o[123] = 1'b0;
  assign data_mem_pkt_o[124] = 1'b0;
  assign data_mem_pkt_o[125] = 1'b0;
  assign data_mem_pkt_o[126] = 1'b0;
  assign data_mem_pkt_o[127] = 1'b0;
  assign data_mem_pkt_o[128] = 1'b0;
  assign data_mem_pkt_o[129] = 1'b0;
  assign data_mem_pkt_o[130] = 1'b0;
  assign data_mem_pkt_o[131] = 1'b0;
  assign data_mem_pkt_o[132] = 1'b0;
  assign data_mem_pkt_o[133] = 1'b0;
  assign data_mem_pkt_o[134] = 1'b0;
  assign data_mem_pkt_o[135] = 1'b0;
  assign data_mem_pkt_o[136] = 1'b0;
  assign data_mem_pkt_o[137] = 1'b0;
  assign data_mem_pkt_o[138] = 1'b0;
  assign data_mem_pkt_o[139] = 1'b0;
  assign data_mem_pkt_o[140] = 1'b0;
  assign data_mem_pkt_o[141] = 1'b0;
  assign data_mem_pkt_o[142] = 1'b0;
  assign data_mem_pkt_o[143] = 1'b0;
  assign data_mem_pkt_o[144] = 1'b0;
  assign data_mem_pkt_o[145] = 1'b0;
  assign data_mem_pkt_o[146] = 1'b0;
  assign data_mem_pkt_o[147] = 1'b0;
  assign data_mem_pkt_o[148] = 1'b0;
  assign data_mem_pkt_o[149] = 1'b0;
  assign data_mem_pkt_o[150] = 1'b0;
  assign data_mem_pkt_o[151] = 1'b0;
  assign data_mem_pkt_o[152] = 1'b0;
  assign data_mem_pkt_o[153] = 1'b0;
  assign data_mem_pkt_o[154] = 1'b0;
  assign data_mem_pkt_o[155] = 1'b0;
  assign data_mem_pkt_o[156] = 1'b0;
  assign data_mem_pkt_o[157] = 1'b0;
  assign data_mem_pkt_o[158] = 1'b0;
  assign data_mem_pkt_o[159] = 1'b0;
  assign data_mem_pkt_o[160] = 1'b0;
  assign data_mem_pkt_o[161] = 1'b0;
  assign data_mem_pkt_o[162] = 1'b0;
  assign data_mem_pkt_o[163] = 1'b0;
  assign data_mem_pkt_o[164] = 1'b0;
  assign data_mem_pkt_o[165] = 1'b0;
  assign data_mem_pkt_o[166] = 1'b0;
  assign data_mem_pkt_o[167] = 1'b0;
  assign data_mem_pkt_o[168] = 1'b0;
  assign data_mem_pkt_o[169] = 1'b0;
  assign data_mem_pkt_o[170] = 1'b0;
  assign data_mem_pkt_o[171] = 1'b0;
  assign data_mem_pkt_o[172] = 1'b0;
  assign data_mem_pkt_o[173] = 1'b0;
  assign data_mem_pkt_o[174] = 1'b0;
  assign data_mem_pkt_o[175] = 1'b0;
  assign data_mem_pkt_o[176] = 1'b0;
  assign data_mem_pkt_o[177] = 1'b0;
  assign data_mem_pkt_o[178] = 1'b0;
  assign data_mem_pkt_o[179] = 1'b0;
  assign data_mem_pkt_o[180] = 1'b0;
  assign data_mem_pkt_o[181] = 1'b0;
  assign data_mem_pkt_o[182] = 1'b0;
  assign data_mem_pkt_o[183] = 1'b0;
  assign data_mem_pkt_o[184] = 1'b0;
  assign data_mem_pkt_o[185] = 1'b0;
  assign data_mem_pkt_o[186] = 1'b0;
  assign data_mem_pkt_o[187] = 1'b0;
  assign data_mem_pkt_o[188] = 1'b0;
  assign data_mem_pkt_o[189] = 1'b0;
  assign data_mem_pkt_o[190] = 1'b0;
  assign data_mem_pkt_o[191] = 1'b0;
  assign data_mem_pkt_o[192] = 1'b0;
  assign data_mem_pkt_o[193] = 1'b0;
  assign data_mem_pkt_o[194] = 1'b0;
  assign data_mem_pkt_o[195] = 1'b0;
  assign data_mem_pkt_o[196] = 1'b0;
  assign data_mem_pkt_o[197] = 1'b0;
  assign data_mem_pkt_o[198] = 1'b0;
  assign data_mem_pkt_o[199] = 1'b0;
  assign data_mem_pkt_o[200] = 1'b0;
  assign data_mem_pkt_o[201] = 1'b0;
  assign data_mem_pkt_o[202] = 1'b0;
  assign data_mem_pkt_o[203] = 1'b0;
  assign data_mem_pkt_o[204] = 1'b0;
  assign data_mem_pkt_o[205] = 1'b0;
  assign data_mem_pkt_o[206] = 1'b0;
  assign data_mem_pkt_o[207] = 1'b0;
  assign data_mem_pkt_o[208] = 1'b0;
  assign data_mem_pkt_o[209] = 1'b0;
  assign data_mem_pkt_o[210] = 1'b0;
  assign data_mem_pkt_o[211] = 1'b0;
  assign data_mem_pkt_o[212] = 1'b0;
  assign data_mem_pkt_o[213] = 1'b0;
  assign data_mem_pkt_o[214] = 1'b0;
  assign data_mem_pkt_o[215] = 1'b0;
  assign data_mem_pkt_o[216] = 1'b0;
  assign data_mem_pkt_o[217] = 1'b0;
  assign data_mem_pkt_o[218] = 1'b0;
  assign data_mem_pkt_o[219] = 1'b0;
  assign data_mem_pkt_o[220] = 1'b0;
  assign data_mem_pkt_o[221] = 1'b0;
  assign data_mem_pkt_o[222] = 1'b0;
  assign data_mem_pkt_o[223] = 1'b0;
  assign data_mem_pkt_o[224] = 1'b0;
  assign data_mem_pkt_o[225] = 1'b0;
  assign data_mem_pkt_o[226] = 1'b0;
  assign data_mem_pkt_o[227] = 1'b0;
  assign data_mem_pkt_o[228] = 1'b0;
  assign data_mem_pkt_o[229] = 1'b0;
  assign data_mem_pkt_o[230] = 1'b0;
  assign data_mem_pkt_o[231] = 1'b0;
  assign data_mem_pkt_o[232] = 1'b0;
  assign data_mem_pkt_o[233] = 1'b0;
  assign data_mem_pkt_o[234] = 1'b0;
  assign data_mem_pkt_o[235] = 1'b0;
  assign data_mem_pkt_o[236] = 1'b0;
  assign data_mem_pkt_o[237] = 1'b0;
  assign data_mem_pkt_o[238] = 1'b0;
  assign data_mem_pkt_o[239] = 1'b0;
  assign data_mem_pkt_o[240] = 1'b0;
  assign data_mem_pkt_o[241] = 1'b0;
  assign data_mem_pkt_o[242] = 1'b0;
  assign data_mem_pkt_o[243] = 1'b0;
  assign data_mem_pkt_o[244] = 1'b0;
  assign data_mem_pkt_o[245] = 1'b0;
  assign data_mem_pkt_o[246] = 1'b0;
  assign data_mem_pkt_o[247] = 1'b0;
  assign data_mem_pkt_o[248] = 1'b0;
  assign data_mem_pkt_o[249] = 1'b0;
  assign data_mem_pkt_o[250] = 1'b0;
  assign data_mem_pkt_o[251] = 1'b0;
  assign data_mem_pkt_o[252] = 1'b0;
  assign data_mem_pkt_o[253] = 1'b0;
  assign data_mem_pkt_o[254] = 1'b0;
  assign data_mem_pkt_o[255] = 1'b0;
  assign data_mem_pkt_o[256] = 1'b0;
  assign data_mem_pkt_o[257] = 1'b0;
  assign data_mem_pkt_o[258] = 1'b0;
  assign data_mem_pkt_o[259] = 1'b0;
  assign data_mem_pkt_o[260] = 1'b0;
  assign data_mem_pkt_o[261] = 1'b0;
  assign data_mem_pkt_o[262] = 1'b0;
  assign data_mem_pkt_o[263] = 1'b0;
  assign data_mem_pkt_o[264] = 1'b0;
  assign data_mem_pkt_o[265] = 1'b0;
  assign data_mem_pkt_o[266] = 1'b0;
  assign data_mem_pkt_o[267] = 1'b0;
  assign data_mem_pkt_o[268] = 1'b0;
  assign data_mem_pkt_o[269] = 1'b0;
  assign data_mem_pkt_o[270] = 1'b0;
  assign data_mem_pkt_o[271] = 1'b0;
  assign data_mem_pkt_o[272] = 1'b0;
  assign data_mem_pkt_o[273] = 1'b0;
  assign data_mem_pkt_o[274] = 1'b0;
  assign data_mem_pkt_o[275] = 1'b0;
  assign data_mem_pkt_o[276] = 1'b0;
  assign data_mem_pkt_o[277] = 1'b0;
  assign data_mem_pkt_o[278] = 1'b0;
  assign data_mem_pkt_o[279] = 1'b0;
  assign data_mem_pkt_o[280] = 1'b0;
  assign data_mem_pkt_o[281] = 1'b0;
  assign data_mem_pkt_o[282] = 1'b0;
  assign data_mem_pkt_o[283] = 1'b0;
  assign data_mem_pkt_o[284] = 1'b0;
  assign data_mem_pkt_o[285] = 1'b0;
  assign data_mem_pkt_o[286] = 1'b0;
  assign data_mem_pkt_o[287] = 1'b0;
  assign data_mem_pkt_o[288] = 1'b0;
  assign data_mem_pkt_o[289] = 1'b0;
  assign data_mem_pkt_o[290] = 1'b0;
  assign data_mem_pkt_o[291] = 1'b0;
  assign data_mem_pkt_o[292] = 1'b0;
  assign data_mem_pkt_o[293] = 1'b0;
  assign data_mem_pkt_o[294] = 1'b0;
  assign data_mem_pkt_o[295] = 1'b0;
  assign data_mem_pkt_o[296] = 1'b0;
  assign data_mem_pkt_o[297] = 1'b0;
  assign data_mem_pkt_o[298] = 1'b0;
  assign data_mem_pkt_o[299] = 1'b0;
  assign data_mem_pkt_o[300] = 1'b0;
  assign data_mem_pkt_o[301] = 1'b0;
  assign data_mem_pkt_o[302] = 1'b0;
  assign data_mem_pkt_o[303] = 1'b0;
  assign data_mem_pkt_o[304] = 1'b0;
  assign data_mem_pkt_o[305] = 1'b0;
  assign data_mem_pkt_o[306] = 1'b0;
  assign data_mem_pkt_o[307] = 1'b0;
  assign data_mem_pkt_o[308] = 1'b0;
  assign data_mem_pkt_o[309] = 1'b0;
  assign data_mem_pkt_o[310] = 1'b0;
  assign data_mem_pkt_o[311] = 1'b0;
  assign data_mem_pkt_o[312] = 1'b0;
  assign data_mem_pkt_o[313] = 1'b0;
  assign data_mem_pkt_o[314] = 1'b0;
  assign data_mem_pkt_o[315] = 1'b0;
  assign data_mem_pkt_o[316] = 1'b0;
  assign data_mem_pkt_o[317] = 1'b0;
  assign data_mem_pkt_o[318] = 1'b0;
  assign data_mem_pkt_o[319] = 1'b0;
  assign data_mem_pkt_o[320] = 1'b0;
  assign data_mem_pkt_o[321] = 1'b0;
  assign data_mem_pkt_o[322] = 1'b0;
  assign data_mem_pkt_o[323] = 1'b0;
  assign data_mem_pkt_o[324] = 1'b0;
  assign data_mem_pkt_o[325] = 1'b0;
  assign data_mem_pkt_o[326] = 1'b0;
  assign data_mem_pkt_o[327] = 1'b0;
  assign data_mem_pkt_o[328] = 1'b0;
  assign data_mem_pkt_o[329] = 1'b0;
  assign data_mem_pkt_o[330] = 1'b0;
  assign data_mem_pkt_o[331] = 1'b0;
  assign data_mem_pkt_o[332] = 1'b0;
  assign data_mem_pkt_o[333] = 1'b0;
  assign data_mem_pkt_o[334] = 1'b0;
  assign data_mem_pkt_o[335] = 1'b0;
  assign data_mem_pkt_o[336] = 1'b0;
  assign data_mem_pkt_o[337] = 1'b0;
  assign data_mem_pkt_o[338] = 1'b0;
  assign data_mem_pkt_o[339] = 1'b0;
  assign data_mem_pkt_o[340] = 1'b0;
  assign data_mem_pkt_o[341] = 1'b0;
  assign data_mem_pkt_o[342] = 1'b0;
  assign data_mem_pkt_o[343] = 1'b0;
  assign data_mem_pkt_o[344] = 1'b0;
  assign data_mem_pkt_o[345] = 1'b0;
  assign data_mem_pkt_o[346] = 1'b0;
  assign data_mem_pkt_o[347] = 1'b0;
  assign data_mem_pkt_o[348] = 1'b0;
  assign data_mem_pkt_o[349] = 1'b0;
  assign data_mem_pkt_o[350] = 1'b0;
  assign data_mem_pkt_o[351] = 1'b0;
  assign data_mem_pkt_o[352] = 1'b0;
  assign data_mem_pkt_o[353] = 1'b0;
  assign data_mem_pkt_o[354] = 1'b0;
  assign data_mem_pkt_o[355] = 1'b0;
  assign data_mem_pkt_o[356] = 1'b0;
  assign data_mem_pkt_o[357] = 1'b0;
  assign data_mem_pkt_o[358] = 1'b0;
  assign data_mem_pkt_o[359] = 1'b0;
  assign data_mem_pkt_o[360] = 1'b0;
  assign data_mem_pkt_o[361] = 1'b0;
  assign data_mem_pkt_o[362] = 1'b0;
  assign data_mem_pkt_o[363] = 1'b0;
  assign data_mem_pkt_o[364] = 1'b0;
  assign data_mem_pkt_o[365] = 1'b0;
  assign data_mem_pkt_o[366] = 1'b0;
  assign data_mem_pkt_o[367] = 1'b0;
  assign data_mem_pkt_o[368] = 1'b0;
  assign data_mem_pkt_o[369] = 1'b0;
  assign data_mem_pkt_o[370] = 1'b0;
  assign data_mem_pkt_o[371] = 1'b0;
  assign data_mem_pkt_o[372] = 1'b0;
  assign data_mem_pkt_o[373] = 1'b0;
  assign data_mem_pkt_o[374] = 1'b0;
  assign data_mem_pkt_o[375] = 1'b0;
  assign data_mem_pkt_o[376] = 1'b0;
  assign data_mem_pkt_o[377] = 1'b0;
  assign data_mem_pkt_o[378] = 1'b0;
  assign data_mem_pkt_o[379] = 1'b0;
  assign data_mem_pkt_o[380] = 1'b0;
  assign data_mem_pkt_o[381] = 1'b0;
  assign data_mem_pkt_o[382] = 1'b0;
  assign data_mem_pkt_o[383] = 1'b0;
  assign data_mem_pkt_o[384] = 1'b0;
  assign data_mem_pkt_o[385] = 1'b0;
  assign data_mem_pkt_o[386] = 1'b0;
  assign data_mem_pkt_o[387] = 1'b0;
  assign data_mem_pkt_o[388] = 1'b0;
  assign data_mem_pkt_o[389] = 1'b0;
  assign data_mem_pkt_o[390] = 1'b0;
  assign data_mem_pkt_o[391] = 1'b0;
  assign data_mem_pkt_o[392] = 1'b0;
  assign data_mem_pkt_o[393] = 1'b0;
  assign data_mem_pkt_o[394] = 1'b0;
  assign data_mem_pkt_o[395] = 1'b0;
  assign data_mem_pkt_o[396] = 1'b0;
  assign data_mem_pkt_o[397] = 1'b0;
  assign data_mem_pkt_o[398] = 1'b0;
  assign data_mem_pkt_o[399] = 1'b0;
  assign data_mem_pkt_o[400] = 1'b0;
  assign data_mem_pkt_o[401] = 1'b0;
  assign data_mem_pkt_o[402] = 1'b0;
  assign data_mem_pkt_o[403] = 1'b0;
  assign data_mem_pkt_o[404] = 1'b0;
  assign data_mem_pkt_o[405] = 1'b0;
  assign data_mem_pkt_o[406] = 1'b0;
  assign data_mem_pkt_o[407] = 1'b0;
  assign data_mem_pkt_o[408] = 1'b0;
  assign data_mem_pkt_o[409] = 1'b0;
  assign data_mem_pkt_o[410] = 1'b0;
  assign data_mem_pkt_o[411] = 1'b0;
  assign data_mem_pkt_o[412] = 1'b0;
  assign data_mem_pkt_o[413] = 1'b0;
  assign data_mem_pkt_o[414] = 1'b0;
  assign data_mem_pkt_o[415] = 1'b0;
  assign data_mem_pkt_o[416] = 1'b0;
  assign data_mem_pkt_o[417] = 1'b0;
  assign data_mem_pkt_o[418] = 1'b0;
  assign data_mem_pkt_o[419] = 1'b0;
  assign data_mem_pkt_o[420] = 1'b0;
  assign data_mem_pkt_o[421] = 1'b0;
  assign data_mem_pkt_o[422] = 1'b0;
  assign data_mem_pkt_o[423] = 1'b0;
  assign data_mem_pkt_o[424] = 1'b0;
  assign data_mem_pkt_o[425] = 1'b0;
  assign data_mem_pkt_o[426] = 1'b0;
  assign data_mem_pkt_o[427] = 1'b0;
  assign data_mem_pkt_o[428] = 1'b0;
  assign data_mem_pkt_o[429] = 1'b0;
  assign data_mem_pkt_o[430] = 1'b0;
  assign data_mem_pkt_o[431] = 1'b0;
  assign data_mem_pkt_o[432] = 1'b0;
  assign data_mem_pkt_o[433] = 1'b0;
  assign data_mem_pkt_o[434] = 1'b0;
  assign data_mem_pkt_o[435] = 1'b0;
  assign data_mem_pkt_o[436] = 1'b0;
  assign data_mem_pkt_o[437] = 1'b0;
  assign data_mem_pkt_o[438] = 1'b0;
  assign data_mem_pkt_o[439] = 1'b0;
  assign data_mem_pkt_o[440] = 1'b0;
  assign data_mem_pkt_o[441] = 1'b0;
  assign data_mem_pkt_o[442] = 1'b0;
  assign data_mem_pkt_o[443] = 1'b0;
  assign data_mem_pkt_o[444] = 1'b0;
  assign data_mem_pkt_o[445] = 1'b0;
  assign data_mem_pkt_o[446] = 1'b0;
  assign data_mem_pkt_o[447] = 1'b0;
  assign data_mem_pkt_o[448] = 1'b0;
  assign data_mem_pkt_o[449] = 1'b0;
  assign data_mem_pkt_o[450] = 1'b0;
  assign data_mem_pkt_o[451] = 1'b0;
  assign data_mem_pkt_o[452] = 1'b0;
  assign data_mem_pkt_o[453] = 1'b0;
  assign data_mem_pkt_o[454] = 1'b0;
  assign data_mem_pkt_o[455] = 1'b0;
  assign data_mem_pkt_o[456] = 1'b0;
  assign data_mem_pkt_o[457] = 1'b0;
  assign data_mem_pkt_o[458] = 1'b0;
  assign data_mem_pkt_o[459] = 1'b0;
  assign data_mem_pkt_o[460] = 1'b0;
  assign data_mem_pkt_o[461] = 1'b0;
  assign data_mem_pkt_o[462] = 1'b0;
  assign data_mem_pkt_o[463] = 1'b0;
  assign data_mem_pkt_o[464] = 1'b0;
  assign data_mem_pkt_o[465] = 1'b0;
  assign data_mem_pkt_o[466] = 1'b0;
  assign data_mem_pkt_o[467] = 1'b0;
  assign data_mem_pkt_o[468] = 1'b0;
  assign data_mem_pkt_o[469] = 1'b0;
  assign data_mem_pkt_o[470] = 1'b0;
  assign data_mem_pkt_o[471] = 1'b0;
  assign data_mem_pkt_o[472] = 1'b0;
  assign data_mem_pkt_o[473] = 1'b0;
  assign data_mem_pkt_o[474] = 1'b0;
  assign data_mem_pkt_o[475] = 1'b0;
  assign data_mem_pkt_o[476] = 1'b0;
  assign data_mem_pkt_o[477] = 1'b0;
  assign data_mem_pkt_o[478] = 1'b0;
  assign data_mem_pkt_o[479] = 1'b0;
  assign data_mem_pkt_o[480] = 1'b0;
  assign data_mem_pkt_o[481] = 1'b0;
  assign data_mem_pkt_o[482] = 1'b0;
  assign data_mem_pkt_o[483] = 1'b0;
  assign data_mem_pkt_o[484] = 1'b0;
  assign data_mem_pkt_o[485] = 1'b0;
  assign data_mem_pkt_o[486] = 1'b0;
  assign data_mem_pkt_o[487] = 1'b0;
  assign data_mem_pkt_o[488] = 1'b0;
  assign data_mem_pkt_o[489] = 1'b0;
  assign data_mem_pkt_o[490] = 1'b0;
  assign data_mem_pkt_o[491] = 1'b0;
  assign data_mem_pkt_o[492] = 1'b0;
  assign data_mem_pkt_o[493] = 1'b0;
  assign data_mem_pkt_o[494] = 1'b0;
  assign data_mem_pkt_o[495] = 1'b0;
  assign data_mem_pkt_o[496] = 1'b0;
  assign data_mem_pkt_o[497] = 1'b0;
  assign data_mem_pkt_o[498] = 1'b0;
  assign data_mem_pkt_o[499] = 1'b0;
  assign data_mem_pkt_o[500] = 1'b0;
  assign data_mem_pkt_o[501] = 1'b0;
  assign data_mem_pkt_o[502] = 1'b0;
  assign data_mem_pkt_o[503] = 1'b0;
  assign data_mem_pkt_o[504] = 1'b0;
  assign data_mem_pkt_o[505] = 1'b0;
  assign data_mem_pkt_o[506] = 1'b0;
  assign data_mem_pkt_o[507] = 1'b0;
  assign data_mem_pkt_o[508] = 1'b0;
  assign data_mem_pkt_o[509] = 1'b0;
  assign data_mem_pkt_o[510] = 1'b0;
  assign data_mem_pkt_o[511] = 1'b0;
  assign data_mem_pkt_o[512] = 1'b0;
  assign lce_data_cmd_o[3] = 1'b0;
  assign lce_data_cmd_o[4] = 1'b0;
  assign lce_data_resp_o[25] = 1'b0;
  assign lce_data_resp_o[26] = 1'b0;
  assign lce_data_resp_o[27] = 1'b0;
  assign lce_data_resp_o[28] = 1'b0;
  assign lce_data_resp_o[29] = 1'b0;
  assign lce_data_resp_o[30] = 1'b0;
  assign lce_data_resp_o[31] = 1'b0;
  assign lce_data_resp_o[32] = 1'b0;
  assign lce_data_resp_o[33] = 1'b0;
  assign lce_data_resp_o[34] = 1'b0;
  assign lce_data_resp_o[35] = 1'b0;
  assign lce_data_resp_o[36] = 1'b0;
  assign lce_data_resp_o[37] = 1'b0;
  assign lce_data_resp_o[38] = 1'b0;
  assign lce_data_resp_o[39] = 1'b0;
  assign lce_data_resp_o[40] = 1'b0;
  assign lce_data_resp_o[41] = 1'b0;
  assign lce_data_resp_o[42] = 1'b0;
  assign lce_data_resp_o[43] = 1'b0;
  assign lce_data_resp_o[44] = 1'b0;
  assign lce_data_resp_o[45] = 1'b0;
  assign lce_data_resp_o[46] = 1'b0;
  assign lce_data_resp_o[47] = 1'b0;
  assign lce_data_resp_o[48] = 1'b0;
  assign lce_data_resp_o[49] = 1'b0;
  assign lce_data_resp_o[50] = 1'b0;
  assign lce_data_resp_o[51] = 1'b0;
  assign lce_data_resp_o[52] = 1'b0;
  assign lce_data_resp_o[53] = 1'b0;
  assign lce_data_resp_o[54] = 1'b0;
  assign lce_data_resp_o[55] = 1'b0;
  assign lce_data_resp_o[56] = 1'b0;
  assign lce_data_resp_o[57] = 1'b0;
  assign lce_data_resp_o[58] = 1'b0;
  assign lce_data_resp_o[59] = 1'b0;
  assign lce_data_resp_o[60] = 1'b0;
  assign lce_data_resp_o[61] = 1'b0;
  assign lce_data_resp_o[62] = 1'b0;
  assign lce_data_resp_o[63] = 1'b0;
  assign lce_data_resp_o[64] = 1'b0;
  assign lce_data_resp_o[65] = 1'b0;
  assign lce_data_resp_o[66] = 1'b0;
  assign lce_data_resp_o[67] = 1'b0;
  assign lce_data_resp_o[68] = 1'b0;
  assign lce_data_resp_o[69] = 1'b0;
  assign lce_data_resp_o[70] = 1'b0;
  assign lce_data_resp_o[71] = 1'b0;
  assign lce_data_resp_o[72] = 1'b0;
  assign lce_data_resp_o[73] = 1'b0;
  assign lce_data_resp_o[74] = 1'b0;
  assign lce_data_resp_o[75] = 1'b0;
  assign lce_data_resp_o[76] = 1'b0;
  assign lce_data_resp_o[77] = 1'b0;
  assign lce_data_resp_o[78] = 1'b0;
  assign lce_data_resp_o[79] = 1'b0;
  assign lce_data_resp_o[80] = 1'b0;
  assign lce_data_resp_o[81] = 1'b0;
  assign lce_data_resp_o[82] = 1'b0;
  assign lce_data_resp_o[83] = 1'b0;
  assign lce_data_resp_o[84] = 1'b0;
  assign lce_data_resp_o[85] = 1'b0;
  assign lce_data_resp_o[86] = 1'b0;
  assign lce_data_resp_o[87] = 1'b0;
  assign lce_data_resp_o[88] = 1'b0;
  assign lce_data_resp_o[89] = 1'b0;
  assign lce_data_resp_o[90] = 1'b0;
  assign lce_data_resp_o[91] = 1'b0;
  assign lce_data_resp_o[92] = 1'b0;
  assign lce_data_resp_o[93] = 1'b0;
  assign lce_data_resp_o[94] = 1'b0;
  assign lce_data_resp_o[95] = 1'b0;
  assign lce_data_resp_o[96] = 1'b0;
  assign lce_data_resp_o[97] = 1'b0;
  assign lce_data_resp_o[98] = 1'b0;
  assign lce_data_resp_o[99] = 1'b0;
  assign lce_data_resp_o[100] = 1'b0;
  assign lce_data_resp_o[101] = 1'b0;
  assign lce_data_resp_o[102] = 1'b0;
  assign lce_data_resp_o[103] = 1'b0;
  assign lce_data_resp_o[104] = 1'b0;
  assign lce_data_resp_o[105] = 1'b0;
  assign lce_data_resp_o[106] = 1'b0;
  assign lce_data_resp_o[107] = 1'b0;
  assign lce_data_resp_o[108] = 1'b0;
  assign lce_data_resp_o[109] = 1'b0;
  assign lce_data_resp_o[110] = 1'b0;
  assign lce_data_resp_o[111] = 1'b0;
  assign lce_data_resp_o[112] = 1'b0;
  assign lce_data_resp_o[113] = 1'b0;
  assign lce_data_resp_o[114] = 1'b0;
  assign lce_data_resp_o[115] = 1'b0;
  assign lce_data_resp_o[116] = 1'b0;
  assign lce_data_resp_o[117] = 1'b0;
  assign lce_data_resp_o[118] = 1'b0;
  assign lce_data_resp_o[119] = 1'b0;
  assign lce_data_resp_o[120] = 1'b0;
  assign lce_data_resp_o[121] = 1'b0;
  assign lce_data_resp_o[122] = 1'b0;
  assign lce_data_resp_o[123] = 1'b0;
  assign lce_data_resp_o[124] = 1'b0;
  assign lce_data_resp_o[125] = 1'b0;
  assign lce_data_resp_o[126] = 1'b0;
  assign lce_data_resp_o[127] = 1'b0;
  assign lce_data_resp_o[128] = 1'b0;
  assign lce_data_resp_o[129] = 1'b0;
  assign lce_data_resp_o[130] = 1'b0;
  assign lce_data_resp_o[131] = 1'b0;
  assign lce_data_resp_o[132] = 1'b0;
  assign lce_data_resp_o[133] = 1'b0;
  assign lce_data_resp_o[134] = 1'b0;
  assign lce_data_resp_o[135] = 1'b0;
  assign lce_data_resp_o[136] = 1'b0;
  assign lce_data_resp_o[137] = 1'b0;
  assign lce_data_resp_o[138] = 1'b0;
  assign lce_data_resp_o[139] = 1'b0;
  assign lce_data_resp_o[140] = 1'b0;
  assign lce_data_resp_o[141] = 1'b0;
  assign lce_data_resp_o[142] = 1'b0;
  assign lce_data_resp_o[143] = 1'b0;
  assign lce_data_resp_o[144] = 1'b0;
  assign lce_data_resp_o[145] = 1'b0;
  assign lce_data_resp_o[146] = 1'b0;
  assign lce_data_resp_o[147] = 1'b0;
  assign lce_data_resp_o[148] = 1'b0;
  assign lce_data_resp_o[149] = 1'b0;
  assign lce_data_resp_o[150] = 1'b0;
  assign lce_data_resp_o[151] = 1'b0;
  assign lce_data_resp_o[152] = 1'b0;
  assign lce_data_resp_o[153] = 1'b0;
  assign lce_data_resp_o[154] = 1'b0;
  assign lce_data_resp_o[155] = 1'b0;
  assign lce_data_resp_o[156] = 1'b0;
  assign lce_data_resp_o[157] = 1'b0;
  assign lce_data_resp_o[158] = 1'b0;
  assign lce_data_resp_o[159] = 1'b0;
  assign lce_data_resp_o[160] = 1'b0;
  assign lce_data_resp_o[161] = 1'b0;
  assign lce_data_resp_o[162] = 1'b0;
  assign lce_data_resp_o[163] = 1'b0;
  assign lce_data_resp_o[164] = 1'b0;
  assign lce_data_resp_o[165] = 1'b0;
  assign lce_data_resp_o[166] = 1'b0;
  assign lce_data_resp_o[167] = 1'b0;
  assign lce_data_resp_o[168] = 1'b0;
  assign lce_data_resp_o[169] = 1'b0;
  assign lce_data_resp_o[170] = 1'b0;
  assign lce_data_resp_o[171] = 1'b0;
  assign lce_data_resp_o[172] = 1'b0;
  assign lce_data_resp_o[173] = 1'b0;
  assign lce_data_resp_o[174] = 1'b0;
  assign lce_data_resp_o[175] = 1'b0;
  assign lce_data_resp_o[176] = 1'b0;
  assign lce_data_resp_o[177] = 1'b0;
  assign lce_data_resp_o[178] = 1'b0;
  assign lce_data_resp_o[179] = 1'b0;
  assign lce_data_resp_o[180] = 1'b0;
  assign lce_data_resp_o[181] = 1'b0;
  assign lce_data_resp_o[182] = 1'b0;
  assign lce_data_resp_o[183] = 1'b0;
  assign lce_data_resp_o[184] = 1'b0;
  assign lce_data_resp_o[185] = 1'b0;
  assign lce_data_resp_o[186] = 1'b0;
  assign lce_data_resp_o[187] = 1'b0;
  assign lce_data_resp_o[188] = 1'b0;
  assign lce_data_resp_o[189] = 1'b0;
  assign lce_data_resp_o[190] = 1'b0;
  assign lce_data_resp_o[191] = 1'b0;
  assign lce_data_resp_o[192] = 1'b0;
  assign lce_data_resp_o[193] = 1'b0;
  assign lce_data_resp_o[194] = 1'b0;
  assign lce_data_resp_o[195] = 1'b0;
  assign lce_data_resp_o[196] = 1'b0;
  assign lce_data_resp_o[197] = 1'b0;
  assign lce_data_resp_o[198] = 1'b0;
  assign lce_data_resp_o[199] = 1'b0;
  assign lce_data_resp_o[200] = 1'b0;
  assign lce_data_resp_o[201] = 1'b0;
  assign lce_data_resp_o[202] = 1'b0;
  assign lce_data_resp_o[203] = 1'b0;
  assign lce_data_resp_o[204] = 1'b0;
  assign lce_data_resp_o[205] = 1'b0;
  assign lce_data_resp_o[206] = 1'b0;
  assign lce_data_resp_o[207] = 1'b0;
  assign lce_data_resp_o[208] = 1'b0;
  assign lce_data_resp_o[209] = 1'b0;
  assign lce_data_resp_o[210] = 1'b0;
  assign lce_data_resp_o[211] = 1'b0;
  assign lce_data_resp_o[212] = 1'b0;
  assign lce_data_resp_o[213] = 1'b0;
  assign lce_data_resp_o[214] = 1'b0;
  assign lce_data_resp_o[215] = 1'b0;
  assign lce_data_resp_o[216] = 1'b0;
  assign lce_data_resp_o[217] = 1'b0;
  assign lce_data_resp_o[218] = 1'b0;
  assign lce_data_resp_o[219] = 1'b0;
  assign lce_data_resp_o[220] = 1'b0;
  assign lce_data_resp_o[221] = 1'b0;
  assign lce_data_resp_o[222] = 1'b0;
  assign lce_data_resp_o[223] = 1'b0;
  assign lce_data_resp_o[224] = 1'b0;
  assign lce_data_resp_o[225] = 1'b0;
  assign lce_data_resp_o[226] = 1'b0;
  assign lce_data_resp_o[227] = 1'b0;
  assign lce_data_resp_o[228] = 1'b0;
  assign lce_data_resp_o[229] = 1'b0;
  assign lce_data_resp_o[230] = 1'b0;
  assign lce_data_resp_o[231] = 1'b0;
  assign lce_data_resp_o[232] = 1'b0;
  assign lce_data_resp_o[233] = 1'b0;
  assign lce_data_resp_o[234] = 1'b0;
  assign lce_data_resp_o[235] = 1'b0;
  assign lce_data_resp_o[236] = 1'b0;
  assign lce_data_resp_o[237] = 1'b0;
  assign lce_data_resp_o[238] = 1'b0;
  assign lce_data_resp_o[239] = 1'b0;
  assign lce_data_resp_o[240] = 1'b0;
  assign lce_data_resp_o[241] = 1'b0;
  assign lce_data_resp_o[242] = 1'b0;
  assign lce_data_resp_o[243] = 1'b0;
  assign lce_data_resp_o[244] = 1'b0;
  assign lce_data_resp_o[245] = 1'b0;
  assign lce_data_resp_o[246] = 1'b0;
  assign lce_data_resp_o[247] = 1'b0;
  assign lce_data_resp_o[248] = 1'b0;
  assign lce_data_resp_o[249] = 1'b0;
  assign lce_data_resp_o[250] = 1'b0;
  assign lce_data_resp_o[251] = 1'b0;
  assign lce_data_resp_o[252] = 1'b0;
  assign lce_data_resp_o[253] = 1'b0;
  assign lce_data_resp_o[254] = 1'b0;
  assign lce_data_resp_o[255] = 1'b0;
  assign lce_data_resp_o[256] = 1'b0;
  assign lce_data_resp_o[257] = 1'b0;
  assign lce_data_resp_o[258] = 1'b0;
  assign lce_data_resp_o[259] = 1'b0;
  assign lce_data_resp_o[260] = 1'b0;
  assign lce_data_resp_o[261] = 1'b0;
  assign lce_data_resp_o[262] = 1'b0;
  assign lce_data_resp_o[263] = 1'b0;
  assign lce_data_resp_o[264] = 1'b0;
  assign lce_data_resp_o[265] = 1'b0;
  assign lce_data_resp_o[266] = 1'b0;
  assign lce_data_resp_o[267] = 1'b0;
  assign lce_data_resp_o[268] = 1'b0;
  assign lce_data_resp_o[269] = 1'b0;
  assign lce_data_resp_o[270] = 1'b0;
  assign lce_data_resp_o[271] = 1'b0;
  assign lce_data_resp_o[272] = 1'b0;
  assign lce_data_resp_o[273] = 1'b0;
  assign lce_data_resp_o[274] = 1'b0;
  assign lce_data_resp_o[275] = 1'b0;
  assign lce_data_resp_o[276] = 1'b0;
  assign lce_data_resp_o[277] = 1'b0;
  assign lce_data_resp_o[278] = 1'b0;
  assign lce_data_resp_o[279] = 1'b0;
  assign lce_data_resp_o[280] = 1'b0;
  assign lce_data_resp_o[281] = 1'b0;
  assign lce_data_resp_o[282] = 1'b0;
  assign lce_data_resp_o[283] = 1'b0;
  assign lce_data_resp_o[284] = 1'b0;
  assign lce_data_resp_o[285] = 1'b0;
  assign lce_data_resp_o[286] = 1'b0;
  assign lce_data_resp_o[287] = 1'b0;
  assign lce_data_resp_o[288] = 1'b0;
  assign lce_data_resp_o[289] = 1'b0;
  assign lce_data_resp_o[290] = 1'b0;
  assign lce_data_resp_o[291] = 1'b0;
  assign lce_data_resp_o[292] = 1'b0;
  assign lce_data_resp_o[293] = 1'b0;
  assign lce_data_resp_o[294] = 1'b0;
  assign lce_data_resp_o[295] = 1'b0;
  assign lce_data_resp_o[296] = 1'b0;
  assign lce_data_resp_o[297] = 1'b0;
  assign lce_data_resp_o[298] = 1'b0;
  assign lce_data_resp_o[299] = 1'b0;
  assign lce_data_resp_o[300] = 1'b0;
  assign lce_data_resp_o[301] = 1'b0;
  assign lce_data_resp_o[302] = 1'b0;
  assign lce_data_resp_o[303] = 1'b0;
  assign lce_data_resp_o[304] = 1'b0;
  assign lce_data_resp_o[305] = 1'b0;
  assign lce_data_resp_o[306] = 1'b0;
  assign lce_data_resp_o[307] = 1'b0;
  assign lce_data_resp_o[308] = 1'b0;
  assign lce_data_resp_o[309] = 1'b0;
  assign lce_data_resp_o[310] = 1'b0;
  assign lce_data_resp_o[311] = 1'b0;
  assign lce_data_resp_o[312] = 1'b0;
  assign lce_data_resp_o[313] = 1'b0;
  assign lce_data_resp_o[314] = 1'b0;
  assign lce_data_resp_o[315] = 1'b0;
  assign lce_data_resp_o[316] = 1'b0;
  assign lce_data_resp_o[317] = 1'b0;
  assign lce_data_resp_o[318] = 1'b0;
  assign lce_data_resp_o[319] = 1'b0;
  assign lce_data_resp_o[320] = 1'b0;
  assign lce_data_resp_o[321] = 1'b0;
  assign lce_data_resp_o[322] = 1'b0;
  assign lce_data_resp_o[323] = 1'b0;
  assign lce_data_resp_o[324] = 1'b0;
  assign lce_data_resp_o[325] = 1'b0;
  assign lce_data_resp_o[326] = 1'b0;
  assign lce_data_resp_o[327] = 1'b0;
  assign lce_data_resp_o[328] = 1'b0;
  assign lce_data_resp_o[329] = 1'b0;
  assign lce_data_resp_o[330] = 1'b0;
  assign lce_data_resp_o[331] = 1'b0;
  assign lce_data_resp_o[332] = 1'b0;
  assign lce_data_resp_o[333] = 1'b0;
  assign lce_data_resp_o[334] = 1'b0;
  assign lce_data_resp_o[335] = 1'b0;
  assign lce_data_resp_o[336] = 1'b0;
  assign lce_data_resp_o[337] = 1'b0;
  assign lce_data_resp_o[338] = 1'b0;
  assign lce_data_resp_o[339] = 1'b0;
  assign lce_data_resp_o[340] = 1'b0;
  assign lce_data_resp_o[341] = 1'b0;
  assign lce_data_resp_o[342] = 1'b0;
  assign lce_data_resp_o[343] = 1'b0;
  assign lce_data_resp_o[344] = 1'b0;
  assign lce_data_resp_o[345] = 1'b0;
  assign lce_data_resp_o[346] = 1'b0;
  assign lce_data_resp_o[347] = 1'b0;
  assign lce_data_resp_o[348] = 1'b0;
  assign lce_data_resp_o[349] = 1'b0;
  assign lce_data_resp_o[350] = 1'b0;
  assign lce_data_resp_o[351] = 1'b0;
  assign lce_data_resp_o[352] = 1'b0;
  assign lce_data_resp_o[353] = 1'b0;
  assign lce_data_resp_o[354] = 1'b0;
  assign lce_data_resp_o[355] = 1'b0;
  assign lce_data_resp_o[356] = 1'b0;
  assign lce_data_resp_o[357] = 1'b0;
  assign lce_data_resp_o[358] = 1'b0;
  assign lce_data_resp_o[359] = 1'b0;
  assign lce_data_resp_o[360] = 1'b0;
  assign lce_data_resp_o[361] = 1'b0;
  assign lce_data_resp_o[362] = 1'b0;
  assign lce_data_resp_o[363] = 1'b0;
  assign lce_data_resp_o[364] = 1'b0;
  assign lce_data_resp_o[365] = 1'b0;
  assign lce_data_resp_o[366] = 1'b0;
  assign lce_data_resp_o[367] = 1'b0;
  assign lce_data_resp_o[368] = 1'b0;
  assign lce_data_resp_o[369] = 1'b0;
  assign lce_data_resp_o[370] = 1'b0;
  assign lce_data_resp_o[371] = 1'b0;
  assign lce_data_resp_o[372] = 1'b0;
  assign lce_data_resp_o[373] = 1'b0;
  assign lce_data_resp_o[374] = 1'b0;
  assign lce_data_resp_o[375] = 1'b0;
  assign lce_data_resp_o[376] = 1'b0;
  assign lce_data_resp_o[377] = 1'b0;
  assign lce_data_resp_o[378] = 1'b0;
  assign lce_data_resp_o[379] = 1'b0;
  assign lce_data_resp_o[380] = 1'b0;
  assign lce_data_resp_o[381] = 1'b0;
  assign lce_data_resp_o[382] = 1'b0;
  assign lce_data_resp_o[383] = 1'b0;
  assign lce_data_resp_o[384] = 1'b0;
  assign lce_data_resp_o[385] = 1'b0;
  assign lce_data_resp_o[386] = 1'b0;
  assign lce_data_resp_o[387] = 1'b0;
  assign lce_data_resp_o[388] = 1'b0;
  assign lce_data_resp_o[389] = 1'b0;
  assign lce_data_resp_o[390] = 1'b0;
  assign lce_data_resp_o[391] = 1'b0;
  assign lce_data_resp_o[392] = 1'b0;
  assign lce_data_resp_o[393] = 1'b0;
  assign lce_data_resp_o[394] = 1'b0;
  assign lce_data_resp_o[395] = 1'b0;
  assign lce_data_resp_o[396] = 1'b0;
  assign lce_data_resp_o[397] = 1'b0;
  assign lce_data_resp_o[398] = 1'b0;
  assign lce_data_resp_o[399] = 1'b0;
  assign lce_data_resp_o[400] = 1'b0;
  assign lce_data_resp_o[401] = 1'b0;
  assign lce_data_resp_o[402] = 1'b0;
  assign lce_data_resp_o[403] = 1'b0;
  assign lce_data_resp_o[404] = 1'b0;
  assign lce_data_resp_o[405] = 1'b0;
  assign lce_data_resp_o[406] = 1'b0;
  assign lce_data_resp_o[407] = 1'b0;
  assign lce_data_resp_o[408] = 1'b0;
  assign lce_data_resp_o[409] = 1'b0;
  assign lce_data_resp_o[410] = 1'b0;
  assign lce_data_resp_o[411] = 1'b0;
  assign lce_data_resp_o[412] = 1'b0;
  assign lce_data_resp_o[413] = 1'b0;
  assign lce_data_resp_o[414] = 1'b0;
  assign lce_data_resp_o[415] = 1'b0;
  assign lce_data_resp_o[416] = 1'b0;
  assign lce_data_resp_o[417] = 1'b0;
  assign lce_data_resp_o[418] = 1'b0;
  assign lce_data_resp_o[419] = 1'b0;
  assign lce_data_resp_o[420] = 1'b0;
  assign lce_data_resp_o[421] = 1'b0;
  assign lce_data_resp_o[422] = 1'b0;
  assign lce_data_resp_o[423] = 1'b0;
  assign lce_data_resp_o[424] = 1'b0;
  assign lce_data_resp_o[425] = 1'b0;
  assign lce_data_resp_o[426] = 1'b0;
  assign lce_data_resp_o[427] = 1'b0;
  assign lce_data_resp_o[428] = 1'b0;
  assign lce_data_resp_o[429] = 1'b0;
  assign lce_data_resp_o[430] = 1'b0;
  assign lce_data_resp_o[431] = 1'b0;
  assign lce_data_resp_o[432] = 1'b0;
  assign lce_data_resp_o[433] = 1'b0;
  assign lce_data_resp_o[434] = 1'b0;
  assign lce_data_resp_o[435] = 1'b0;
  assign lce_data_resp_o[436] = 1'b0;
  assign lce_data_resp_o[437] = 1'b0;
  assign lce_data_resp_o[438] = 1'b0;
  assign lce_data_resp_o[439] = 1'b0;
  assign lce_data_resp_o[440] = 1'b0;
  assign lce_data_resp_o[441] = 1'b0;
  assign lce_data_resp_o[442] = 1'b0;
  assign lce_data_resp_o[443] = 1'b0;
  assign lce_data_resp_o[444] = 1'b0;
  assign lce_data_resp_o[445] = 1'b0;
  assign lce_data_resp_o[446] = 1'b0;
  assign lce_data_resp_o[447] = 1'b0;
  assign lce_data_resp_o[448] = 1'b0;
  assign lce_data_resp_o[449] = 1'b0;
  assign lce_data_resp_o[450] = 1'b0;
  assign lce_data_resp_o[451] = 1'b0;
  assign lce_data_resp_o[452] = 1'b0;
  assign lce_data_resp_o[453] = 1'b0;
  assign lce_data_resp_o[454] = 1'b0;
  assign lce_data_resp_o[455] = 1'b0;
  assign lce_data_resp_o[456] = 1'b0;
  assign lce_data_resp_o[457] = 1'b0;
  assign lce_data_resp_o[458] = 1'b0;
  assign lce_data_resp_o[459] = 1'b0;
  assign lce_data_resp_o[460] = 1'b0;
  assign lce_data_resp_o[461] = 1'b0;
  assign lce_data_resp_o[462] = 1'b0;
  assign lce_data_resp_o[463] = 1'b0;
  assign lce_data_resp_o[464] = 1'b0;
  assign lce_data_resp_o[465] = 1'b0;
  assign lce_data_resp_o[466] = 1'b0;
  assign lce_data_resp_o[467] = 1'b0;
  assign lce_data_resp_o[468] = 1'b0;
  assign lce_data_resp_o[469] = 1'b0;
  assign lce_data_resp_o[470] = 1'b0;
  assign lce_data_resp_o[471] = 1'b0;
  assign lce_data_resp_o[472] = 1'b0;
  assign lce_data_resp_o[473] = 1'b0;
  assign lce_data_resp_o[474] = 1'b0;
  assign lce_data_resp_o[475] = 1'b0;
  assign lce_data_resp_o[476] = 1'b0;
  assign lce_data_resp_o[477] = 1'b0;
  assign lce_data_resp_o[478] = 1'b0;
  assign lce_data_resp_o[479] = 1'b0;
  assign lce_data_resp_o[480] = 1'b0;
  assign lce_data_resp_o[481] = 1'b0;
  assign lce_data_resp_o[482] = 1'b0;
  assign lce_data_resp_o[483] = 1'b0;
  assign lce_data_resp_o[484] = 1'b0;
  assign lce_data_resp_o[485] = 1'b0;
  assign lce_data_resp_o[486] = 1'b0;
  assign lce_data_resp_o[487] = 1'b0;
  assign lce_data_resp_o[488] = 1'b0;
  assign lce_data_resp_o[489] = 1'b0;
  assign lce_data_resp_o[490] = 1'b0;
  assign lce_data_resp_o[491] = 1'b0;
  assign lce_data_resp_o[492] = 1'b0;
  assign lce_data_resp_o[493] = 1'b0;
  assign lce_data_resp_o[494] = 1'b0;
  assign lce_data_resp_o[495] = 1'b0;
  assign lce_data_resp_o[496] = 1'b0;
  assign lce_data_resp_o[497] = 1'b0;
  assign lce_data_resp_o[498] = 1'b0;
  assign lce_data_resp_o[499] = 1'b0;
  assign lce_data_resp_o[500] = 1'b0;
  assign lce_data_resp_o[501] = 1'b0;
  assign lce_data_resp_o[502] = 1'b0;
  assign lce_data_resp_o[503] = 1'b0;
  assign lce_data_resp_o[504] = 1'b0;
  assign lce_data_resp_o[505] = 1'b0;
  assign lce_data_resp_o[506] = 1'b0;
  assign lce_data_resp_o[507] = 1'b0;
  assign lce_data_resp_o[508] = 1'b0;
  assign lce_data_resp_o[509] = 1'b0;
  assign lce_data_resp_o[510] = 1'b0;
  assign lce_data_resp_o[511] = 1'b0;
  assign lce_data_resp_o[512] = 1'b0;
  assign lce_data_resp_o[513] = 1'b0;
  assign lce_data_resp_o[514] = 1'b0;
  assign lce_data_resp_o[515] = 1'b0;
  assign lce_data_resp_o[516] = 1'b0;
  assign lce_data_resp_o[517] = 1'b0;
  assign lce_data_resp_o[518] = 1'b0;
  assign lce_data_resp_o[519] = 1'b0;
  assign lce_data_resp_o[520] = 1'b0;
  assign lce_data_resp_o[521] = 1'b0;
  assign lce_data_resp_o[522] = 1'b0;
  assign lce_data_resp_o[523] = 1'b0;
  assign lce_data_resp_o[524] = 1'b0;
  assign lce_data_resp_o[525] = 1'b0;
  assign lce_data_resp_o[526] = 1'b0;
  assign lce_data_resp_o[527] = 1'b0;
  assign lce_data_resp_o[528] = 1'b0;
  assign lce_data_resp_o[529] = 1'b0;
  assign lce_data_resp_o[530] = 1'b0;
  assign lce_data_resp_o[531] = 1'b0;
  assign lce_data_resp_o[532] = 1'b0;
  assign lce_data_resp_o[533] = 1'b0;
  assign lce_data_resp_o[534] = 1'b0;
  assign lce_data_resp_o[535] = 1'b0;
  assign lce_data_resp_o[536] = 1'b0;
  assign lce_resp_o[23] = 1'b0;
  assign lce_data_resp_o[23] = id_i[0];
  assign lce_resp_o[24] = id_i[0];
  assign N22 = state_r[1] | N21;
  assign N25 = N24 | state_r[0];
  assign N27 = N24 & N21;
  assign N28 = state_r[1] & state_r[0];
  assign lce_ready_o = state_r[0] | state_r[1];
  assign N811 = ~lce_cmd_i[31];
  assign N812 = lce_cmd_i[32] | lce_cmd_i[33];
  assign N813 = N811 | N812;
  assign N814 = ~N813;
  assign N815 = ~lce_cmd_i[33];
  assign N816 = ~lce_cmd_i[32];
  assign N817 = N816 | N815;
  assign N818 = lce_cmd_i[31] | N817;
  assign N819 = ~N818;
  assign N820 = ~syn_ack_cnt_r[0];
  assign N821 = lce_cmd_i[32] | N815;
  assign N822 = N811 | N821;
  assign N823 = ~N822;
  assign N824 = lce_cmd_i[31] | N812;
  assign N825 = ~N824;
  assign N826 = lce_cmd_i[31] | N821;
  assign N827 = ~N826;
  assign N828 = N811 | N830;
  assign N829 = ~N828;
  assign N830 = N816 | lce_cmd_i[33];
  assign N831 = lce_cmd_i[31] | N830;
  assign N832 = ~N831;
  assign N651 = syn_ack_cnt_r[0] ^ 1'b1;
  assign N37 = (N0)? 1'b0 :
               (N1)? lce_cmd_v_i : 1'b0;
  assign N0 = flag_invalidate_r;
  assign N1 = N36;
  assign N40 = (N2)? 1'b0 :
               (N667)? 1'b1 :
               (N39)? tag_mem_pkt_yumi_i : 1'b0;
  assign N2 = lce_resp_yumi_i;
  assign { N50, N49, N48, N47, N46, N45, N44, N43, N42 } = (N3)? { lce_cmd_i[20:15], lce_cmd_i[8:6] } :
                                                           (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                           (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                           (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                           (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                           (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N3 = N832;
  assign N4 = N831;
  assign N5 = 1'b0;
  assign N51 = (N3)? lce_cmd_v_i :
               (N4)? 1'b0 :
               (N5)? 1'b0 :
               (N5)? 1'b0 :
               (N5)? 1'b0 :
               (N5)? 1'b0 : 1'b0;
  assign { N53, N52 } = (N3)? { data_mem_pkt_yumi_i, N34 } :
                        (N4)? state_r : 1'b0;
  assign { N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55 } = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                      (N6)? { lce_cmd_i[34:34], 1'b1, lce_cmd_i[30:9] } :
                                                                                                                                      (N54)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                      (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                      (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                      (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N6 = N829;
  assign N79 = (N3)? 1'b0 :
               (N6)? lce_cmd_v_i :
               (N54)? 1'b0 :
               (N5)? 1'b0 :
               (N5)? 1'b0 :
               (N5)? 1'b0 : 1'b0;
  assign N80 = (N3)? 1'b0 :
               (N6)? N35 :
               (N7)? tag_mem_pkt_yumi_i :
               (N8)? tag_mem_pkt_yumi_i :
               (N9)? lce_resp_yumi_i :
               (N33)? 1'b0 : 1'b0;
  assign N7 = N827;
  assign N8 = N823;
  assign N9 = N819;
  assign { N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82 } = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                               (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                               (N7)? { lce_cmd_i[5:4], lce_cmd_i[30:21], 1'b1 } :
                                                                               (N8)? { lce_cmd_i[5:4], lce_cmd_i[30:21], 1'b1 } :
                                                                               (N81)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                               (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N103, N102, N101, N100, N99, N98, N97, N96, N95 } = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                               (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                               (N7)? { lce_cmd_i[20:15], lce_cmd_i[8:6] } :
                                                               (N8)? { lce_cmd_i[20:15], lce_cmd_i[8:6] } :
                                                               (N9)? { lce_cmd_i[20:15], lce_cmd_i[8:6] } :
                                                               (N33)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N104 = (N3)? 1'b0 :
                (N6)? 1'b0 :
                (N7)? lce_cmd_v_i :
                (N8)? lce_cmd_v_i :
                (N9)? N37 :
                (N33)? 1'b0 : 1'b0;
  assign N106 = (N3)? 1'b0 :
                (N6)? 1'b0 :
                (N7)? tag_mem_pkt_yumi_i :
                (N105)? 1'b0 :
                (N5)? 1'b0 :
                (N5)? 1'b0 : 1'b0;
  assign N107 = (N3)? 1'b0 :
                (N6)? 1'b0 :
                (N7)? 1'b0 :
                (N8)? tag_mem_pkt_yumi_i :
                (N81)? 1'b0 :
                (N5)? 1'b0 : 1'b0;
  assign N108 = (N9)? N40 :
                (N33)? flag_invalidate_r : 1'b0;
  assign { N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109 } = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                              (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                              (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                              (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                              (N9)? { lce_cmd_i[34:34], 1'b1, lce_cmd_i[30:9] } :
                                                                                                                                                              (N33)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N133 = (N3)? 1'b0 :
                (N6)? 1'b0 :
                (N7)? 1'b0 :
                (N8)? 1'b0 :
                (N9)? N41 :
                (N33)? 1'b0 : 1'b0;
  assign { N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136 } = (N10)? data_r :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N11)? data_mem_data_i : 1'b0;
  assign N10 = flag_data_buffered_r;
  assign N11 = N135;
  assign { N658, N657, N656, N655, N654, N653 } = (N12)? lce_cmd_i[20:15] :
                                                  (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                  (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = N814;
  assign N13 = N813;
  assign N659 = (N12)? lce_cmd_v_i :
                (N13)? 1'b0 :
                (N5)? 1'b0 : 1'b0;
  assign N660 = (N12)? tag_mem_pkt_yumi_i :
                (N14)? lce_resp_yumi_i :
                (N649)? 1'b0 : 1'b0;
  assign N14 = N825;
  assign N661 = (N12)? 1'b0 :
                (N14)? lce_cmd_i[34] :
                (N649)? 1'b0 : 1'b0;
  assign N662 = (N12)? 1'b0 :
                (N14)? lce_cmd_v_i :
                (N649)? 1'b0 : 1'b0;
  assign N663 = (N14)? N651 :
                (N649)? syn_ack_cnt_r[0] : 1'b0;
  assign { N665, N664 } = (N14)? { 1'b0, N652 } :
                          (N649)? state_r : 1'b0;
  assign lce_resp_v_o = (N15)? N133 :
                        (N16)? 1'b0 :
                        (N17)? N662 :
                        (N18)? 1'b0 : 1'b0;
  assign N15 = N23;
  assign N16 = N26;
  assign N17 = N27;
  assign N18 = N28;
  assign data_mem_pkt_o[521:513] = (N15)? { N50, N49, N48, N47, N46, N45, N44, N43, N42 } :
                                   (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                   (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                   (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign data_mem_pkt_v_o = (N15)? N51 :
                            (N16)? 1'b0 :
                            (N17)? 1'b0 :
                            (N18)? 1'b0 : 1'b0;
  assign state_n = (N15)? { N53, N52 } :
                   (N16)? { N134, lce_data_cmd_ready_i } :
                   (N17)? { N665, N664 } : 1'b0;
  assign { lce_data_resp_o[24:24], lce_data_resp_o[22:0] } = (N15)? { N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55 } :
                                                             (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                             (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                             (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_data_resp_v_o = (N15)? N79 :
                             (N16)? 1'b0 :
                             (N17)? 1'b0 :
                             (N18)? 1'b0 : 1'b0;
  assign lce_cmd_yumi_o = (N15)? N80 :
                          (N16)? lce_data_cmd_ready_i :
                          (N17)? N660 :
                          (N18)? 1'b0 : 1'b0;
  assign tag_mem_pkt_o = (N15)? { N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N819 } :
                         (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                         (N17)? { N658, N657, N656, N655, N654, N653, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                         (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_mem_pkt_v_o = (N15)? N104 :
                           (N16)? 1'b0 :
                           (N17)? N659 :
                           (N18)? 1'b0 : 1'b0;
  assign set_tag_received_o = (N15)? N106 :
                              (N16)? 1'b0 :
                              (N17)? 1'b0 :
                              (N18)? 1'b0 : 1'b0;
  assign set_tag_wakeup_received_o = (N15)? N107 :
                                     (N16)? 1'b0 :
                                     (N17)? 1'b0 :
                                     (N18)? 1'b0 : 1'b0;
  assign { lce_resp_o[25:25], lce_resp_o[22:0] } = (N15)? { N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109 } :
                                                   (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                   (N17)? { N661, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                   (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { lce_data_cmd_o[517:5], lce_data_cmd_o[2:0] } = (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                          (N16)? { N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, lce_cmd_i[3:0] } :
                                                          (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                          (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_data_cmd_v_o = (N15)? 1'b0 :
                            (N16)? 1'b1 :
                            (N17)? 1'b0 :
                            (N18)? 1'b0 : 1'b0;
  assign metadata_mem_pkt_o[9:4] = (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                   (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                   (N17)? { N658, N657, N656, N655, N654, N653 } :
                                   (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign metadata_mem_pkt_v_o = (N15)? 1'b0 :
                                (N16)? 1'b0 :
                                (N17)? N659 :
                                (N18)? 1'b0 : 1'b0;
  assign { N670, N669 } = (N19)? { 1'b0, 1'b0 } :
                          (N20)? state_n : 1'b0;
  assign N19 = reset_i;
  assign N20 = N668;
  assign N671 = (N19)? 1'b0 :
                (N20)? N663 : 1'b0;
  assign N672 = (N19)? 1'b0 :
                (N20)? N134 : 1'b0;
  assign N673 = (N19)? 1'b0 :
                (N20)? N108 : 1'b0;
  assign N21 = ~state_r[0];
  assign N23 = ~N22;
  assign N24 = ~state_r[1];
  assign N26 = ~N25;
  assign N29 = N829 | N832;
  assign N30 = N827 | N29;
  assign N31 = N823 | N30;
  assign N32 = N819 | N31;
  assign N33 = ~N32;
  assign N34 = ~data_mem_pkt_yumi_i;
  assign N35 = lce_data_resp_ready_i & lce_cmd_v_i;
  assign N36 = ~flag_invalidate_r;
  assign N38 = flag_invalidate_r | lce_resp_yumi_i;
  assign N39 = ~N38;
  assign N41 = flag_invalidate_r | tag_mem_pkt_yumi_i;
  assign N54 = ~N29;
  assign N81 = ~N31;
  assign N105 = ~N30;
  assign N134 = ~lce_data_cmd_ready_i;
  assign N135 = ~flag_data_buffered_r;
  assign N648 = N825 | N814;
  assign N649 = ~N648;
  assign N650 = ~lce_resp_yumi_i;
  assign N652 = N820 & lce_resp_yumi_i;
  assign N666 = ~lce_resp_yumi_i;
  assign N667 = flag_invalidate_r & N666;
  assign N668 = ~reset_i;
  assign N674 = N23 & N668;
  assign N675 = N26 & N668;
  assign N676 = flag_data_buffered_r & N675;
  assign N677 = N674 | N676;
  assign N678 = N27 & N668;
  assign N679 = N677 | N678;
  assign N680 = N28 & N668;
  assign N681 = N679 | N680;
  assign N682 = ~N681;
  assign N683 = N668 & N682;
  assign N684 = N23 & N668;
  assign N685 = N26 & N668;
  assign N686 = flag_data_buffered_r & N685;
  assign N687 = N684 | N686;
  assign N688 = N27 & N668;
  assign N689 = N687 | N688;
  assign N690 = N28 & N668;
  assign N691 = N689 | N690;
  assign N692 = ~N691;
  assign N693 = N668 & N692;
  assign N694 = N23 & N668;
  assign N695 = N26 & N668;
  assign N696 = flag_data_buffered_r & N695;
  assign N697 = N694 | N696;
  assign N698 = N27 & N668;
  assign N699 = N697 | N698;
  assign N700 = N28 & N668;
  assign N701 = N699 | N700;
  assign N702 = ~N701;
  assign N703 = N668 & N702;
  assign N704 = N23 & N668;
  assign N705 = N26 & N668;
  assign N706 = flag_data_buffered_r & N705;
  assign N707 = N704 | N706;
  assign N708 = N27 & N668;
  assign N709 = N707 | N708;
  assign N710 = N28 & N668;
  assign N711 = N709 | N710;
  assign N712 = ~N711;
  assign N713 = N668 & N712;
  assign N714 = N23 & N668;
  assign N715 = N26 & N668;
  assign N716 = flag_data_buffered_r & N715;
  assign N717 = N714 | N716;
  assign N718 = N27 & N668;
  assign N719 = N717 | N718;
  assign N720 = N28 & N668;
  assign N721 = N719 | N720;
  assign N722 = ~N721;
  assign N723 = N668 & N722;
  assign N724 = N23 & N668;
  assign N725 = N26 & N668;
  assign N726 = flag_data_buffered_r & N725;
  assign N727 = N724 | N726;
  assign N728 = N27 & N668;
  assign N729 = N727 | N728;
  assign N730 = N28 & N668;
  assign N731 = N729 | N730;
  assign N732 = ~N731;
  assign N733 = N668 & N732;
  assign N734 = N724 | N716;
  assign N735 = N734 | N728;
  assign N736 = N735 | N730;
  assign N737 = ~N736;
  assign N738 = N668 & N737;
  assign N739 = N735 | N720;
  assign N740 = ~N739;
  assign N741 = N668 & N740;
  assign N742 = N668 & N722;
  assign N743 = N714 | N706;
  assign N744 = N743 | N718;
  assign N745 = N744 | N720;
  assign N746 = ~N745;
  assign N747 = N668 & N746;
  assign N748 = N744 | N710;
  assign N749 = ~N748;
  assign N750 = N668 & N749;
  assign N751 = N668 & N712;
  assign N752 = N668 & N712;
  assign N753 = N704 | N696;
  assign N754 = N753 | N708;
  assign N755 = N754 | N710;
  assign N756 = ~N755;
  assign N757 = N668 & N756;
  assign N758 = N754 | N700;
  assign N759 = ~N758;
  assign N760 = N668 & N759;
  assign N761 = N668 & N702;
  assign N762 = N668 & N702;
  assign N763 = N694 | N686;
  assign N764 = N763 | N698;
  assign N765 = N764 | N700;
  assign N766 = ~N765;
  assign N767 = N668 & N766;
  assign N768 = N764 | N690;
  assign N769 = ~N768;
  assign N770 = N668 & N769;
  assign N771 = N668 & N692;
  assign N772 = N668 & N692;
  assign N773 = N684 | N676;
  assign N774 = N773 | N688;
  assign N775 = N774 | N690;
  assign N776 = ~N775;
  assign N777 = N668 & N776;
  assign N778 = N774 | N680;
  assign N779 = ~N778;
  assign N780 = N668 & N779;
  assign N781 = N668 & N682;
  assign N782 = N668 & N682;
  assign N783 = N668 & N682;
  assign N784 = N668 & N682;
  assign N785 = N668 & N682;
  assign N786 = N814 & N678;
  assign N787 = N786 | N680;
  assign N788 = ~N787;
  assign N789 = N674 | N675;
  assign N790 = N789 | N786;
  assign N791 = N825 & N678;
  assign N792 = N650 & N791;
  assign N793 = N790 | N792;
  assign N794 = N793 | N680;
  assign N795 = ~N794;
  assign N796 = N674 | N678;
  assign N797 = N796 | N680;
  assign N798 = ~N797;
  assign N799 = N832 & N674;
  assign N800 = N829 & N674;
  assign N801 = N799 | N800;
  assign N802 = N827 & N674;
  assign N803 = N801 | N802;
  assign N804 = N823 & N674;
  assign N805 = N803 | N804;
  assign N806 = N805 | N675;
  assign N807 = N806 | N678;
  assign N808 = N807 | N680;
  assign N809 = ~N808;

  always @(posedge clk_i) begin
    if(N683) begin
      { data_r[511:511], data_r[0:0] } <= { data_mem_data_i[511:511], data_mem_data_i[0:0] };
    end
    if(N693) begin
      { data_r[510:510] } <= { data_mem_data_i[510:510] };
    end
    if(N703) begin
      { data_r[509:509] } <= { data_mem_data_i[509:509] };
    end
    if(N713) begin
      { data_r[508:508] } <= { data_mem_data_i[508:508] };
    end
    if(N723) begin
      { data_r[507:507], data_r[488:413] } <= { data_mem_data_i[507:507], data_mem_data_i[488:413] };
    end
    if(N733) begin
      { data_r[506:493] } <= { data_mem_data_i[506:493] };
    end
    if(N738) begin
      { data_r[492:490] } <= { data_mem_data_i[492:490] };
    end
    if(N741) begin
      { data_r[489:489] } <= { data_mem_data_i[489:489] };
    end
    if(N742) begin
      { data_r[412:394] } <= { data_mem_data_i[412:394] };
    end
    if(N747) begin
      { data_r[393:391] } <= { data_mem_data_i[393:391] };
    end
    if(N750) begin
      { data_r[390:390] } <= { data_mem_data_i[390:390] };
    end
    if(N751) begin
      { data_r[389:314] } <= { data_mem_data_i[389:314] };
    end
    if(N752) begin
      { data_r[313:295] } <= { data_mem_data_i[313:295] };
    end
    if(N757) begin
      { data_r[294:292] } <= { data_mem_data_i[294:292] };
    end
    if(N760) begin
      { data_r[291:291] } <= { data_mem_data_i[291:291] };
    end
    if(N761) begin
      { data_r[290:215] } <= { data_mem_data_i[290:215] };
    end
    if(N762) begin
      { data_r[214:196] } <= { data_mem_data_i[214:196] };
    end
    if(N767) begin
      { data_r[195:193] } <= { data_mem_data_i[195:193] };
    end
    if(N770) begin
      { data_r[192:192] } <= { data_mem_data_i[192:192] };
    end
    if(N771) begin
      { data_r[191:116] } <= { data_mem_data_i[191:116] };
    end
    if(N772) begin
      { data_r[115:97] } <= { data_mem_data_i[115:97] };
    end
    if(N777) begin
      { data_r[96:94] } <= { data_mem_data_i[96:94] };
    end
    if(N780) begin
      { data_r[93:93] } <= { data_mem_data_i[93:93] };
    end
    if(N781) begin
      { data_r[92:17], data_r[4:4] } <= { data_mem_data_i[92:17], data_mem_data_i[4:4] };
    end
    if(N782) begin
      { data_r[16:5] } <= { data_mem_data_i[16:5] };
    end
    if(N783) begin
      { data_r[3:3] } <= { data_mem_data_i[3:3] };
    end
    if(N784) begin
      { data_r[2:2] } <= { data_mem_data_i[2:2] };
    end
    if(N785) begin
      { data_r[1:1] } <= { data_mem_data_i[1:1] };
    end
    if(N788) begin
      { state_r[1:0] } <= { N670, N669 };
    end
    if(N795) begin
      { syn_ack_cnt_r[0:0] } <= { N671 };
    end
    if(N798) begin
      flag_data_buffered_r <= N672;
    end
    if(N809) begin
      flag_invalidate_r <= N673;
    end
  end


endmodule



module bp_fe_lce_data_cmd_data_width_p64_paddr_width_p22_lce_data_width_p512_num_cce_p1_num_lce_p2_sets_p64_ways_p8
(
  cce_data_received_o,
  tr_data_received_o,
  miss_addr_i,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_yumi_o,
  data_mem_pkt_v_o,
  data_mem_pkt_o,
  data_mem_pkt_yumi_i
);

  input [21:0] miss_addr_i;
  input [517:0] lce_data_cmd_i;
  output [521:0] data_mem_pkt_o;
  input lce_data_cmd_v_i;
  input data_mem_pkt_yumi_i;
  output cce_data_received_o;
  output tr_data_received_o;
  output lce_data_cmd_yumi_o;
  output data_mem_pkt_v_o;
  wire [521:0] data_mem_pkt_o;
  wire cce_data_received_o,tr_data_received_o,lce_data_cmd_yumi_o,data_mem_pkt_v_o,
  data_mem_pkt_yumi_i,lce_data_cmd_v_i,N0,N1,N2,N3,N4;
  assign data_mem_pkt_o[512] = 1'b1;
  assign data_mem_pkt_o[515] = lce_data_cmd_i[2];
  assign data_mem_pkt_o[514] = lce_data_cmd_i[1];
  assign data_mem_pkt_o[513] = lce_data_cmd_i[0];
  assign data_mem_pkt_o[511] = lce_data_cmd_i[517];
  assign data_mem_pkt_o[510] = lce_data_cmd_i[516];
  assign data_mem_pkt_o[509] = lce_data_cmd_i[515];
  assign data_mem_pkt_o[508] = lce_data_cmd_i[514];
  assign data_mem_pkt_o[507] = lce_data_cmd_i[513];
  assign data_mem_pkt_o[506] = lce_data_cmd_i[512];
  assign data_mem_pkt_o[505] = lce_data_cmd_i[511];
  assign data_mem_pkt_o[504] = lce_data_cmd_i[510];
  assign data_mem_pkt_o[503] = lce_data_cmd_i[509];
  assign data_mem_pkt_o[502] = lce_data_cmd_i[508];
  assign data_mem_pkt_o[501] = lce_data_cmd_i[507];
  assign data_mem_pkt_o[500] = lce_data_cmd_i[506];
  assign data_mem_pkt_o[499] = lce_data_cmd_i[505];
  assign data_mem_pkt_o[498] = lce_data_cmd_i[504];
  assign data_mem_pkt_o[497] = lce_data_cmd_i[503];
  assign data_mem_pkt_o[496] = lce_data_cmd_i[502];
  assign data_mem_pkt_o[495] = lce_data_cmd_i[501];
  assign data_mem_pkt_o[494] = lce_data_cmd_i[500];
  assign data_mem_pkt_o[493] = lce_data_cmd_i[499];
  assign data_mem_pkt_o[492] = lce_data_cmd_i[498];
  assign data_mem_pkt_o[491] = lce_data_cmd_i[497];
  assign data_mem_pkt_o[490] = lce_data_cmd_i[496];
  assign data_mem_pkt_o[489] = lce_data_cmd_i[495];
  assign data_mem_pkt_o[488] = lce_data_cmd_i[494];
  assign data_mem_pkt_o[487] = lce_data_cmd_i[493];
  assign data_mem_pkt_o[486] = lce_data_cmd_i[492];
  assign data_mem_pkt_o[485] = lce_data_cmd_i[491];
  assign data_mem_pkt_o[484] = lce_data_cmd_i[490];
  assign data_mem_pkt_o[483] = lce_data_cmd_i[489];
  assign data_mem_pkt_o[482] = lce_data_cmd_i[488];
  assign data_mem_pkt_o[481] = lce_data_cmd_i[487];
  assign data_mem_pkt_o[480] = lce_data_cmd_i[486];
  assign data_mem_pkt_o[479] = lce_data_cmd_i[485];
  assign data_mem_pkt_o[478] = lce_data_cmd_i[484];
  assign data_mem_pkt_o[477] = lce_data_cmd_i[483];
  assign data_mem_pkt_o[476] = lce_data_cmd_i[482];
  assign data_mem_pkt_o[475] = lce_data_cmd_i[481];
  assign data_mem_pkt_o[474] = lce_data_cmd_i[480];
  assign data_mem_pkt_o[473] = lce_data_cmd_i[479];
  assign data_mem_pkt_o[472] = lce_data_cmd_i[478];
  assign data_mem_pkt_o[471] = lce_data_cmd_i[477];
  assign data_mem_pkt_o[470] = lce_data_cmd_i[476];
  assign data_mem_pkt_o[469] = lce_data_cmd_i[475];
  assign data_mem_pkt_o[468] = lce_data_cmd_i[474];
  assign data_mem_pkt_o[467] = lce_data_cmd_i[473];
  assign data_mem_pkt_o[466] = lce_data_cmd_i[472];
  assign data_mem_pkt_o[465] = lce_data_cmd_i[471];
  assign data_mem_pkt_o[464] = lce_data_cmd_i[470];
  assign data_mem_pkt_o[463] = lce_data_cmd_i[469];
  assign data_mem_pkt_o[462] = lce_data_cmd_i[468];
  assign data_mem_pkt_o[461] = lce_data_cmd_i[467];
  assign data_mem_pkt_o[460] = lce_data_cmd_i[466];
  assign data_mem_pkt_o[459] = lce_data_cmd_i[465];
  assign data_mem_pkt_o[458] = lce_data_cmd_i[464];
  assign data_mem_pkt_o[457] = lce_data_cmd_i[463];
  assign data_mem_pkt_o[456] = lce_data_cmd_i[462];
  assign data_mem_pkt_o[455] = lce_data_cmd_i[461];
  assign data_mem_pkt_o[454] = lce_data_cmd_i[460];
  assign data_mem_pkt_o[453] = lce_data_cmd_i[459];
  assign data_mem_pkt_o[452] = lce_data_cmd_i[458];
  assign data_mem_pkt_o[451] = lce_data_cmd_i[457];
  assign data_mem_pkt_o[450] = lce_data_cmd_i[456];
  assign data_mem_pkt_o[449] = lce_data_cmd_i[455];
  assign data_mem_pkt_o[448] = lce_data_cmd_i[454];
  assign data_mem_pkt_o[447] = lce_data_cmd_i[453];
  assign data_mem_pkt_o[446] = lce_data_cmd_i[452];
  assign data_mem_pkt_o[445] = lce_data_cmd_i[451];
  assign data_mem_pkt_o[444] = lce_data_cmd_i[450];
  assign data_mem_pkt_o[443] = lce_data_cmd_i[449];
  assign data_mem_pkt_o[442] = lce_data_cmd_i[448];
  assign data_mem_pkt_o[441] = lce_data_cmd_i[447];
  assign data_mem_pkt_o[440] = lce_data_cmd_i[446];
  assign data_mem_pkt_o[439] = lce_data_cmd_i[445];
  assign data_mem_pkt_o[438] = lce_data_cmd_i[444];
  assign data_mem_pkt_o[437] = lce_data_cmd_i[443];
  assign data_mem_pkt_o[436] = lce_data_cmd_i[442];
  assign data_mem_pkt_o[435] = lce_data_cmd_i[441];
  assign data_mem_pkt_o[434] = lce_data_cmd_i[440];
  assign data_mem_pkt_o[433] = lce_data_cmd_i[439];
  assign data_mem_pkt_o[432] = lce_data_cmd_i[438];
  assign data_mem_pkt_o[431] = lce_data_cmd_i[437];
  assign data_mem_pkt_o[430] = lce_data_cmd_i[436];
  assign data_mem_pkt_o[429] = lce_data_cmd_i[435];
  assign data_mem_pkt_o[428] = lce_data_cmd_i[434];
  assign data_mem_pkt_o[427] = lce_data_cmd_i[433];
  assign data_mem_pkt_o[426] = lce_data_cmd_i[432];
  assign data_mem_pkt_o[425] = lce_data_cmd_i[431];
  assign data_mem_pkt_o[424] = lce_data_cmd_i[430];
  assign data_mem_pkt_o[423] = lce_data_cmd_i[429];
  assign data_mem_pkt_o[422] = lce_data_cmd_i[428];
  assign data_mem_pkt_o[421] = lce_data_cmd_i[427];
  assign data_mem_pkt_o[420] = lce_data_cmd_i[426];
  assign data_mem_pkt_o[419] = lce_data_cmd_i[425];
  assign data_mem_pkt_o[418] = lce_data_cmd_i[424];
  assign data_mem_pkt_o[417] = lce_data_cmd_i[423];
  assign data_mem_pkt_o[416] = lce_data_cmd_i[422];
  assign data_mem_pkt_o[415] = lce_data_cmd_i[421];
  assign data_mem_pkt_o[414] = lce_data_cmd_i[420];
  assign data_mem_pkt_o[413] = lce_data_cmd_i[419];
  assign data_mem_pkt_o[412] = lce_data_cmd_i[418];
  assign data_mem_pkt_o[411] = lce_data_cmd_i[417];
  assign data_mem_pkt_o[410] = lce_data_cmd_i[416];
  assign data_mem_pkt_o[409] = lce_data_cmd_i[415];
  assign data_mem_pkt_o[408] = lce_data_cmd_i[414];
  assign data_mem_pkt_o[407] = lce_data_cmd_i[413];
  assign data_mem_pkt_o[406] = lce_data_cmd_i[412];
  assign data_mem_pkt_o[405] = lce_data_cmd_i[411];
  assign data_mem_pkt_o[404] = lce_data_cmd_i[410];
  assign data_mem_pkt_o[403] = lce_data_cmd_i[409];
  assign data_mem_pkt_o[402] = lce_data_cmd_i[408];
  assign data_mem_pkt_o[401] = lce_data_cmd_i[407];
  assign data_mem_pkt_o[400] = lce_data_cmd_i[406];
  assign data_mem_pkt_o[399] = lce_data_cmd_i[405];
  assign data_mem_pkt_o[398] = lce_data_cmd_i[404];
  assign data_mem_pkt_o[397] = lce_data_cmd_i[403];
  assign data_mem_pkt_o[396] = lce_data_cmd_i[402];
  assign data_mem_pkt_o[395] = lce_data_cmd_i[401];
  assign data_mem_pkt_o[394] = lce_data_cmd_i[400];
  assign data_mem_pkt_o[393] = lce_data_cmd_i[399];
  assign data_mem_pkt_o[392] = lce_data_cmd_i[398];
  assign data_mem_pkt_o[391] = lce_data_cmd_i[397];
  assign data_mem_pkt_o[390] = lce_data_cmd_i[396];
  assign data_mem_pkt_o[389] = lce_data_cmd_i[395];
  assign data_mem_pkt_o[388] = lce_data_cmd_i[394];
  assign data_mem_pkt_o[387] = lce_data_cmd_i[393];
  assign data_mem_pkt_o[386] = lce_data_cmd_i[392];
  assign data_mem_pkt_o[385] = lce_data_cmd_i[391];
  assign data_mem_pkt_o[384] = lce_data_cmd_i[390];
  assign data_mem_pkt_o[383] = lce_data_cmd_i[389];
  assign data_mem_pkt_o[382] = lce_data_cmd_i[388];
  assign data_mem_pkt_o[381] = lce_data_cmd_i[387];
  assign data_mem_pkt_o[380] = lce_data_cmd_i[386];
  assign data_mem_pkt_o[379] = lce_data_cmd_i[385];
  assign data_mem_pkt_o[378] = lce_data_cmd_i[384];
  assign data_mem_pkt_o[377] = lce_data_cmd_i[383];
  assign data_mem_pkt_o[376] = lce_data_cmd_i[382];
  assign data_mem_pkt_o[375] = lce_data_cmd_i[381];
  assign data_mem_pkt_o[374] = lce_data_cmd_i[380];
  assign data_mem_pkt_o[373] = lce_data_cmd_i[379];
  assign data_mem_pkt_o[372] = lce_data_cmd_i[378];
  assign data_mem_pkt_o[371] = lce_data_cmd_i[377];
  assign data_mem_pkt_o[370] = lce_data_cmd_i[376];
  assign data_mem_pkt_o[369] = lce_data_cmd_i[375];
  assign data_mem_pkt_o[368] = lce_data_cmd_i[374];
  assign data_mem_pkt_o[367] = lce_data_cmd_i[373];
  assign data_mem_pkt_o[366] = lce_data_cmd_i[372];
  assign data_mem_pkt_o[365] = lce_data_cmd_i[371];
  assign data_mem_pkt_o[364] = lce_data_cmd_i[370];
  assign data_mem_pkt_o[363] = lce_data_cmd_i[369];
  assign data_mem_pkt_o[362] = lce_data_cmd_i[368];
  assign data_mem_pkt_o[361] = lce_data_cmd_i[367];
  assign data_mem_pkt_o[360] = lce_data_cmd_i[366];
  assign data_mem_pkt_o[359] = lce_data_cmd_i[365];
  assign data_mem_pkt_o[358] = lce_data_cmd_i[364];
  assign data_mem_pkt_o[357] = lce_data_cmd_i[363];
  assign data_mem_pkt_o[356] = lce_data_cmd_i[362];
  assign data_mem_pkt_o[355] = lce_data_cmd_i[361];
  assign data_mem_pkt_o[354] = lce_data_cmd_i[360];
  assign data_mem_pkt_o[353] = lce_data_cmd_i[359];
  assign data_mem_pkt_o[352] = lce_data_cmd_i[358];
  assign data_mem_pkt_o[351] = lce_data_cmd_i[357];
  assign data_mem_pkt_o[350] = lce_data_cmd_i[356];
  assign data_mem_pkt_o[349] = lce_data_cmd_i[355];
  assign data_mem_pkt_o[348] = lce_data_cmd_i[354];
  assign data_mem_pkt_o[347] = lce_data_cmd_i[353];
  assign data_mem_pkt_o[346] = lce_data_cmd_i[352];
  assign data_mem_pkt_o[345] = lce_data_cmd_i[351];
  assign data_mem_pkt_o[344] = lce_data_cmd_i[350];
  assign data_mem_pkt_o[343] = lce_data_cmd_i[349];
  assign data_mem_pkt_o[342] = lce_data_cmd_i[348];
  assign data_mem_pkt_o[341] = lce_data_cmd_i[347];
  assign data_mem_pkt_o[340] = lce_data_cmd_i[346];
  assign data_mem_pkt_o[339] = lce_data_cmd_i[345];
  assign data_mem_pkt_o[338] = lce_data_cmd_i[344];
  assign data_mem_pkt_o[337] = lce_data_cmd_i[343];
  assign data_mem_pkt_o[336] = lce_data_cmd_i[342];
  assign data_mem_pkt_o[335] = lce_data_cmd_i[341];
  assign data_mem_pkt_o[334] = lce_data_cmd_i[340];
  assign data_mem_pkt_o[333] = lce_data_cmd_i[339];
  assign data_mem_pkt_o[332] = lce_data_cmd_i[338];
  assign data_mem_pkt_o[331] = lce_data_cmd_i[337];
  assign data_mem_pkt_o[330] = lce_data_cmd_i[336];
  assign data_mem_pkt_o[329] = lce_data_cmd_i[335];
  assign data_mem_pkt_o[328] = lce_data_cmd_i[334];
  assign data_mem_pkt_o[327] = lce_data_cmd_i[333];
  assign data_mem_pkt_o[326] = lce_data_cmd_i[332];
  assign data_mem_pkt_o[325] = lce_data_cmd_i[331];
  assign data_mem_pkt_o[324] = lce_data_cmd_i[330];
  assign data_mem_pkt_o[323] = lce_data_cmd_i[329];
  assign data_mem_pkt_o[322] = lce_data_cmd_i[328];
  assign data_mem_pkt_o[321] = lce_data_cmd_i[327];
  assign data_mem_pkt_o[320] = lce_data_cmd_i[326];
  assign data_mem_pkt_o[319] = lce_data_cmd_i[325];
  assign data_mem_pkt_o[318] = lce_data_cmd_i[324];
  assign data_mem_pkt_o[317] = lce_data_cmd_i[323];
  assign data_mem_pkt_o[316] = lce_data_cmd_i[322];
  assign data_mem_pkt_o[315] = lce_data_cmd_i[321];
  assign data_mem_pkt_o[314] = lce_data_cmd_i[320];
  assign data_mem_pkt_o[313] = lce_data_cmd_i[319];
  assign data_mem_pkt_o[312] = lce_data_cmd_i[318];
  assign data_mem_pkt_o[311] = lce_data_cmd_i[317];
  assign data_mem_pkt_o[310] = lce_data_cmd_i[316];
  assign data_mem_pkt_o[309] = lce_data_cmd_i[315];
  assign data_mem_pkt_o[308] = lce_data_cmd_i[314];
  assign data_mem_pkt_o[307] = lce_data_cmd_i[313];
  assign data_mem_pkt_o[306] = lce_data_cmd_i[312];
  assign data_mem_pkt_o[305] = lce_data_cmd_i[311];
  assign data_mem_pkt_o[304] = lce_data_cmd_i[310];
  assign data_mem_pkt_o[303] = lce_data_cmd_i[309];
  assign data_mem_pkt_o[302] = lce_data_cmd_i[308];
  assign data_mem_pkt_o[301] = lce_data_cmd_i[307];
  assign data_mem_pkt_o[300] = lce_data_cmd_i[306];
  assign data_mem_pkt_o[299] = lce_data_cmd_i[305];
  assign data_mem_pkt_o[298] = lce_data_cmd_i[304];
  assign data_mem_pkt_o[297] = lce_data_cmd_i[303];
  assign data_mem_pkt_o[296] = lce_data_cmd_i[302];
  assign data_mem_pkt_o[295] = lce_data_cmd_i[301];
  assign data_mem_pkt_o[294] = lce_data_cmd_i[300];
  assign data_mem_pkt_o[293] = lce_data_cmd_i[299];
  assign data_mem_pkt_o[292] = lce_data_cmd_i[298];
  assign data_mem_pkt_o[291] = lce_data_cmd_i[297];
  assign data_mem_pkt_o[290] = lce_data_cmd_i[296];
  assign data_mem_pkt_o[289] = lce_data_cmd_i[295];
  assign data_mem_pkt_o[288] = lce_data_cmd_i[294];
  assign data_mem_pkt_o[287] = lce_data_cmd_i[293];
  assign data_mem_pkt_o[286] = lce_data_cmd_i[292];
  assign data_mem_pkt_o[285] = lce_data_cmd_i[291];
  assign data_mem_pkt_o[284] = lce_data_cmd_i[290];
  assign data_mem_pkt_o[283] = lce_data_cmd_i[289];
  assign data_mem_pkt_o[282] = lce_data_cmd_i[288];
  assign data_mem_pkt_o[281] = lce_data_cmd_i[287];
  assign data_mem_pkt_o[280] = lce_data_cmd_i[286];
  assign data_mem_pkt_o[279] = lce_data_cmd_i[285];
  assign data_mem_pkt_o[278] = lce_data_cmd_i[284];
  assign data_mem_pkt_o[277] = lce_data_cmd_i[283];
  assign data_mem_pkt_o[276] = lce_data_cmd_i[282];
  assign data_mem_pkt_o[275] = lce_data_cmd_i[281];
  assign data_mem_pkt_o[274] = lce_data_cmd_i[280];
  assign data_mem_pkt_o[273] = lce_data_cmd_i[279];
  assign data_mem_pkt_o[272] = lce_data_cmd_i[278];
  assign data_mem_pkt_o[271] = lce_data_cmd_i[277];
  assign data_mem_pkt_o[270] = lce_data_cmd_i[276];
  assign data_mem_pkt_o[269] = lce_data_cmd_i[275];
  assign data_mem_pkt_o[268] = lce_data_cmd_i[274];
  assign data_mem_pkt_o[267] = lce_data_cmd_i[273];
  assign data_mem_pkt_o[266] = lce_data_cmd_i[272];
  assign data_mem_pkt_o[265] = lce_data_cmd_i[271];
  assign data_mem_pkt_o[264] = lce_data_cmd_i[270];
  assign data_mem_pkt_o[263] = lce_data_cmd_i[269];
  assign data_mem_pkt_o[262] = lce_data_cmd_i[268];
  assign data_mem_pkt_o[261] = lce_data_cmd_i[267];
  assign data_mem_pkt_o[260] = lce_data_cmd_i[266];
  assign data_mem_pkt_o[259] = lce_data_cmd_i[265];
  assign data_mem_pkt_o[258] = lce_data_cmd_i[264];
  assign data_mem_pkt_o[257] = lce_data_cmd_i[263];
  assign data_mem_pkt_o[256] = lce_data_cmd_i[262];
  assign data_mem_pkt_o[255] = lce_data_cmd_i[261];
  assign data_mem_pkt_o[254] = lce_data_cmd_i[260];
  assign data_mem_pkt_o[253] = lce_data_cmd_i[259];
  assign data_mem_pkt_o[252] = lce_data_cmd_i[258];
  assign data_mem_pkt_o[251] = lce_data_cmd_i[257];
  assign data_mem_pkt_o[250] = lce_data_cmd_i[256];
  assign data_mem_pkt_o[249] = lce_data_cmd_i[255];
  assign data_mem_pkt_o[248] = lce_data_cmd_i[254];
  assign data_mem_pkt_o[247] = lce_data_cmd_i[253];
  assign data_mem_pkt_o[246] = lce_data_cmd_i[252];
  assign data_mem_pkt_o[245] = lce_data_cmd_i[251];
  assign data_mem_pkt_o[244] = lce_data_cmd_i[250];
  assign data_mem_pkt_o[243] = lce_data_cmd_i[249];
  assign data_mem_pkt_o[242] = lce_data_cmd_i[248];
  assign data_mem_pkt_o[241] = lce_data_cmd_i[247];
  assign data_mem_pkt_o[240] = lce_data_cmd_i[246];
  assign data_mem_pkt_o[239] = lce_data_cmd_i[245];
  assign data_mem_pkt_o[238] = lce_data_cmd_i[244];
  assign data_mem_pkt_o[237] = lce_data_cmd_i[243];
  assign data_mem_pkt_o[236] = lce_data_cmd_i[242];
  assign data_mem_pkt_o[235] = lce_data_cmd_i[241];
  assign data_mem_pkt_o[234] = lce_data_cmd_i[240];
  assign data_mem_pkt_o[233] = lce_data_cmd_i[239];
  assign data_mem_pkt_o[232] = lce_data_cmd_i[238];
  assign data_mem_pkt_o[231] = lce_data_cmd_i[237];
  assign data_mem_pkt_o[230] = lce_data_cmd_i[236];
  assign data_mem_pkt_o[229] = lce_data_cmd_i[235];
  assign data_mem_pkt_o[228] = lce_data_cmd_i[234];
  assign data_mem_pkt_o[227] = lce_data_cmd_i[233];
  assign data_mem_pkt_o[226] = lce_data_cmd_i[232];
  assign data_mem_pkt_o[225] = lce_data_cmd_i[231];
  assign data_mem_pkt_o[224] = lce_data_cmd_i[230];
  assign data_mem_pkt_o[223] = lce_data_cmd_i[229];
  assign data_mem_pkt_o[222] = lce_data_cmd_i[228];
  assign data_mem_pkt_o[221] = lce_data_cmd_i[227];
  assign data_mem_pkt_o[220] = lce_data_cmd_i[226];
  assign data_mem_pkt_o[219] = lce_data_cmd_i[225];
  assign data_mem_pkt_o[218] = lce_data_cmd_i[224];
  assign data_mem_pkt_o[217] = lce_data_cmd_i[223];
  assign data_mem_pkt_o[216] = lce_data_cmd_i[222];
  assign data_mem_pkt_o[215] = lce_data_cmd_i[221];
  assign data_mem_pkt_o[214] = lce_data_cmd_i[220];
  assign data_mem_pkt_o[213] = lce_data_cmd_i[219];
  assign data_mem_pkt_o[212] = lce_data_cmd_i[218];
  assign data_mem_pkt_o[211] = lce_data_cmd_i[217];
  assign data_mem_pkt_o[210] = lce_data_cmd_i[216];
  assign data_mem_pkt_o[209] = lce_data_cmd_i[215];
  assign data_mem_pkt_o[208] = lce_data_cmd_i[214];
  assign data_mem_pkt_o[207] = lce_data_cmd_i[213];
  assign data_mem_pkt_o[206] = lce_data_cmd_i[212];
  assign data_mem_pkt_o[205] = lce_data_cmd_i[211];
  assign data_mem_pkt_o[204] = lce_data_cmd_i[210];
  assign data_mem_pkt_o[203] = lce_data_cmd_i[209];
  assign data_mem_pkt_o[202] = lce_data_cmd_i[208];
  assign data_mem_pkt_o[201] = lce_data_cmd_i[207];
  assign data_mem_pkt_o[200] = lce_data_cmd_i[206];
  assign data_mem_pkt_o[199] = lce_data_cmd_i[205];
  assign data_mem_pkt_o[198] = lce_data_cmd_i[204];
  assign data_mem_pkt_o[197] = lce_data_cmd_i[203];
  assign data_mem_pkt_o[196] = lce_data_cmd_i[202];
  assign data_mem_pkt_o[195] = lce_data_cmd_i[201];
  assign data_mem_pkt_o[194] = lce_data_cmd_i[200];
  assign data_mem_pkt_o[193] = lce_data_cmd_i[199];
  assign data_mem_pkt_o[192] = lce_data_cmd_i[198];
  assign data_mem_pkt_o[191] = lce_data_cmd_i[197];
  assign data_mem_pkt_o[190] = lce_data_cmd_i[196];
  assign data_mem_pkt_o[189] = lce_data_cmd_i[195];
  assign data_mem_pkt_o[188] = lce_data_cmd_i[194];
  assign data_mem_pkt_o[187] = lce_data_cmd_i[193];
  assign data_mem_pkt_o[186] = lce_data_cmd_i[192];
  assign data_mem_pkt_o[185] = lce_data_cmd_i[191];
  assign data_mem_pkt_o[184] = lce_data_cmd_i[190];
  assign data_mem_pkt_o[183] = lce_data_cmd_i[189];
  assign data_mem_pkt_o[182] = lce_data_cmd_i[188];
  assign data_mem_pkt_o[181] = lce_data_cmd_i[187];
  assign data_mem_pkt_o[180] = lce_data_cmd_i[186];
  assign data_mem_pkt_o[179] = lce_data_cmd_i[185];
  assign data_mem_pkt_o[178] = lce_data_cmd_i[184];
  assign data_mem_pkt_o[177] = lce_data_cmd_i[183];
  assign data_mem_pkt_o[176] = lce_data_cmd_i[182];
  assign data_mem_pkt_o[175] = lce_data_cmd_i[181];
  assign data_mem_pkt_o[174] = lce_data_cmd_i[180];
  assign data_mem_pkt_o[173] = lce_data_cmd_i[179];
  assign data_mem_pkt_o[172] = lce_data_cmd_i[178];
  assign data_mem_pkt_o[171] = lce_data_cmd_i[177];
  assign data_mem_pkt_o[170] = lce_data_cmd_i[176];
  assign data_mem_pkt_o[169] = lce_data_cmd_i[175];
  assign data_mem_pkt_o[168] = lce_data_cmd_i[174];
  assign data_mem_pkt_o[167] = lce_data_cmd_i[173];
  assign data_mem_pkt_o[166] = lce_data_cmd_i[172];
  assign data_mem_pkt_o[165] = lce_data_cmd_i[171];
  assign data_mem_pkt_o[164] = lce_data_cmd_i[170];
  assign data_mem_pkt_o[163] = lce_data_cmd_i[169];
  assign data_mem_pkt_o[162] = lce_data_cmd_i[168];
  assign data_mem_pkt_o[161] = lce_data_cmd_i[167];
  assign data_mem_pkt_o[160] = lce_data_cmd_i[166];
  assign data_mem_pkt_o[159] = lce_data_cmd_i[165];
  assign data_mem_pkt_o[158] = lce_data_cmd_i[164];
  assign data_mem_pkt_o[157] = lce_data_cmd_i[163];
  assign data_mem_pkt_o[156] = lce_data_cmd_i[162];
  assign data_mem_pkt_o[155] = lce_data_cmd_i[161];
  assign data_mem_pkt_o[154] = lce_data_cmd_i[160];
  assign data_mem_pkt_o[153] = lce_data_cmd_i[159];
  assign data_mem_pkt_o[152] = lce_data_cmd_i[158];
  assign data_mem_pkt_o[151] = lce_data_cmd_i[157];
  assign data_mem_pkt_o[150] = lce_data_cmd_i[156];
  assign data_mem_pkt_o[149] = lce_data_cmd_i[155];
  assign data_mem_pkt_o[148] = lce_data_cmd_i[154];
  assign data_mem_pkt_o[147] = lce_data_cmd_i[153];
  assign data_mem_pkt_o[146] = lce_data_cmd_i[152];
  assign data_mem_pkt_o[145] = lce_data_cmd_i[151];
  assign data_mem_pkt_o[144] = lce_data_cmd_i[150];
  assign data_mem_pkt_o[143] = lce_data_cmd_i[149];
  assign data_mem_pkt_o[142] = lce_data_cmd_i[148];
  assign data_mem_pkt_o[141] = lce_data_cmd_i[147];
  assign data_mem_pkt_o[140] = lce_data_cmd_i[146];
  assign data_mem_pkt_o[139] = lce_data_cmd_i[145];
  assign data_mem_pkt_o[138] = lce_data_cmd_i[144];
  assign data_mem_pkt_o[137] = lce_data_cmd_i[143];
  assign data_mem_pkt_o[136] = lce_data_cmd_i[142];
  assign data_mem_pkt_o[135] = lce_data_cmd_i[141];
  assign data_mem_pkt_o[134] = lce_data_cmd_i[140];
  assign data_mem_pkt_o[133] = lce_data_cmd_i[139];
  assign data_mem_pkt_o[132] = lce_data_cmd_i[138];
  assign data_mem_pkt_o[131] = lce_data_cmd_i[137];
  assign data_mem_pkt_o[130] = lce_data_cmd_i[136];
  assign data_mem_pkt_o[129] = lce_data_cmd_i[135];
  assign data_mem_pkt_o[128] = lce_data_cmd_i[134];
  assign data_mem_pkt_o[127] = lce_data_cmd_i[133];
  assign data_mem_pkt_o[126] = lce_data_cmd_i[132];
  assign data_mem_pkt_o[125] = lce_data_cmd_i[131];
  assign data_mem_pkt_o[124] = lce_data_cmd_i[130];
  assign data_mem_pkt_o[123] = lce_data_cmd_i[129];
  assign data_mem_pkt_o[122] = lce_data_cmd_i[128];
  assign data_mem_pkt_o[121] = lce_data_cmd_i[127];
  assign data_mem_pkt_o[120] = lce_data_cmd_i[126];
  assign data_mem_pkt_o[119] = lce_data_cmd_i[125];
  assign data_mem_pkt_o[118] = lce_data_cmd_i[124];
  assign data_mem_pkt_o[117] = lce_data_cmd_i[123];
  assign data_mem_pkt_o[116] = lce_data_cmd_i[122];
  assign data_mem_pkt_o[115] = lce_data_cmd_i[121];
  assign data_mem_pkt_o[114] = lce_data_cmd_i[120];
  assign data_mem_pkt_o[113] = lce_data_cmd_i[119];
  assign data_mem_pkt_o[112] = lce_data_cmd_i[118];
  assign data_mem_pkt_o[111] = lce_data_cmd_i[117];
  assign data_mem_pkt_o[110] = lce_data_cmd_i[116];
  assign data_mem_pkt_o[109] = lce_data_cmd_i[115];
  assign data_mem_pkt_o[108] = lce_data_cmd_i[114];
  assign data_mem_pkt_o[107] = lce_data_cmd_i[113];
  assign data_mem_pkt_o[106] = lce_data_cmd_i[112];
  assign data_mem_pkt_o[105] = lce_data_cmd_i[111];
  assign data_mem_pkt_o[104] = lce_data_cmd_i[110];
  assign data_mem_pkt_o[103] = lce_data_cmd_i[109];
  assign data_mem_pkt_o[102] = lce_data_cmd_i[108];
  assign data_mem_pkt_o[101] = lce_data_cmd_i[107];
  assign data_mem_pkt_o[100] = lce_data_cmd_i[106];
  assign data_mem_pkt_o[99] = lce_data_cmd_i[105];
  assign data_mem_pkt_o[98] = lce_data_cmd_i[104];
  assign data_mem_pkt_o[97] = lce_data_cmd_i[103];
  assign data_mem_pkt_o[96] = lce_data_cmd_i[102];
  assign data_mem_pkt_o[95] = lce_data_cmd_i[101];
  assign data_mem_pkt_o[94] = lce_data_cmd_i[100];
  assign data_mem_pkt_o[93] = lce_data_cmd_i[99];
  assign data_mem_pkt_o[92] = lce_data_cmd_i[98];
  assign data_mem_pkt_o[91] = lce_data_cmd_i[97];
  assign data_mem_pkt_o[90] = lce_data_cmd_i[96];
  assign data_mem_pkt_o[89] = lce_data_cmd_i[95];
  assign data_mem_pkt_o[88] = lce_data_cmd_i[94];
  assign data_mem_pkt_o[87] = lce_data_cmd_i[93];
  assign data_mem_pkt_o[86] = lce_data_cmd_i[92];
  assign data_mem_pkt_o[85] = lce_data_cmd_i[91];
  assign data_mem_pkt_o[84] = lce_data_cmd_i[90];
  assign data_mem_pkt_o[83] = lce_data_cmd_i[89];
  assign data_mem_pkt_o[82] = lce_data_cmd_i[88];
  assign data_mem_pkt_o[81] = lce_data_cmd_i[87];
  assign data_mem_pkt_o[80] = lce_data_cmd_i[86];
  assign data_mem_pkt_o[79] = lce_data_cmd_i[85];
  assign data_mem_pkt_o[78] = lce_data_cmd_i[84];
  assign data_mem_pkt_o[77] = lce_data_cmd_i[83];
  assign data_mem_pkt_o[76] = lce_data_cmd_i[82];
  assign data_mem_pkt_o[75] = lce_data_cmd_i[81];
  assign data_mem_pkt_o[74] = lce_data_cmd_i[80];
  assign data_mem_pkt_o[73] = lce_data_cmd_i[79];
  assign data_mem_pkt_o[72] = lce_data_cmd_i[78];
  assign data_mem_pkt_o[71] = lce_data_cmd_i[77];
  assign data_mem_pkt_o[70] = lce_data_cmd_i[76];
  assign data_mem_pkt_o[69] = lce_data_cmd_i[75];
  assign data_mem_pkt_o[68] = lce_data_cmd_i[74];
  assign data_mem_pkt_o[67] = lce_data_cmd_i[73];
  assign data_mem_pkt_o[66] = lce_data_cmd_i[72];
  assign data_mem_pkt_o[65] = lce_data_cmd_i[71];
  assign data_mem_pkt_o[64] = lce_data_cmd_i[70];
  assign data_mem_pkt_o[63] = lce_data_cmd_i[69];
  assign data_mem_pkt_o[62] = lce_data_cmd_i[68];
  assign data_mem_pkt_o[61] = lce_data_cmd_i[67];
  assign data_mem_pkt_o[60] = lce_data_cmd_i[66];
  assign data_mem_pkt_o[59] = lce_data_cmd_i[65];
  assign data_mem_pkt_o[58] = lce_data_cmd_i[64];
  assign data_mem_pkt_o[57] = lce_data_cmd_i[63];
  assign data_mem_pkt_o[56] = lce_data_cmd_i[62];
  assign data_mem_pkt_o[55] = lce_data_cmd_i[61];
  assign data_mem_pkt_o[54] = lce_data_cmd_i[60];
  assign data_mem_pkt_o[53] = lce_data_cmd_i[59];
  assign data_mem_pkt_o[52] = lce_data_cmd_i[58];
  assign data_mem_pkt_o[51] = lce_data_cmd_i[57];
  assign data_mem_pkt_o[50] = lce_data_cmd_i[56];
  assign data_mem_pkt_o[49] = lce_data_cmd_i[55];
  assign data_mem_pkt_o[48] = lce_data_cmd_i[54];
  assign data_mem_pkt_o[47] = lce_data_cmd_i[53];
  assign data_mem_pkt_o[46] = lce_data_cmd_i[52];
  assign data_mem_pkt_o[45] = lce_data_cmd_i[51];
  assign data_mem_pkt_o[44] = lce_data_cmd_i[50];
  assign data_mem_pkt_o[43] = lce_data_cmd_i[49];
  assign data_mem_pkt_o[42] = lce_data_cmd_i[48];
  assign data_mem_pkt_o[41] = lce_data_cmd_i[47];
  assign data_mem_pkt_o[40] = lce_data_cmd_i[46];
  assign data_mem_pkt_o[39] = lce_data_cmd_i[45];
  assign data_mem_pkt_o[38] = lce_data_cmd_i[44];
  assign data_mem_pkt_o[37] = lce_data_cmd_i[43];
  assign data_mem_pkt_o[36] = lce_data_cmd_i[42];
  assign data_mem_pkt_o[35] = lce_data_cmd_i[41];
  assign data_mem_pkt_o[34] = lce_data_cmd_i[40];
  assign data_mem_pkt_o[33] = lce_data_cmd_i[39];
  assign data_mem_pkt_o[32] = lce_data_cmd_i[38];
  assign data_mem_pkt_o[31] = lce_data_cmd_i[37];
  assign data_mem_pkt_o[30] = lce_data_cmd_i[36];
  assign data_mem_pkt_o[29] = lce_data_cmd_i[35];
  assign data_mem_pkt_o[28] = lce_data_cmd_i[34];
  assign data_mem_pkt_o[27] = lce_data_cmd_i[33];
  assign data_mem_pkt_o[26] = lce_data_cmd_i[32];
  assign data_mem_pkt_o[25] = lce_data_cmd_i[31];
  assign data_mem_pkt_o[24] = lce_data_cmd_i[30];
  assign data_mem_pkt_o[23] = lce_data_cmd_i[29];
  assign data_mem_pkt_o[22] = lce_data_cmd_i[28];
  assign data_mem_pkt_o[21] = lce_data_cmd_i[27];
  assign data_mem_pkt_o[20] = lce_data_cmd_i[26];
  assign data_mem_pkt_o[19] = lce_data_cmd_i[25];
  assign data_mem_pkt_o[18] = lce_data_cmd_i[24];
  assign data_mem_pkt_o[17] = lce_data_cmd_i[23];
  assign data_mem_pkt_o[16] = lce_data_cmd_i[22];
  assign data_mem_pkt_o[15] = lce_data_cmd_i[21];
  assign data_mem_pkt_o[14] = lce_data_cmd_i[20];
  assign data_mem_pkt_o[13] = lce_data_cmd_i[19];
  assign data_mem_pkt_o[12] = lce_data_cmd_i[18];
  assign data_mem_pkt_o[11] = lce_data_cmd_i[17];
  assign data_mem_pkt_o[10] = lce_data_cmd_i[16];
  assign data_mem_pkt_o[9] = lce_data_cmd_i[15];
  assign data_mem_pkt_o[8] = lce_data_cmd_i[14];
  assign data_mem_pkt_o[7] = lce_data_cmd_i[13];
  assign data_mem_pkt_o[6] = lce_data_cmd_i[12];
  assign data_mem_pkt_o[5] = lce_data_cmd_i[11];
  assign data_mem_pkt_o[4] = lce_data_cmd_i[10];
  assign data_mem_pkt_o[3] = lce_data_cmd_i[9];
  assign data_mem_pkt_o[2] = lce_data_cmd_i[8];
  assign data_mem_pkt_o[1] = lce_data_cmd_i[7];
  assign data_mem_pkt_o[0] = lce_data_cmd_i[6];
  assign lce_data_cmd_yumi_o = data_mem_pkt_yumi_i;
  assign data_mem_pkt_v_o = lce_data_cmd_v_i;
  assign data_mem_pkt_o[521] = miss_addr_i[11];
  assign data_mem_pkt_o[520] = miss_addr_i[10];
  assign data_mem_pkt_o[519] = miss_addr_i[9];
  assign data_mem_pkt_o[518] = miss_addr_i[8];
  assign data_mem_pkt_o[517] = miss_addr_i[7];
  assign data_mem_pkt_o[516] = miss_addr_i[6];
  assign N0 = ~lce_data_cmd_i[3];
  assign N1 = N0 | lce_data_cmd_i[4];
  assign N2 = ~N1;
  assign N3 = lce_data_cmd_i[3] | lce_data_cmd_i[4];
  assign N4 = ~N3;
  assign cce_data_received_o = data_mem_pkt_yumi_i & N2;
  assign tr_data_received_o = data_mem_pkt_yumi_i & N4;

endmodule



module bp_fe_lce_data_width_p64_paddr_width_p22_lce_data_width_p512_sets_p64_ways_p8_num_cce_p1_num_lce_p2
(
  clk_i,
  reset_i,
  id_i,
  ready_o,
  cache_miss_o,
  miss_i,
  miss_addr_i,
  data_mem_data_i,
  data_mem_pkt_o,
  data_mem_pkt_v_o,
  data_mem_pkt_yumi_i,
  tag_mem_pkt_o,
  tag_mem_pkt_v_o,
  tag_mem_pkt_yumi_i,
  metadata_mem_pkt_v_o,
  metadata_mem_pkt_o,
  lru_way_i,
  metadata_mem_pkt_yumi_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i
);

  input [0:0] id_i;
  input [21:0] miss_addr_i;
  input [511:0] data_mem_data_i;
  output [521:0] data_mem_pkt_o;
  output [22:0] tag_mem_pkt_o;
  output [9:0] metadata_mem_pkt_o;
  input [2:0] lru_way_i;
  output [96:0] lce_req_o;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  input [35:0] lce_cmd_i;
  input [517:0] lce_data_cmd_i;
  output [517:0] lce_data_cmd_o;
  input clk_i;
  input reset_i;
  input miss_i;
  input data_mem_pkt_yumi_i;
  input tag_mem_pkt_yumi_i;
  input metadata_mem_pkt_yumi_i;
  input lce_req_ready_i;
  input lce_resp_ready_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_v_i;
  input lce_data_cmd_ready_i;
  output ready_o;
  output cache_miss_o;
  output data_mem_pkt_v_o;
  output tag_mem_pkt_v_o;
  output metadata_mem_pkt_v_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_ready_o;
  output lce_data_cmd_ready_o;
  output lce_data_cmd_v_o;
  wire [521:0] data_mem_pkt_o,lce_cmd_data_mem_pkt_lo,lce_data_cmd_data_mem_pkt_lo;
  wire [22:0] tag_mem_pkt_o;
  wire [9:0] metadata_mem_pkt_o;
  wire [96:0] lce_req_o;
  wire [25:0] lce_resp_o,lce_req_lce_resp_lo,lce_cmd_lce_resp_lo;
  wire [536:0] lce_data_resp_o;
  wire [517:0] lce_data_cmd_o;
  wire ready_o,cache_miss_o,data_mem_pkt_v_o,tag_mem_pkt_v_o,metadata_mem_pkt_v_o,
  lce_req_v_o,lce_resp_v_o,lce_data_resp_v_o,lce_cmd_ready_o,lce_data_cmd_ready_o,
  lce_data_cmd_v_o,N0,N1,N2,N3,tr_data_received,cce_data_received,set_tag_received,
  set_tag_wakeup_received,lce_req_lce_resp_v_lo,lce_req_lce_resp_yumi_li,lce_ready_lo,
  lce_cmd_data_mem_pkt_v_lo,lce_cmd_data_mem_pkt_yumi_li,lce_cmd_lce_resp_v_lo,
  lce_cmd_lce_resp_yumi_li,lce_data_cmd_data_mem_pkt_v_lo,
  lce_data_cmd_data_mem_pkt_yumi_li,N4,N5,N6,N7,N8,N9;
  wire [21:0] miss_addr_lo;

  bp_fe_lce_req_data_width_p64_paddr_width_p22_num_cce_p1_num_lce_p2_sets_p64_ways_p8
  lce_req_inst
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .id_i(id_i[0]),
    .miss_i(miss_i),
    .miss_addr_i(miss_addr_i),
    .lru_way_i(lru_way_i),
    .cache_miss_o(cache_miss_o),
    .miss_addr_o(miss_addr_lo),
    .tr_data_received_i(tr_data_received),
    .cce_data_received_i(cce_data_received),
    .set_tag_received_i(set_tag_received),
    .set_tag_wakeup_received_i(set_tag_wakeup_received),
    .lce_req_o(lce_req_o),
    .lce_req_v_o(lce_req_v_o),
    .lce_req_ready_i(lce_req_ready_i),
    .lce_resp_o(lce_req_lce_resp_lo),
    .lce_resp_v_o(lce_req_lce_resp_v_lo),
    .lce_resp_yumi_i(lce_req_lce_resp_yumi_li)
  );


  bp_fe_lce_cmd_data_width_p64_paddr_width_p22_lce_data_width_p512_sets_p64_ways_p8_num_cce_p1_num_lce_p2
  lce_cmd_inst
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .id_i(id_i[0]),
    .lce_ready_o(lce_ready_lo),
    .set_tag_received_o(set_tag_received),
    .set_tag_wakeup_received_o(set_tag_wakeup_received),
    .data_mem_data_i(data_mem_data_i),
    .data_mem_pkt_o(lce_cmd_data_mem_pkt_lo),
    .data_mem_pkt_v_o(lce_cmd_data_mem_pkt_v_lo),
    .data_mem_pkt_yumi_i(lce_cmd_data_mem_pkt_yumi_li),
    .tag_mem_pkt_o(tag_mem_pkt_o),
    .tag_mem_pkt_v_o(tag_mem_pkt_v_o),
    .tag_mem_pkt_yumi_i(tag_mem_pkt_yumi_i),
    .metadata_mem_pkt_v_o(metadata_mem_pkt_v_o),
    .metadata_mem_pkt_o(metadata_mem_pkt_o),
    .metadata_mem_pkt_yumi_i(metadata_mem_pkt_yumi_i),
    .lce_resp_o(lce_cmd_lce_resp_lo),
    .lce_resp_v_o(lce_cmd_lce_resp_v_lo),
    .lce_resp_yumi_i(lce_cmd_lce_resp_yumi_li),
    .lce_data_resp_o(lce_data_resp_o),
    .lce_data_resp_v_o(lce_data_resp_v_o),
    .lce_data_resp_ready_i(lce_data_resp_ready_i),
    .lce_cmd_i(lce_cmd_i),
    .lce_cmd_v_i(lce_cmd_v_i),
    .lce_cmd_yumi_o(lce_cmd_ready_o),
    .lce_data_cmd_o(lce_data_cmd_o),
    .lce_data_cmd_v_o(lce_data_cmd_v_o),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_i)
  );


  bp_fe_lce_data_cmd_data_width_p64_paddr_width_p22_lce_data_width_p512_num_cce_p1_num_lce_p2_sets_p64_ways_p8
  lce_data_cmd
  (
    .cce_data_received_o(cce_data_received),
    .tr_data_received_o(tr_data_received),
    .miss_addr_i(miss_addr_lo),
    .lce_data_cmd_i(lce_data_cmd_i),
    .lce_data_cmd_v_i(lce_data_cmd_v_i),
    .lce_data_cmd_yumi_o(lce_data_cmd_ready_o),
    .data_mem_pkt_v_o(lce_data_cmd_data_mem_pkt_v_lo),
    .data_mem_pkt_o(lce_data_cmd_data_mem_pkt_lo),
    .data_mem_pkt_yumi_i(lce_data_cmd_data_mem_pkt_yumi_li)
  );

  assign data_mem_pkt_v_o = (N0)? 1'b1 :
                            (N1)? lce_cmd_data_mem_pkt_v_lo : 1'b0;
  assign N0 = lce_data_cmd_data_mem_pkt_v_lo;
  assign N1 = N4;
  assign data_mem_pkt_o = (N0)? lce_data_cmd_data_mem_pkt_lo :
                          (N1)? lce_cmd_data_mem_pkt_lo : 1'b0;
  assign lce_data_cmd_data_mem_pkt_yumi_li = (N0)? data_mem_pkt_yumi_i :
                                             (N1)? 1'b0 : 1'b0;
  assign lce_cmd_data_mem_pkt_yumi_li = (N0)? 1'b0 :
                                        (N1)? data_mem_pkt_yumi_i : 1'b0;
  assign lce_resp_v_o = (N2)? 1'b1 :
                        (N3)? lce_cmd_lce_resp_v_lo : 1'b0;
  assign N2 = lce_req_lce_resp_v_lo;
  assign N3 = N5;
  assign lce_resp_o = (N2)? lce_req_lce_resp_lo :
                      (N3)? lce_cmd_lce_resp_lo : 1'b0;
  assign lce_req_lce_resp_yumi_li = (N2)? lce_resp_ready_i :
                                    (N3)? 1'b0 : 1'b0;
  assign lce_cmd_lce_resp_yumi_li = (N2)? 1'b0 :
                                    (N3)? N6 : 1'b0;
  assign N4 = ~lce_data_cmd_data_mem_pkt_v_lo;
  assign N5 = ~lce_req_lce_resp_v_lo;
  assign N6 = lce_cmd_lce_resp_v_lo & lce_resp_ready_i;
  assign ready_o = N8 & N9;
  assign N8 = lce_ready_lo & N7;
  assign N7 = ~1'b0;
  assign N9 = ~cache_miss_o;

endmodule



module bsg_mux_width_p64_els_p8
(
  data_i,
  sel_i,
  data_o
);

  input [511:0] data_i;
  input [2:0] sel_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;
  assign data_o[63] = (N7)? data_i[63] :
                      (N9)? data_i[127] :
                      (N11)? data_i[191] :
                      (N13)? data_i[255] :
                      (N8)? data_i[319] :
                      (N10)? data_i[383] :
                      (N12)? data_i[447] :
                      (N14)? data_i[511] : 1'b0;
  assign data_o[62] = (N7)? data_i[62] :
                      (N9)? data_i[126] :
                      (N11)? data_i[190] :
                      (N13)? data_i[254] :
                      (N8)? data_i[318] :
                      (N10)? data_i[382] :
                      (N12)? data_i[446] :
                      (N14)? data_i[510] : 1'b0;
  assign data_o[61] = (N7)? data_i[61] :
                      (N9)? data_i[125] :
                      (N11)? data_i[189] :
                      (N13)? data_i[253] :
                      (N8)? data_i[317] :
                      (N10)? data_i[381] :
                      (N12)? data_i[445] :
                      (N14)? data_i[509] : 1'b0;
  assign data_o[60] = (N7)? data_i[60] :
                      (N9)? data_i[124] :
                      (N11)? data_i[188] :
                      (N13)? data_i[252] :
                      (N8)? data_i[316] :
                      (N10)? data_i[380] :
                      (N12)? data_i[444] :
                      (N14)? data_i[508] : 1'b0;
  assign data_o[59] = (N7)? data_i[59] :
                      (N9)? data_i[123] :
                      (N11)? data_i[187] :
                      (N13)? data_i[251] :
                      (N8)? data_i[315] :
                      (N10)? data_i[379] :
                      (N12)? data_i[443] :
                      (N14)? data_i[507] : 1'b0;
  assign data_o[58] = (N7)? data_i[58] :
                      (N9)? data_i[122] :
                      (N11)? data_i[186] :
                      (N13)? data_i[250] :
                      (N8)? data_i[314] :
                      (N10)? data_i[378] :
                      (N12)? data_i[442] :
                      (N14)? data_i[506] : 1'b0;
  assign data_o[57] = (N7)? data_i[57] :
                      (N9)? data_i[121] :
                      (N11)? data_i[185] :
                      (N13)? data_i[249] :
                      (N8)? data_i[313] :
                      (N10)? data_i[377] :
                      (N12)? data_i[441] :
                      (N14)? data_i[505] : 1'b0;
  assign data_o[56] = (N7)? data_i[56] :
                      (N9)? data_i[120] :
                      (N11)? data_i[184] :
                      (N13)? data_i[248] :
                      (N8)? data_i[312] :
                      (N10)? data_i[376] :
                      (N12)? data_i[440] :
                      (N14)? data_i[504] : 1'b0;
  assign data_o[55] = (N7)? data_i[55] :
                      (N9)? data_i[119] :
                      (N11)? data_i[183] :
                      (N13)? data_i[247] :
                      (N8)? data_i[311] :
                      (N10)? data_i[375] :
                      (N12)? data_i[439] :
                      (N14)? data_i[503] : 1'b0;
  assign data_o[54] = (N7)? data_i[54] :
                      (N9)? data_i[118] :
                      (N11)? data_i[182] :
                      (N13)? data_i[246] :
                      (N8)? data_i[310] :
                      (N10)? data_i[374] :
                      (N12)? data_i[438] :
                      (N14)? data_i[502] : 1'b0;
  assign data_o[53] = (N7)? data_i[53] :
                      (N9)? data_i[117] :
                      (N11)? data_i[181] :
                      (N13)? data_i[245] :
                      (N8)? data_i[309] :
                      (N10)? data_i[373] :
                      (N12)? data_i[437] :
                      (N14)? data_i[501] : 1'b0;
  assign data_o[52] = (N7)? data_i[52] :
                      (N9)? data_i[116] :
                      (N11)? data_i[180] :
                      (N13)? data_i[244] :
                      (N8)? data_i[308] :
                      (N10)? data_i[372] :
                      (N12)? data_i[436] :
                      (N14)? data_i[500] : 1'b0;
  assign data_o[51] = (N7)? data_i[51] :
                      (N9)? data_i[115] :
                      (N11)? data_i[179] :
                      (N13)? data_i[243] :
                      (N8)? data_i[307] :
                      (N10)? data_i[371] :
                      (N12)? data_i[435] :
                      (N14)? data_i[499] : 1'b0;
  assign data_o[50] = (N7)? data_i[50] :
                      (N9)? data_i[114] :
                      (N11)? data_i[178] :
                      (N13)? data_i[242] :
                      (N8)? data_i[306] :
                      (N10)? data_i[370] :
                      (N12)? data_i[434] :
                      (N14)? data_i[498] : 1'b0;
  assign data_o[49] = (N7)? data_i[49] :
                      (N9)? data_i[113] :
                      (N11)? data_i[177] :
                      (N13)? data_i[241] :
                      (N8)? data_i[305] :
                      (N10)? data_i[369] :
                      (N12)? data_i[433] :
                      (N14)? data_i[497] : 1'b0;
  assign data_o[48] = (N7)? data_i[48] :
                      (N9)? data_i[112] :
                      (N11)? data_i[176] :
                      (N13)? data_i[240] :
                      (N8)? data_i[304] :
                      (N10)? data_i[368] :
                      (N12)? data_i[432] :
                      (N14)? data_i[496] : 1'b0;
  assign data_o[47] = (N7)? data_i[47] :
                      (N9)? data_i[111] :
                      (N11)? data_i[175] :
                      (N13)? data_i[239] :
                      (N8)? data_i[303] :
                      (N10)? data_i[367] :
                      (N12)? data_i[431] :
                      (N14)? data_i[495] : 1'b0;
  assign data_o[46] = (N7)? data_i[46] :
                      (N9)? data_i[110] :
                      (N11)? data_i[174] :
                      (N13)? data_i[238] :
                      (N8)? data_i[302] :
                      (N10)? data_i[366] :
                      (N12)? data_i[430] :
                      (N14)? data_i[494] : 1'b0;
  assign data_o[45] = (N7)? data_i[45] :
                      (N9)? data_i[109] :
                      (N11)? data_i[173] :
                      (N13)? data_i[237] :
                      (N8)? data_i[301] :
                      (N10)? data_i[365] :
                      (N12)? data_i[429] :
                      (N14)? data_i[493] : 1'b0;
  assign data_o[44] = (N7)? data_i[44] :
                      (N9)? data_i[108] :
                      (N11)? data_i[172] :
                      (N13)? data_i[236] :
                      (N8)? data_i[300] :
                      (N10)? data_i[364] :
                      (N12)? data_i[428] :
                      (N14)? data_i[492] : 1'b0;
  assign data_o[43] = (N7)? data_i[43] :
                      (N9)? data_i[107] :
                      (N11)? data_i[171] :
                      (N13)? data_i[235] :
                      (N8)? data_i[299] :
                      (N10)? data_i[363] :
                      (N12)? data_i[427] :
                      (N14)? data_i[491] : 1'b0;
  assign data_o[42] = (N7)? data_i[42] :
                      (N9)? data_i[106] :
                      (N11)? data_i[170] :
                      (N13)? data_i[234] :
                      (N8)? data_i[298] :
                      (N10)? data_i[362] :
                      (N12)? data_i[426] :
                      (N14)? data_i[490] : 1'b0;
  assign data_o[41] = (N7)? data_i[41] :
                      (N9)? data_i[105] :
                      (N11)? data_i[169] :
                      (N13)? data_i[233] :
                      (N8)? data_i[297] :
                      (N10)? data_i[361] :
                      (N12)? data_i[425] :
                      (N14)? data_i[489] : 1'b0;
  assign data_o[40] = (N7)? data_i[40] :
                      (N9)? data_i[104] :
                      (N11)? data_i[168] :
                      (N13)? data_i[232] :
                      (N8)? data_i[296] :
                      (N10)? data_i[360] :
                      (N12)? data_i[424] :
                      (N14)? data_i[488] : 1'b0;
  assign data_o[39] = (N7)? data_i[39] :
                      (N9)? data_i[103] :
                      (N11)? data_i[167] :
                      (N13)? data_i[231] :
                      (N8)? data_i[295] :
                      (N10)? data_i[359] :
                      (N12)? data_i[423] :
                      (N14)? data_i[487] : 1'b0;
  assign data_o[38] = (N7)? data_i[38] :
                      (N9)? data_i[102] :
                      (N11)? data_i[166] :
                      (N13)? data_i[230] :
                      (N8)? data_i[294] :
                      (N10)? data_i[358] :
                      (N12)? data_i[422] :
                      (N14)? data_i[486] : 1'b0;
  assign data_o[37] = (N7)? data_i[37] :
                      (N9)? data_i[101] :
                      (N11)? data_i[165] :
                      (N13)? data_i[229] :
                      (N8)? data_i[293] :
                      (N10)? data_i[357] :
                      (N12)? data_i[421] :
                      (N14)? data_i[485] : 1'b0;
  assign data_o[36] = (N7)? data_i[36] :
                      (N9)? data_i[100] :
                      (N11)? data_i[164] :
                      (N13)? data_i[228] :
                      (N8)? data_i[292] :
                      (N10)? data_i[356] :
                      (N12)? data_i[420] :
                      (N14)? data_i[484] : 1'b0;
  assign data_o[35] = (N7)? data_i[35] :
                      (N9)? data_i[99] :
                      (N11)? data_i[163] :
                      (N13)? data_i[227] :
                      (N8)? data_i[291] :
                      (N10)? data_i[355] :
                      (N12)? data_i[419] :
                      (N14)? data_i[483] : 1'b0;
  assign data_o[34] = (N7)? data_i[34] :
                      (N9)? data_i[98] :
                      (N11)? data_i[162] :
                      (N13)? data_i[226] :
                      (N8)? data_i[290] :
                      (N10)? data_i[354] :
                      (N12)? data_i[418] :
                      (N14)? data_i[482] : 1'b0;
  assign data_o[33] = (N7)? data_i[33] :
                      (N9)? data_i[97] :
                      (N11)? data_i[161] :
                      (N13)? data_i[225] :
                      (N8)? data_i[289] :
                      (N10)? data_i[353] :
                      (N12)? data_i[417] :
                      (N14)? data_i[481] : 1'b0;
  assign data_o[32] = (N7)? data_i[32] :
                      (N9)? data_i[96] :
                      (N11)? data_i[160] :
                      (N13)? data_i[224] :
                      (N8)? data_i[288] :
                      (N10)? data_i[352] :
                      (N12)? data_i[416] :
                      (N14)? data_i[480] : 1'b0;
  assign data_o[31] = (N7)? data_i[31] :
                      (N9)? data_i[95] :
                      (N11)? data_i[159] :
                      (N13)? data_i[223] :
                      (N8)? data_i[287] :
                      (N10)? data_i[351] :
                      (N12)? data_i[415] :
                      (N14)? data_i[479] : 1'b0;
  assign data_o[30] = (N7)? data_i[30] :
                      (N9)? data_i[94] :
                      (N11)? data_i[158] :
                      (N13)? data_i[222] :
                      (N8)? data_i[286] :
                      (N10)? data_i[350] :
                      (N12)? data_i[414] :
                      (N14)? data_i[478] : 1'b0;
  assign data_o[29] = (N7)? data_i[29] :
                      (N9)? data_i[93] :
                      (N11)? data_i[157] :
                      (N13)? data_i[221] :
                      (N8)? data_i[285] :
                      (N10)? data_i[349] :
                      (N12)? data_i[413] :
                      (N14)? data_i[477] : 1'b0;
  assign data_o[28] = (N7)? data_i[28] :
                      (N9)? data_i[92] :
                      (N11)? data_i[156] :
                      (N13)? data_i[220] :
                      (N8)? data_i[284] :
                      (N10)? data_i[348] :
                      (N12)? data_i[412] :
                      (N14)? data_i[476] : 1'b0;
  assign data_o[27] = (N7)? data_i[27] :
                      (N9)? data_i[91] :
                      (N11)? data_i[155] :
                      (N13)? data_i[219] :
                      (N8)? data_i[283] :
                      (N10)? data_i[347] :
                      (N12)? data_i[411] :
                      (N14)? data_i[475] : 1'b0;
  assign data_o[26] = (N7)? data_i[26] :
                      (N9)? data_i[90] :
                      (N11)? data_i[154] :
                      (N13)? data_i[218] :
                      (N8)? data_i[282] :
                      (N10)? data_i[346] :
                      (N12)? data_i[410] :
                      (N14)? data_i[474] : 1'b0;
  assign data_o[25] = (N7)? data_i[25] :
                      (N9)? data_i[89] :
                      (N11)? data_i[153] :
                      (N13)? data_i[217] :
                      (N8)? data_i[281] :
                      (N10)? data_i[345] :
                      (N12)? data_i[409] :
                      (N14)? data_i[473] : 1'b0;
  assign data_o[24] = (N7)? data_i[24] :
                      (N9)? data_i[88] :
                      (N11)? data_i[152] :
                      (N13)? data_i[216] :
                      (N8)? data_i[280] :
                      (N10)? data_i[344] :
                      (N12)? data_i[408] :
                      (N14)? data_i[472] : 1'b0;
  assign data_o[23] = (N7)? data_i[23] :
                      (N9)? data_i[87] :
                      (N11)? data_i[151] :
                      (N13)? data_i[215] :
                      (N8)? data_i[279] :
                      (N10)? data_i[343] :
                      (N12)? data_i[407] :
                      (N14)? data_i[471] : 1'b0;
  assign data_o[22] = (N7)? data_i[22] :
                      (N9)? data_i[86] :
                      (N11)? data_i[150] :
                      (N13)? data_i[214] :
                      (N8)? data_i[278] :
                      (N10)? data_i[342] :
                      (N12)? data_i[406] :
                      (N14)? data_i[470] : 1'b0;
  assign data_o[21] = (N7)? data_i[21] :
                      (N9)? data_i[85] :
                      (N11)? data_i[149] :
                      (N13)? data_i[213] :
                      (N8)? data_i[277] :
                      (N10)? data_i[341] :
                      (N12)? data_i[405] :
                      (N14)? data_i[469] : 1'b0;
  assign data_o[20] = (N7)? data_i[20] :
                      (N9)? data_i[84] :
                      (N11)? data_i[148] :
                      (N13)? data_i[212] :
                      (N8)? data_i[276] :
                      (N10)? data_i[340] :
                      (N12)? data_i[404] :
                      (N14)? data_i[468] : 1'b0;
  assign data_o[19] = (N7)? data_i[19] :
                      (N9)? data_i[83] :
                      (N11)? data_i[147] :
                      (N13)? data_i[211] :
                      (N8)? data_i[275] :
                      (N10)? data_i[339] :
                      (N12)? data_i[403] :
                      (N14)? data_i[467] : 1'b0;
  assign data_o[18] = (N7)? data_i[18] :
                      (N9)? data_i[82] :
                      (N11)? data_i[146] :
                      (N13)? data_i[210] :
                      (N8)? data_i[274] :
                      (N10)? data_i[338] :
                      (N12)? data_i[402] :
                      (N14)? data_i[466] : 1'b0;
  assign data_o[17] = (N7)? data_i[17] :
                      (N9)? data_i[81] :
                      (N11)? data_i[145] :
                      (N13)? data_i[209] :
                      (N8)? data_i[273] :
                      (N10)? data_i[337] :
                      (N12)? data_i[401] :
                      (N14)? data_i[465] : 1'b0;
  assign data_o[16] = (N7)? data_i[16] :
                      (N9)? data_i[80] :
                      (N11)? data_i[144] :
                      (N13)? data_i[208] :
                      (N8)? data_i[272] :
                      (N10)? data_i[336] :
                      (N12)? data_i[400] :
                      (N14)? data_i[464] : 1'b0;
  assign data_o[15] = (N7)? data_i[15] :
                      (N9)? data_i[79] :
                      (N11)? data_i[143] :
                      (N13)? data_i[207] :
                      (N8)? data_i[271] :
                      (N10)? data_i[335] :
                      (N12)? data_i[399] :
                      (N14)? data_i[463] : 1'b0;
  assign data_o[14] = (N7)? data_i[14] :
                      (N9)? data_i[78] :
                      (N11)? data_i[142] :
                      (N13)? data_i[206] :
                      (N8)? data_i[270] :
                      (N10)? data_i[334] :
                      (N12)? data_i[398] :
                      (N14)? data_i[462] : 1'b0;
  assign data_o[13] = (N7)? data_i[13] :
                      (N9)? data_i[77] :
                      (N11)? data_i[141] :
                      (N13)? data_i[205] :
                      (N8)? data_i[269] :
                      (N10)? data_i[333] :
                      (N12)? data_i[397] :
                      (N14)? data_i[461] : 1'b0;
  assign data_o[12] = (N7)? data_i[12] :
                      (N9)? data_i[76] :
                      (N11)? data_i[140] :
                      (N13)? data_i[204] :
                      (N8)? data_i[268] :
                      (N10)? data_i[332] :
                      (N12)? data_i[396] :
                      (N14)? data_i[460] : 1'b0;
  assign data_o[11] = (N7)? data_i[11] :
                      (N9)? data_i[75] :
                      (N11)? data_i[139] :
                      (N13)? data_i[203] :
                      (N8)? data_i[267] :
                      (N10)? data_i[331] :
                      (N12)? data_i[395] :
                      (N14)? data_i[459] : 1'b0;
  assign data_o[10] = (N7)? data_i[10] :
                      (N9)? data_i[74] :
                      (N11)? data_i[138] :
                      (N13)? data_i[202] :
                      (N8)? data_i[266] :
                      (N10)? data_i[330] :
                      (N12)? data_i[394] :
                      (N14)? data_i[458] : 1'b0;
  assign data_o[9] = (N7)? data_i[9] :
                     (N9)? data_i[73] :
                     (N11)? data_i[137] :
                     (N13)? data_i[201] :
                     (N8)? data_i[265] :
                     (N10)? data_i[329] :
                     (N12)? data_i[393] :
                     (N14)? data_i[457] : 1'b0;
  assign data_o[8] = (N7)? data_i[8] :
                     (N9)? data_i[72] :
                     (N11)? data_i[136] :
                     (N13)? data_i[200] :
                     (N8)? data_i[264] :
                     (N10)? data_i[328] :
                     (N12)? data_i[392] :
                     (N14)? data_i[456] : 1'b0;
  assign data_o[7] = (N7)? data_i[7] :
                     (N9)? data_i[71] :
                     (N11)? data_i[135] :
                     (N13)? data_i[199] :
                     (N8)? data_i[263] :
                     (N10)? data_i[327] :
                     (N12)? data_i[391] :
                     (N14)? data_i[455] : 1'b0;
  assign data_o[6] = (N7)? data_i[6] :
                     (N9)? data_i[70] :
                     (N11)? data_i[134] :
                     (N13)? data_i[198] :
                     (N8)? data_i[262] :
                     (N10)? data_i[326] :
                     (N12)? data_i[390] :
                     (N14)? data_i[454] : 1'b0;
  assign data_o[5] = (N7)? data_i[5] :
                     (N9)? data_i[69] :
                     (N11)? data_i[133] :
                     (N13)? data_i[197] :
                     (N8)? data_i[261] :
                     (N10)? data_i[325] :
                     (N12)? data_i[389] :
                     (N14)? data_i[453] : 1'b0;
  assign data_o[4] = (N7)? data_i[4] :
                     (N9)? data_i[68] :
                     (N11)? data_i[132] :
                     (N13)? data_i[196] :
                     (N8)? data_i[260] :
                     (N10)? data_i[324] :
                     (N12)? data_i[388] :
                     (N14)? data_i[452] : 1'b0;
  assign data_o[3] = (N7)? data_i[3] :
                     (N9)? data_i[67] :
                     (N11)? data_i[131] :
                     (N13)? data_i[195] :
                     (N8)? data_i[259] :
                     (N10)? data_i[323] :
                     (N12)? data_i[387] :
                     (N14)? data_i[451] : 1'b0;
  assign data_o[2] = (N7)? data_i[2] :
                     (N9)? data_i[66] :
                     (N11)? data_i[130] :
                     (N13)? data_i[194] :
                     (N8)? data_i[258] :
                     (N10)? data_i[322] :
                     (N12)? data_i[386] :
                     (N14)? data_i[450] : 1'b0;
  assign data_o[1] = (N7)? data_i[1] :
                     (N9)? data_i[65] :
                     (N11)? data_i[129] :
                     (N13)? data_i[193] :
                     (N8)? data_i[257] :
                     (N10)? data_i[321] :
                     (N12)? data_i[385] :
                     (N14)? data_i[449] : 1'b0;
  assign data_o[0] = (N7)? data_i[0] :
                     (N9)? data_i[64] :
                     (N11)? data_i[128] :
                     (N13)? data_i[192] :
                     (N8)? data_i[256] :
                     (N10)? data_i[320] :
                     (N12)? data_i[384] :
                     (N14)? data_i[448] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];
  assign N6 = ~sel_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & sel_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & sel_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & sel_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & sel_i[2];

endmodule



module bsg_swap_width_p64
(
  data_i,
  swap_i,
  data_o
);

  input [127:0] data_i;
  output [127:0] data_o;
  input swap_i;
  wire [127:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[63:0], data_i[127:64] } :
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p128
(
  data_i,
  swap_i,
  data_o
);

  input [255:0] data_i;
  output [255:0] data_o;
  input swap_i;
  wire [255:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[127:0], data_i[255:128] } :
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p256
(
  data_i,
  swap_i,
  data_o
);

  input [511:0] data_i;
  output [511:0] data_o;
  input swap_i;
  wire [511:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[255:0], data_i[511:256] } :
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_mux_butterfly_width_p64_els_p8
(
  data_i,
  sel_i,
  data_o
);

  input [511:0] data_i;
  input [2:0] sel_i;
  output [511:0] data_o;
  wire [511:0] data_o;
  wire data_stage_1__511_,data_stage_1__510_,data_stage_1__509_,data_stage_1__508_,
  data_stage_1__507_,data_stage_1__506_,data_stage_1__505_,data_stage_1__504_,
  data_stage_1__503_,data_stage_1__502_,data_stage_1__501_,data_stage_1__500_,
  data_stage_1__499_,data_stage_1__498_,data_stage_1__497_,data_stage_1__496_,
  data_stage_1__495_,data_stage_1__494_,data_stage_1__493_,data_stage_1__492_,data_stage_1__491_,
  data_stage_1__490_,data_stage_1__489_,data_stage_1__488_,data_stage_1__487_,
  data_stage_1__486_,data_stage_1__485_,data_stage_1__484_,data_stage_1__483_,
  data_stage_1__482_,data_stage_1__481_,data_stage_1__480_,data_stage_1__479_,
  data_stage_1__478_,data_stage_1__477_,data_stage_1__476_,data_stage_1__475_,
  data_stage_1__474_,data_stage_1__473_,data_stage_1__472_,data_stage_1__471_,data_stage_1__470_,
  data_stage_1__469_,data_stage_1__468_,data_stage_1__467_,data_stage_1__466_,
  data_stage_1__465_,data_stage_1__464_,data_stage_1__463_,data_stage_1__462_,
  data_stage_1__461_,data_stage_1__460_,data_stage_1__459_,data_stage_1__458_,
  data_stage_1__457_,data_stage_1__456_,data_stage_1__455_,data_stage_1__454_,
  data_stage_1__453_,data_stage_1__452_,data_stage_1__451_,data_stage_1__450_,data_stage_1__449_,
  data_stage_1__448_,data_stage_1__447_,data_stage_1__446_,data_stage_1__445_,
  data_stage_1__444_,data_stage_1__443_,data_stage_1__442_,data_stage_1__441_,
  data_stage_1__440_,data_stage_1__439_,data_stage_1__438_,data_stage_1__437_,
  data_stage_1__436_,data_stage_1__435_,data_stage_1__434_,data_stage_1__433_,data_stage_1__432_,
  data_stage_1__431_,data_stage_1__430_,data_stage_1__429_,data_stage_1__428_,
  data_stage_1__427_,data_stage_1__426_,data_stage_1__425_,data_stage_1__424_,
  data_stage_1__423_,data_stage_1__422_,data_stage_1__421_,data_stage_1__420_,
  data_stage_1__419_,data_stage_1__418_,data_stage_1__417_,data_stage_1__416_,
  data_stage_1__415_,data_stage_1__414_,data_stage_1__413_,data_stage_1__412_,data_stage_1__411_,
  data_stage_1__410_,data_stage_1__409_,data_stage_1__408_,data_stage_1__407_,
  data_stage_1__406_,data_stage_1__405_,data_stage_1__404_,data_stage_1__403_,
  data_stage_1__402_,data_stage_1__401_,data_stage_1__400_,data_stage_1__399_,
  data_stage_1__398_,data_stage_1__397_,data_stage_1__396_,data_stage_1__395_,
  data_stage_1__394_,data_stage_1__393_,data_stage_1__392_,data_stage_1__391_,data_stage_1__390_,
  data_stage_1__389_,data_stage_1__388_,data_stage_1__387_,data_stage_1__386_,
  data_stage_1__385_,data_stage_1__384_,data_stage_1__383_,data_stage_1__382_,
  data_stage_1__381_,data_stage_1__380_,data_stage_1__379_,data_stage_1__378_,
  data_stage_1__377_,data_stage_1__376_,data_stage_1__375_,data_stage_1__374_,
  data_stage_1__373_,data_stage_1__372_,data_stage_1__371_,data_stage_1__370_,data_stage_1__369_,
  data_stage_1__368_,data_stage_1__367_,data_stage_1__366_,data_stage_1__365_,
  data_stage_1__364_,data_stage_1__363_,data_stage_1__362_,data_stage_1__361_,
  data_stage_1__360_,data_stage_1__359_,data_stage_1__358_,data_stage_1__357_,
  data_stage_1__356_,data_stage_1__355_,data_stage_1__354_,data_stage_1__353_,data_stage_1__352_,
  data_stage_1__351_,data_stage_1__350_,data_stage_1__349_,data_stage_1__348_,
  data_stage_1__347_,data_stage_1__346_,data_stage_1__345_,data_stage_1__344_,
  data_stage_1__343_,data_stage_1__342_,data_stage_1__341_,data_stage_1__340_,
  data_stage_1__339_,data_stage_1__338_,data_stage_1__337_,data_stage_1__336_,
  data_stage_1__335_,data_stage_1__334_,data_stage_1__333_,data_stage_1__332_,data_stage_1__331_,
  data_stage_1__330_,data_stage_1__329_,data_stage_1__328_,data_stage_1__327_,
  data_stage_1__326_,data_stage_1__325_,data_stage_1__324_,data_stage_1__323_,
  data_stage_1__322_,data_stage_1__321_,data_stage_1__320_,data_stage_1__319_,
  data_stage_1__318_,data_stage_1__317_,data_stage_1__316_,data_stage_1__315_,
  data_stage_1__314_,data_stage_1__313_,data_stage_1__312_,data_stage_1__311_,data_stage_1__310_,
  data_stage_1__309_,data_stage_1__308_,data_stage_1__307_,data_stage_1__306_,
  data_stage_1__305_,data_stage_1__304_,data_stage_1__303_,data_stage_1__302_,
  data_stage_1__301_,data_stage_1__300_,data_stage_1__299_,data_stage_1__298_,
  data_stage_1__297_,data_stage_1__296_,data_stage_1__295_,data_stage_1__294_,
  data_stage_1__293_,data_stage_1__292_,data_stage_1__291_,data_stage_1__290_,data_stage_1__289_,
  data_stage_1__288_,data_stage_1__287_,data_stage_1__286_,data_stage_1__285_,
  data_stage_1__284_,data_stage_1__283_,data_stage_1__282_,data_stage_1__281_,
  data_stage_1__280_,data_stage_1__279_,data_stage_1__278_,data_stage_1__277_,
  data_stage_1__276_,data_stage_1__275_,data_stage_1__274_,data_stage_1__273_,data_stage_1__272_,
  data_stage_1__271_,data_stage_1__270_,data_stage_1__269_,data_stage_1__268_,
  data_stage_1__267_,data_stage_1__266_,data_stage_1__265_,data_stage_1__264_,
  data_stage_1__263_,data_stage_1__262_,data_stage_1__261_,data_stage_1__260_,
  data_stage_1__259_,data_stage_1__258_,data_stage_1__257_,data_stage_1__256_,
  data_stage_1__255_,data_stage_1__254_,data_stage_1__253_,data_stage_1__252_,data_stage_1__251_,
  data_stage_1__250_,data_stage_1__249_,data_stage_1__248_,data_stage_1__247_,
  data_stage_1__246_,data_stage_1__245_,data_stage_1__244_,data_stage_1__243_,
  data_stage_1__242_,data_stage_1__241_,data_stage_1__240_,data_stage_1__239_,
  data_stage_1__238_,data_stage_1__237_,data_stage_1__236_,data_stage_1__235_,
  data_stage_1__234_,data_stage_1__233_,data_stage_1__232_,data_stage_1__231_,data_stage_1__230_,
  data_stage_1__229_,data_stage_1__228_,data_stage_1__227_,data_stage_1__226_,
  data_stage_1__225_,data_stage_1__224_,data_stage_1__223_,data_stage_1__222_,
  data_stage_1__221_,data_stage_1__220_,data_stage_1__219_,data_stage_1__218_,
  data_stage_1__217_,data_stage_1__216_,data_stage_1__215_,data_stage_1__214_,
  data_stage_1__213_,data_stage_1__212_,data_stage_1__211_,data_stage_1__210_,data_stage_1__209_,
  data_stage_1__208_,data_stage_1__207_,data_stage_1__206_,data_stage_1__205_,
  data_stage_1__204_,data_stage_1__203_,data_stage_1__202_,data_stage_1__201_,
  data_stage_1__200_,data_stage_1__199_,data_stage_1__198_,data_stage_1__197_,
  data_stage_1__196_,data_stage_1__195_,data_stage_1__194_,data_stage_1__193_,data_stage_1__192_,
  data_stage_1__191_,data_stage_1__190_,data_stage_1__189_,data_stage_1__188_,
  data_stage_1__187_,data_stage_1__186_,data_stage_1__185_,data_stage_1__184_,
  data_stage_1__183_,data_stage_1__182_,data_stage_1__181_,data_stage_1__180_,
  data_stage_1__179_,data_stage_1__178_,data_stage_1__177_,data_stage_1__176_,
  data_stage_1__175_,data_stage_1__174_,data_stage_1__173_,data_stage_1__172_,data_stage_1__171_,
  data_stage_1__170_,data_stage_1__169_,data_stage_1__168_,data_stage_1__167_,
  data_stage_1__166_,data_stage_1__165_,data_stage_1__164_,data_stage_1__163_,
  data_stage_1__162_,data_stage_1__161_,data_stage_1__160_,data_stage_1__159_,
  data_stage_1__158_,data_stage_1__157_,data_stage_1__156_,data_stage_1__155_,
  data_stage_1__154_,data_stage_1__153_,data_stage_1__152_,data_stage_1__151_,data_stage_1__150_,
  data_stage_1__149_,data_stage_1__148_,data_stage_1__147_,data_stage_1__146_,
  data_stage_1__145_,data_stage_1__144_,data_stage_1__143_,data_stage_1__142_,
  data_stage_1__141_,data_stage_1__140_,data_stage_1__139_,data_stage_1__138_,
  data_stage_1__137_,data_stage_1__136_,data_stage_1__135_,data_stage_1__134_,
  data_stage_1__133_,data_stage_1__132_,data_stage_1__131_,data_stage_1__130_,data_stage_1__129_,
  data_stage_1__128_,data_stage_1__127_,data_stage_1__126_,data_stage_1__125_,
  data_stage_1__124_,data_stage_1__123_,data_stage_1__122_,data_stage_1__121_,
  data_stage_1__120_,data_stage_1__119_,data_stage_1__118_,data_stage_1__117_,
  data_stage_1__116_,data_stage_1__115_,data_stage_1__114_,data_stage_1__113_,data_stage_1__112_,
  data_stage_1__111_,data_stage_1__110_,data_stage_1__109_,data_stage_1__108_,
  data_stage_1__107_,data_stage_1__106_,data_stage_1__105_,data_stage_1__104_,
  data_stage_1__103_,data_stage_1__102_,data_stage_1__101_,data_stage_1__100_,
  data_stage_1__99_,data_stage_1__98_,data_stage_1__97_,data_stage_1__96_,data_stage_1__95_,
  data_stage_1__94_,data_stage_1__93_,data_stage_1__92_,data_stage_1__91_,
  data_stage_1__90_,data_stage_1__89_,data_stage_1__88_,data_stage_1__87_,data_stage_1__86_,
  data_stage_1__85_,data_stage_1__84_,data_stage_1__83_,data_stage_1__82_,
  data_stage_1__81_,data_stage_1__80_,data_stage_1__79_,data_stage_1__78_,
  data_stage_1__77_,data_stage_1__76_,data_stage_1__75_,data_stage_1__74_,data_stage_1__73_,
  data_stage_1__72_,data_stage_1__71_,data_stage_1__70_,data_stage_1__69_,
  data_stage_1__68_,data_stage_1__67_,data_stage_1__66_,data_stage_1__65_,data_stage_1__64_,
  data_stage_1__63_,data_stage_1__62_,data_stage_1__61_,data_stage_1__60_,
  data_stage_1__59_,data_stage_1__58_,data_stage_1__57_,data_stage_1__56_,data_stage_1__55_,
  data_stage_1__54_,data_stage_1__53_,data_stage_1__52_,data_stage_1__51_,
  data_stage_1__50_,data_stage_1__49_,data_stage_1__48_,data_stage_1__47_,data_stage_1__46_,
  data_stage_1__45_,data_stage_1__44_,data_stage_1__43_,data_stage_1__42_,
  data_stage_1__41_,data_stage_1__40_,data_stage_1__39_,data_stage_1__38_,
  data_stage_1__37_,data_stage_1__36_,data_stage_1__35_,data_stage_1__34_,data_stage_1__33_,
  data_stage_1__32_,data_stage_1__31_,data_stage_1__30_,data_stage_1__29_,
  data_stage_1__28_,data_stage_1__27_,data_stage_1__26_,data_stage_1__25_,data_stage_1__24_,
  data_stage_1__23_,data_stage_1__22_,data_stage_1__21_,data_stage_1__20_,
  data_stage_1__19_,data_stage_1__18_,data_stage_1__17_,data_stage_1__16_,data_stage_1__15_,
  data_stage_1__14_,data_stage_1__13_,data_stage_1__12_,data_stage_1__11_,
  data_stage_1__10_,data_stage_1__9_,data_stage_1__8_,data_stage_1__7_,data_stage_1__6_,
  data_stage_1__5_,data_stage_1__4_,data_stage_1__3_,data_stage_1__2_,
  data_stage_1__1_,data_stage_1__0_,data_stage_2__511_,data_stage_2__510_,data_stage_2__509_,
  data_stage_2__508_,data_stage_2__507_,data_stage_2__506_,data_stage_2__505_,
  data_stage_2__504_,data_stage_2__503_,data_stage_2__502_,data_stage_2__501_,
  data_stage_2__500_,data_stage_2__499_,data_stage_2__498_,data_stage_2__497_,
  data_stage_2__496_,data_stage_2__495_,data_stage_2__494_,data_stage_2__493_,data_stage_2__492_,
  data_stage_2__491_,data_stage_2__490_,data_stage_2__489_,data_stage_2__488_,
  data_stage_2__487_,data_stage_2__486_,data_stage_2__485_,data_stage_2__484_,
  data_stage_2__483_,data_stage_2__482_,data_stage_2__481_,data_stage_2__480_,
  data_stage_2__479_,data_stage_2__478_,data_stage_2__477_,data_stage_2__476_,
  data_stage_2__475_,data_stage_2__474_,data_stage_2__473_,data_stage_2__472_,data_stage_2__471_,
  data_stage_2__470_,data_stage_2__469_,data_stage_2__468_,data_stage_2__467_,
  data_stage_2__466_,data_stage_2__465_,data_stage_2__464_,data_stage_2__463_,
  data_stage_2__462_,data_stage_2__461_,data_stage_2__460_,data_stage_2__459_,
  data_stage_2__458_,data_stage_2__457_,data_stage_2__456_,data_stage_2__455_,data_stage_2__454_,
  data_stage_2__453_,data_stage_2__452_,data_stage_2__451_,data_stage_2__450_,
  data_stage_2__449_,data_stage_2__448_,data_stage_2__447_,data_stage_2__446_,
  data_stage_2__445_,data_stage_2__444_,data_stage_2__443_,data_stage_2__442_,
  data_stage_2__441_,data_stage_2__440_,data_stage_2__439_,data_stage_2__438_,
  data_stage_2__437_,data_stage_2__436_,data_stage_2__435_,data_stage_2__434_,data_stage_2__433_,
  data_stage_2__432_,data_stage_2__431_,data_stage_2__430_,data_stage_2__429_,
  data_stage_2__428_,data_stage_2__427_,data_stage_2__426_,data_stage_2__425_,
  data_stage_2__424_,data_stage_2__423_,data_stage_2__422_,data_stage_2__421_,
  data_stage_2__420_,data_stage_2__419_,data_stage_2__418_,data_stage_2__417_,
  data_stage_2__416_,data_stage_2__415_,data_stage_2__414_,data_stage_2__413_,data_stage_2__412_,
  data_stage_2__411_,data_stage_2__410_,data_stage_2__409_,data_stage_2__408_,
  data_stage_2__407_,data_stage_2__406_,data_stage_2__405_,data_stage_2__404_,
  data_stage_2__403_,data_stage_2__402_,data_stage_2__401_,data_stage_2__400_,
  data_stage_2__399_,data_stage_2__398_,data_stage_2__397_,data_stage_2__396_,
  data_stage_2__395_,data_stage_2__394_,data_stage_2__393_,data_stage_2__392_,data_stage_2__391_,
  data_stage_2__390_,data_stage_2__389_,data_stage_2__388_,data_stage_2__387_,
  data_stage_2__386_,data_stage_2__385_,data_stage_2__384_,data_stage_2__383_,
  data_stage_2__382_,data_stage_2__381_,data_stage_2__380_,data_stage_2__379_,
  data_stage_2__378_,data_stage_2__377_,data_stage_2__376_,data_stage_2__375_,data_stage_2__374_,
  data_stage_2__373_,data_stage_2__372_,data_stage_2__371_,data_stage_2__370_,
  data_stage_2__369_,data_stage_2__368_,data_stage_2__367_,data_stage_2__366_,
  data_stage_2__365_,data_stage_2__364_,data_stage_2__363_,data_stage_2__362_,
  data_stage_2__361_,data_stage_2__360_,data_stage_2__359_,data_stage_2__358_,
  data_stage_2__357_,data_stage_2__356_,data_stage_2__355_,data_stage_2__354_,data_stage_2__353_,
  data_stage_2__352_,data_stage_2__351_,data_stage_2__350_,data_stage_2__349_,
  data_stage_2__348_,data_stage_2__347_,data_stage_2__346_,data_stage_2__345_,
  data_stage_2__344_,data_stage_2__343_,data_stage_2__342_,data_stage_2__341_,
  data_stage_2__340_,data_stage_2__339_,data_stage_2__338_,data_stage_2__337_,
  data_stage_2__336_,data_stage_2__335_,data_stage_2__334_,data_stage_2__333_,data_stage_2__332_,
  data_stage_2__331_,data_stage_2__330_,data_stage_2__329_,data_stage_2__328_,
  data_stage_2__327_,data_stage_2__326_,data_stage_2__325_,data_stage_2__324_,
  data_stage_2__323_,data_stage_2__322_,data_stage_2__321_,data_stage_2__320_,
  data_stage_2__319_,data_stage_2__318_,data_stage_2__317_,data_stage_2__316_,
  data_stage_2__315_,data_stage_2__314_,data_stage_2__313_,data_stage_2__312_,data_stage_2__311_,
  data_stage_2__310_,data_stage_2__309_,data_stage_2__308_,data_stage_2__307_,
  data_stage_2__306_,data_stage_2__305_,data_stage_2__304_,data_stage_2__303_,
  data_stage_2__302_,data_stage_2__301_,data_stage_2__300_,data_stage_2__299_,
  data_stage_2__298_,data_stage_2__297_,data_stage_2__296_,data_stage_2__295_,data_stage_2__294_,
  data_stage_2__293_,data_stage_2__292_,data_stage_2__291_,data_stage_2__290_,
  data_stage_2__289_,data_stage_2__288_,data_stage_2__287_,data_stage_2__286_,
  data_stage_2__285_,data_stage_2__284_,data_stage_2__283_,data_stage_2__282_,
  data_stage_2__281_,data_stage_2__280_,data_stage_2__279_,data_stage_2__278_,
  data_stage_2__277_,data_stage_2__276_,data_stage_2__275_,data_stage_2__274_,data_stage_2__273_,
  data_stage_2__272_,data_stage_2__271_,data_stage_2__270_,data_stage_2__269_,
  data_stage_2__268_,data_stage_2__267_,data_stage_2__266_,data_stage_2__265_,
  data_stage_2__264_,data_stage_2__263_,data_stage_2__262_,data_stage_2__261_,
  data_stage_2__260_,data_stage_2__259_,data_stage_2__258_,data_stage_2__257_,
  data_stage_2__256_,data_stage_2__255_,data_stage_2__254_,data_stage_2__253_,data_stage_2__252_,
  data_stage_2__251_,data_stage_2__250_,data_stage_2__249_,data_stage_2__248_,
  data_stage_2__247_,data_stage_2__246_,data_stage_2__245_,data_stage_2__244_,
  data_stage_2__243_,data_stage_2__242_,data_stage_2__241_,data_stage_2__240_,
  data_stage_2__239_,data_stage_2__238_,data_stage_2__237_,data_stage_2__236_,
  data_stage_2__235_,data_stage_2__234_,data_stage_2__233_,data_stage_2__232_,data_stage_2__231_,
  data_stage_2__230_,data_stage_2__229_,data_stage_2__228_,data_stage_2__227_,
  data_stage_2__226_,data_stage_2__225_,data_stage_2__224_,data_stage_2__223_,
  data_stage_2__222_,data_stage_2__221_,data_stage_2__220_,data_stage_2__219_,
  data_stage_2__218_,data_stage_2__217_,data_stage_2__216_,data_stage_2__215_,data_stage_2__214_,
  data_stage_2__213_,data_stage_2__212_,data_stage_2__211_,data_stage_2__210_,
  data_stage_2__209_,data_stage_2__208_,data_stage_2__207_,data_stage_2__206_,
  data_stage_2__205_,data_stage_2__204_,data_stage_2__203_,data_stage_2__202_,
  data_stage_2__201_,data_stage_2__200_,data_stage_2__199_,data_stage_2__198_,
  data_stage_2__197_,data_stage_2__196_,data_stage_2__195_,data_stage_2__194_,data_stage_2__193_,
  data_stage_2__192_,data_stage_2__191_,data_stage_2__190_,data_stage_2__189_,
  data_stage_2__188_,data_stage_2__187_,data_stage_2__186_,data_stage_2__185_,
  data_stage_2__184_,data_stage_2__183_,data_stage_2__182_,data_stage_2__181_,
  data_stage_2__180_,data_stage_2__179_,data_stage_2__178_,data_stage_2__177_,
  data_stage_2__176_,data_stage_2__175_,data_stage_2__174_,data_stage_2__173_,data_stage_2__172_,
  data_stage_2__171_,data_stage_2__170_,data_stage_2__169_,data_stage_2__168_,
  data_stage_2__167_,data_stage_2__166_,data_stage_2__165_,data_stage_2__164_,
  data_stage_2__163_,data_stage_2__162_,data_stage_2__161_,data_stage_2__160_,
  data_stage_2__159_,data_stage_2__158_,data_stage_2__157_,data_stage_2__156_,
  data_stage_2__155_,data_stage_2__154_,data_stage_2__153_,data_stage_2__152_,data_stage_2__151_,
  data_stage_2__150_,data_stage_2__149_,data_stage_2__148_,data_stage_2__147_,
  data_stage_2__146_,data_stage_2__145_,data_stage_2__144_,data_stage_2__143_,
  data_stage_2__142_,data_stage_2__141_,data_stage_2__140_,data_stage_2__139_,
  data_stage_2__138_,data_stage_2__137_,data_stage_2__136_,data_stage_2__135_,data_stage_2__134_,
  data_stage_2__133_,data_stage_2__132_,data_stage_2__131_,data_stage_2__130_,
  data_stage_2__129_,data_stage_2__128_,data_stage_2__127_,data_stage_2__126_,
  data_stage_2__125_,data_stage_2__124_,data_stage_2__123_,data_stage_2__122_,
  data_stage_2__121_,data_stage_2__120_,data_stage_2__119_,data_stage_2__118_,
  data_stage_2__117_,data_stage_2__116_,data_stage_2__115_,data_stage_2__114_,data_stage_2__113_,
  data_stage_2__112_,data_stage_2__111_,data_stage_2__110_,data_stage_2__109_,
  data_stage_2__108_,data_stage_2__107_,data_stage_2__106_,data_stage_2__105_,
  data_stage_2__104_,data_stage_2__103_,data_stage_2__102_,data_stage_2__101_,
  data_stage_2__100_,data_stage_2__99_,data_stage_2__98_,data_stage_2__97_,data_stage_2__96_,
  data_stage_2__95_,data_stage_2__94_,data_stage_2__93_,data_stage_2__92_,
  data_stage_2__91_,data_stage_2__90_,data_stage_2__89_,data_stage_2__88_,data_stage_2__87_,
  data_stage_2__86_,data_stage_2__85_,data_stage_2__84_,data_stage_2__83_,
  data_stage_2__82_,data_stage_2__81_,data_stage_2__80_,data_stage_2__79_,
  data_stage_2__78_,data_stage_2__77_,data_stage_2__76_,data_stage_2__75_,data_stage_2__74_,
  data_stage_2__73_,data_stage_2__72_,data_stage_2__71_,data_stage_2__70_,
  data_stage_2__69_,data_stage_2__68_,data_stage_2__67_,data_stage_2__66_,data_stage_2__65_,
  data_stage_2__64_,data_stage_2__63_,data_stage_2__62_,data_stage_2__61_,
  data_stage_2__60_,data_stage_2__59_,data_stage_2__58_,data_stage_2__57_,data_stage_2__56_,
  data_stage_2__55_,data_stage_2__54_,data_stage_2__53_,data_stage_2__52_,
  data_stage_2__51_,data_stage_2__50_,data_stage_2__49_,data_stage_2__48_,data_stage_2__47_,
  data_stage_2__46_,data_stage_2__45_,data_stage_2__44_,data_stage_2__43_,
  data_stage_2__42_,data_stage_2__41_,data_stage_2__40_,data_stage_2__39_,
  data_stage_2__38_,data_stage_2__37_,data_stage_2__36_,data_stage_2__35_,data_stage_2__34_,
  data_stage_2__33_,data_stage_2__32_,data_stage_2__31_,data_stage_2__30_,
  data_stage_2__29_,data_stage_2__28_,data_stage_2__27_,data_stage_2__26_,data_stage_2__25_,
  data_stage_2__24_,data_stage_2__23_,data_stage_2__22_,data_stage_2__21_,
  data_stage_2__20_,data_stage_2__19_,data_stage_2__18_,data_stage_2__17_,data_stage_2__16_,
  data_stage_2__15_,data_stage_2__14_,data_stage_2__13_,data_stage_2__12_,
  data_stage_2__11_,data_stage_2__10_,data_stage_2__9_,data_stage_2__8_,data_stage_2__7_,
  data_stage_2__6_,data_stage_2__5_,data_stage_2__4_,data_stage_2__3_,
  data_stage_2__2_,data_stage_2__1_,data_stage_2__0_;

  bsg_swap_width_p64
  mux_stage_0__mux_swap_0__swap_inst
  (
    .data_i(data_i[127:0]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__127_, data_stage_1__126_, data_stage_1__125_, data_stage_1__124_, data_stage_1__123_, data_stage_1__122_, data_stage_1__121_, data_stage_1__120_, data_stage_1__119_, data_stage_1__118_, data_stage_1__117_, data_stage_1__116_, data_stage_1__115_, data_stage_1__114_, data_stage_1__113_, data_stage_1__112_, data_stage_1__111_, data_stage_1__110_, data_stage_1__109_, data_stage_1__108_, data_stage_1__107_, data_stage_1__106_, data_stage_1__105_, data_stage_1__104_, data_stage_1__103_, data_stage_1__102_, data_stage_1__101_, data_stage_1__100_, data_stage_1__99_, data_stage_1__98_, data_stage_1__97_, data_stage_1__96_, data_stage_1__95_, data_stage_1__94_, data_stage_1__93_, data_stage_1__92_, data_stage_1__91_, data_stage_1__90_, data_stage_1__89_, data_stage_1__88_, data_stage_1__87_, data_stage_1__86_, data_stage_1__85_, data_stage_1__84_, data_stage_1__83_, data_stage_1__82_, data_stage_1__81_, data_stage_1__80_, data_stage_1__79_, data_stage_1__78_, data_stage_1__77_, data_stage_1__76_, data_stage_1__75_, data_stage_1__74_, data_stage_1__73_, data_stage_1__72_, data_stage_1__71_, data_stage_1__70_, data_stage_1__69_, data_stage_1__68_, data_stage_1__67_, data_stage_1__66_, data_stage_1__65_, data_stage_1__64_, data_stage_1__63_, data_stage_1__62_, data_stage_1__61_, data_stage_1__60_, data_stage_1__59_, data_stage_1__58_, data_stage_1__57_, data_stage_1__56_, data_stage_1__55_, data_stage_1__54_, data_stage_1__53_, data_stage_1__52_, data_stage_1__51_, data_stage_1__50_, data_stage_1__49_, data_stage_1__48_, data_stage_1__47_, data_stage_1__46_, data_stage_1__45_, data_stage_1__44_, data_stage_1__43_, data_stage_1__42_, data_stage_1__41_, data_stage_1__40_, data_stage_1__39_, data_stage_1__38_, data_stage_1__37_, data_stage_1__36_, data_stage_1__35_, data_stage_1__34_, data_stage_1__33_, data_stage_1__32_, data_stage_1__31_, data_stage_1__30_, data_stage_1__29_, data_stage_1__28_, data_stage_1__27_, data_stage_1__26_, data_stage_1__25_, data_stage_1__24_, data_stage_1__23_, data_stage_1__22_, data_stage_1__21_, data_stage_1__20_, data_stage_1__19_, data_stage_1__18_, data_stage_1__17_, data_stage_1__16_, data_stage_1__15_, data_stage_1__14_, data_stage_1__13_, data_stage_1__12_, data_stage_1__11_, data_stage_1__10_, data_stage_1__9_, data_stage_1__8_, data_stage_1__7_, data_stage_1__6_, data_stage_1__5_, data_stage_1__4_, data_stage_1__3_, data_stage_1__2_, data_stage_1__1_, data_stage_1__0_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_1__swap_inst
  (
    .data_i(data_i[255:128]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__255_, data_stage_1__254_, data_stage_1__253_, data_stage_1__252_, data_stage_1__251_, data_stage_1__250_, data_stage_1__249_, data_stage_1__248_, data_stage_1__247_, data_stage_1__246_, data_stage_1__245_, data_stage_1__244_, data_stage_1__243_, data_stage_1__242_, data_stage_1__241_, data_stage_1__240_, data_stage_1__239_, data_stage_1__238_, data_stage_1__237_, data_stage_1__236_, data_stage_1__235_, data_stage_1__234_, data_stage_1__233_, data_stage_1__232_, data_stage_1__231_, data_stage_1__230_, data_stage_1__229_, data_stage_1__228_, data_stage_1__227_, data_stage_1__226_, data_stage_1__225_, data_stage_1__224_, data_stage_1__223_, data_stage_1__222_, data_stage_1__221_, data_stage_1__220_, data_stage_1__219_, data_stage_1__218_, data_stage_1__217_, data_stage_1__216_, data_stage_1__215_, data_stage_1__214_, data_stage_1__213_, data_stage_1__212_, data_stage_1__211_, data_stage_1__210_, data_stage_1__209_, data_stage_1__208_, data_stage_1__207_, data_stage_1__206_, data_stage_1__205_, data_stage_1__204_, data_stage_1__203_, data_stage_1__202_, data_stage_1__201_, data_stage_1__200_, data_stage_1__199_, data_stage_1__198_, data_stage_1__197_, data_stage_1__196_, data_stage_1__195_, data_stage_1__194_, data_stage_1__193_, data_stage_1__192_, data_stage_1__191_, data_stage_1__190_, data_stage_1__189_, data_stage_1__188_, data_stage_1__187_, data_stage_1__186_, data_stage_1__185_, data_stage_1__184_, data_stage_1__183_, data_stage_1__182_, data_stage_1__181_, data_stage_1__180_, data_stage_1__179_, data_stage_1__178_, data_stage_1__177_, data_stage_1__176_, data_stage_1__175_, data_stage_1__174_, data_stage_1__173_, data_stage_1__172_, data_stage_1__171_, data_stage_1__170_, data_stage_1__169_, data_stage_1__168_, data_stage_1__167_, data_stage_1__166_, data_stage_1__165_, data_stage_1__164_, data_stage_1__163_, data_stage_1__162_, data_stage_1__161_, data_stage_1__160_, data_stage_1__159_, data_stage_1__158_, data_stage_1__157_, data_stage_1__156_, data_stage_1__155_, data_stage_1__154_, data_stage_1__153_, data_stage_1__152_, data_stage_1__151_, data_stage_1__150_, data_stage_1__149_, data_stage_1__148_, data_stage_1__147_, data_stage_1__146_, data_stage_1__145_, data_stage_1__144_, data_stage_1__143_, data_stage_1__142_, data_stage_1__141_, data_stage_1__140_, data_stage_1__139_, data_stage_1__138_, data_stage_1__137_, data_stage_1__136_, data_stage_1__135_, data_stage_1__134_, data_stage_1__133_, data_stage_1__132_, data_stage_1__131_, data_stage_1__130_, data_stage_1__129_, data_stage_1__128_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_2__swap_inst
  (
    .data_i(data_i[383:256]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__383_, data_stage_1__382_, data_stage_1__381_, data_stage_1__380_, data_stage_1__379_, data_stage_1__378_, data_stage_1__377_, data_stage_1__376_, data_stage_1__375_, data_stage_1__374_, data_stage_1__373_, data_stage_1__372_, data_stage_1__371_, data_stage_1__370_, data_stage_1__369_, data_stage_1__368_, data_stage_1__367_, data_stage_1__366_, data_stage_1__365_, data_stage_1__364_, data_stage_1__363_, data_stage_1__362_, data_stage_1__361_, data_stage_1__360_, data_stage_1__359_, data_stage_1__358_, data_stage_1__357_, data_stage_1__356_, data_stage_1__355_, data_stage_1__354_, data_stage_1__353_, data_stage_1__352_, data_stage_1__351_, data_stage_1__350_, data_stage_1__349_, data_stage_1__348_, data_stage_1__347_, data_stage_1__346_, data_stage_1__345_, data_stage_1__344_, data_stage_1__343_, data_stage_1__342_, data_stage_1__341_, data_stage_1__340_, data_stage_1__339_, data_stage_1__338_, data_stage_1__337_, data_stage_1__336_, data_stage_1__335_, data_stage_1__334_, data_stage_1__333_, data_stage_1__332_, data_stage_1__331_, data_stage_1__330_, data_stage_1__329_, data_stage_1__328_, data_stage_1__327_, data_stage_1__326_, data_stage_1__325_, data_stage_1__324_, data_stage_1__323_, data_stage_1__322_, data_stage_1__321_, data_stage_1__320_, data_stage_1__319_, data_stage_1__318_, data_stage_1__317_, data_stage_1__316_, data_stage_1__315_, data_stage_1__314_, data_stage_1__313_, data_stage_1__312_, data_stage_1__311_, data_stage_1__310_, data_stage_1__309_, data_stage_1__308_, data_stage_1__307_, data_stage_1__306_, data_stage_1__305_, data_stage_1__304_, data_stage_1__303_, data_stage_1__302_, data_stage_1__301_, data_stage_1__300_, data_stage_1__299_, data_stage_1__298_, data_stage_1__297_, data_stage_1__296_, data_stage_1__295_, data_stage_1__294_, data_stage_1__293_, data_stage_1__292_, data_stage_1__291_, data_stage_1__290_, data_stage_1__289_, data_stage_1__288_, data_stage_1__287_, data_stage_1__286_, data_stage_1__285_, data_stage_1__284_, data_stage_1__283_, data_stage_1__282_, data_stage_1__281_, data_stage_1__280_, data_stage_1__279_, data_stage_1__278_, data_stage_1__277_, data_stage_1__276_, data_stage_1__275_, data_stage_1__274_, data_stage_1__273_, data_stage_1__272_, data_stage_1__271_, data_stage_1__270_, data_stage_1__269_, data_stage_1__268_, data_stage_1__267_, data_stage_1__266_, data_stage_1__265_, data_stage_1__264_, data_stage_1__263_, data_stage_1__262_, data_stage_1__261_, data_stage_1__260_, data_stage_1__259_, data_stage_1__258_, data_stage_1__257_, data_stage_1__256_ })
  );


  bsg_swap_width_p64
  mux_stage_0__mux_swap_3__swap_inst
  (
    .data_i(data_i[511:384]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__511_, data_stage_1__510_, data_stage_1__509_, data_stage_1__508_, data_stage_1__507_, data_stage_1__506_, data_stage_1__505_, data_stage_1__504_, data_stage_1__503_, data_stage_1__502_, data_stage_1__501_, data_stage_1__500_, data_stage_1__499_, data_stage_1__498_, data_stage_1__497_, data_stage_1__496_, data_stage_1__495_, data_stage_1__494_, data_stage_1__493_, data_stage_1__492_, data_stage_1__491_, data_stage_1__490_, data_stage_1__489_, data_stage_1__488_, data_stage_1__487_, data_stage_1__486_, data_stage_1__485_, data_stage_1__484_, data_stage_1__483_, data_stage_1__482_, data_stage_1__481_, data_stage_1__480_, data_stage_1__479_, data_stage_1__478_, data_stage_1__477_, data_stage_1__476_, data_stage_1__475_, data_stage_1__474_, data_stage_1__473_, data_stage_1__472_, data_stage_1__471_, data_stage_1__470_, data_stage_1__469_, data_stage_1__468_, data_stage_1__467_, data_stage_1__466_, data_stage_1__465_, data_stage_1__464_, data_stage_1__463_, data_stage_1__462_, data_stage_1__461_, data_stage_1__460_, data_stage_1__459_, data_stage_1__458_, data_stage_1__457_, data_stage_1__456_, data_stage_1__455_, data_stage_1__454_, data_stage_1__453_, data_stage_1__452_, data_stage_1__451_, data_stage_1__450_, data_stage_1__449_, data_stage_1__448_, data_stage_1__447_, data_stage_1__446_, data_stage_1__445_, data_stage_1__444_, data_stage_1__443_, data_stage_1__442_, data_stage_1__441_, data_stage_1__440_, data_stage_1__439_, data_stage_1__438_, data_stage_1__437_, data_stage_1__436_, data_stage_1__435_, data_stage_1__434_, data_stage_1__433_, data_stage_1__432_, data_stage_1__431_, data_stage_1__430_, data_stage_1__429_, data_stage_1__428_, data_stage_1__427_, data_stage_1__426_, data_stage_1__425_, data_stage_1__424_, data_stage_1__423_, data_stage_1__422_, data_stage_1__421_, data_stage_1__420_, data_stage_1__419_, data_stage_1__418_, data_stage_1__417_, data_stage_1__416_, data_stage_1__415_, data_stage_1__414_, data_stage_1__413_, data_stage_1__412_, data_stage_1__411_, data_stage_1__410_, data_stage_1__409_, data_stage_1__408_, data_stage_1__407_, data_stage_1__406_, data_stage_1__405_, data_stage_1__404_, data_stage_1__403_, data_stage_1__402_, data_stage_1__401_, data_stage_1__400_, data_stage_1__399_, data_stage_1__398_, data_stage_1__397_, data_stage_1__396_, data_stage_1__395_, data_stage_1__394_, data_stage_1__393_, data_stage_1__392_, data_stage_1__391_, data_stage_1__390_, data_stage_1__389_, data_stage_1__388_, data_stage_1__387_, data_stage_1__386_, data_stage_1__385_, data_stage_1__384_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_1__255_, data_stage_1__254_, data_stage_1__253_, data_stage_1__252_, data_stage_1__251_, data_stage_1__250_, data_stage_1__249_, data_stage_1__248_, data_stage_1__247_, data_stage_1__246_, data_stage_1__245_, data_stage_1__244_, data_stage_1__243_, data_stage_1__242_, data_stage_1__241_, data_stage_1__240_, data_stage_1__239_, data_stage_1__238_, data_stage_1__237_, data_stage_1__236_, data_stage_1__235_, data_stage_1__234_, data_stage_1__233_, data_stage_1__232_, data_stage_1__231_, data_stage_1__230_, data_stage_1__229_, data_stage_1__228_, data_stage_1__227_, data_stage_1__226_, data_stage_1__225_, data_stage_1__224_, data_stage_1__223_, data_stage_1__222_, data_stage_1__221_, data_stage_1__220_, data_stage_1__219_, data_stage_1__218_, data_stage_1__217_, data_stage_1__216_, data_stage_1__215_, data_stage_1__214_, data_stage_1__213_, data_stage_1__212_, data_stage_1__211_, data_stage_1__210_, data_stage_1__209_, data_stage_1__208_, data_stage_1__207_, data_stage_1__206_, data_stage_1__205_, data_stage_1__204_, data_stage_1__203_, data_stage_1__202_, data_stage_1__201_, data_stage_1__200_, data_stage_1__199_, data_stage_1__198_, data_stage_1__197_, data_stage_1__196_, data_stage_1__195_, data_stage_1__194_, data_stage_1__193_, data_stage_1__192_, data_stage_1__191_, data_stage_1__190_, data_stage_1__189_, data_stage_1__188_, data_stage_1__187_, data_stage_1__186_, data_stage_1__185_, data_stage_1__184_, data_stage_1__183_, data_stage_1__182_, data_stage_1__181_, data_stage_1__180_, data_stage_1__179_, data_stage_1__178_, data_stage_1__177_, data_stage_1__176_, data_stage_1__175_, data_stage_1__174_, data_stage_1__173_, data_stage_1__172_, data_stage_1__171_, data_stage_1__170_, data_stage_1__169_, data_stage_1__168_, data_stage_1__167_, data_stage_1__166_, data_stage_1__165_, data_stage_1__164_, data_stage_1__163_, data_stage_1__162_, data_stage_1__161_, data_stage_1__160_, data_stage_1__159_, data_stage_1__158_, data_stage_1__157_, data_stage_1__156_, data_stage_1__155_, data_stage_1__154_, data_stage_1__153_, data_stage_1__152_, data_stage_1__151_, data_stage_1__150_, data_stage_1__149_, data_stage_1__148_, data_stage_1__147_, data_stage_1__146_, data_stage_1__145_, data_stage_1__144_, data_stage_1__143_, data_stage_1__142_, data_stage_1__141_, data_stage_1__140_, data_stage_1__139_, data_stage_1__138_, data_stage_1__137_, data_stage_1__136_, data_stage_1__135_, data_stage_1__134_, data_stage_1__133_, data_stage_1__132_, data_stage_1__131_, data_stage_1__130_, data_stage_1__129_, data_stage_1__128_, data_stage_1__127_, data_stage_1__126_, data_stage_1__125_, data_stage_1__124_, data_stage_1__123_, data_stage_1__122_, data_stage_1__121_, data_stage_1__120_, data_stage_1__119_, data_stage_1__118_, data_stage_1__117_, data_stage_1__116_, data_stage_1__115_, data_stage_1__114_, data_stage_1__113_, data_stage_1__112_, data_stage_1__111_, data_stage_1__110_, data_stage_1__109_, data_stage_1__108_, data_stage_1__107_, data_stage_1__106_, data_stage_1__105_, data_stage_1__104_, data_stage_1__103_, data_stage_1__102_, data_stage_1__101_, data_stage_1__100_, data_stage_1__99_, data_stage_1__98_, data_stage_1__97_, data_stage_1__96_, data_stage_1__95_, data_stage_1__94_, data_stage_1__93_, data_stage_1__92_, data_stage_1__91_, data_stage_1__90_, data_stage_1__89_, data_stage_1__88_, data_stage_1__87_, data_stage_1__86_, data_stage_1__85_, data_stage_1__84_, data_stage_1__83_, data_stage_1__82_, data_stage_1__81_, data_stage_1__80_, data_stage_1__79_, data_stage_1__78_, data_stage_1__77_, data_stage_1__76_, data_stage_1__75_, data_stage_1__74_, data_stage_1__73_, data_stage_1__72_, data_stage_1__71_, data_stage_1__70_, data_stage_1__69_, data_stage_1__68_, data_stage_1__67_, data_stage_1__66_, data_stage_1__65_, data_stage_1__64_, data_stage_1__63_, data_stage_1__62_, data_stage_1__61_, data_stage_1__60_, data_stage_1__59_, data_stage_1__58_, data_stage_1__57_, data_stage_1__56_, data_stage_1__55_, data_stage_1__54_, data_stage_1__53_, data_stage_1__52_, data_stage_1__51_, data_stage_1__50_, data_stage_1__49_, data_stage_1__48_, data_stage_1__47_, data_stage_1__46_, data_stage_1__45_, data_stage_1__44_, data_stage_1__43_, data_stage_1__42_, data_stage_1__41_, data_stage_1__40_, data_stage_1__39_, data_stage_1__38_, data_stage_1__37_, data_stage_1__36_, data_stage_1__35_, data_stage_1__34_, data_stage_1__33_, data_stage_1__32_, data_stage_1__31_, data_stage_1__30_, data_stage_1__29_, data_stage_1__28_, data_stage_1__27_, data_stage_1__26_, data_stage_1__25_, data_stage_1__24_, data_stage_1__23_, data_stage_1__22_, data_stage_1__21_, data_stage_1__20_, data_stage_1__19_, data_stage_1__18_, data_stage_1__17_, data_stage_1__16_, data_stage_1__15_, data_stage_1__14_, data_stage_1__13_, data_stage_1__12_, data_stage_1__11_, data_stage_1__10_, data_stage_1__9_, data_stage_1__8_, data_stage_1__7_, data_stage_1__6_, data_stage_1__5_, data_stage_1__4_, data_stage_1__3_, data_stage_1__2_, data_stage_1__1_, data_stage_1__0_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__255_, data_stage_2__254_, data_stage_2__253_, data_stage_2__252_, data_stage_2__251_, data_stage_2__250_, data_stage_2__249_, data_stage_2__248_, data_stage_2__247_, data_stage_2__246_, data_stage_2__245_, data_stage_2__244_, data_stage_2__243_, data_stage_2__242_, data_stage_2__241_, data_stage_2__240_, data_stage_2__239_, data_stage_2__238_, data_stage_2__237_, data_stage_2__236_, data_stage_2__235_, data_stage_2__234_, data_stage_2__233_, data_stage_2__232_, data_stage_2__231_, data_stage_2__230_, data_stage_2__229_, data_stage_2__228_, data_stage_2__227_, data_stage_2__226_, data_stage_2__225_, data_stage_2__224_, data_stage_2__223_, data_stage_2__222_, data_stage_2__221_, data_stage_2__220_, data_stage_2__219_, data_stage_2__218_, data_stage_2__217_, data_stage_2__216_, data_stage_2__215_, data_stage_2__214_, data_stage_2__213_, data_stage_2__212_, data_stage_2__211_, data_stage_2__210_, data_stage_2__209_, data_stage_2__208_, data_stage_2__207_, data_stage_2__206_, data_stage_2__205_, data_stage_2__204_, data_stage_2__203_, data_stage_2__202_, data_stage_2__201_, data_stage_2__200_, data_stage_2__199_, data_stage_2__198_, data_stage_2__197_, data_stage_2__196_, data_stage_2__195_, data_stage_2__194_, data_stage_2__193_, data_stage_2__192_, data_stage_2__191_, data_stage_2__190_, data_stage_2__189_, data_stage_2__188_, data_stage_2__187_, data_stage_2__186_, data_stage_2__185_, data_stage_2__184_, data_stage_2__183_, data_stage_2__182_, data_stage_2__181_, data_stage_2__180_, data_stage_2__179_, data_stage_2__178_, data_stage_2__177_, data_stage_2__176_, data_stage_2__175_, data_stage_2__174_, data_stage_2__173_, data_stage_2__172_, data_stage_2__171_, data_stage_2__170_, data_stage_2__169_, data_stage_2__168_, data_stage_2__167_, data_stage_2__166_, data_stage_2__165_, data_stage_2__164_, data_stage_2__163_, data_stage_2__162_, data_stage_2__161_, data_stage_2__160_, data_stage_2__159_, data_stage_2__158_, data_stage_2__157_, data_stage_2__156_, data_stage_2__155_, data_stage_2__154_, data_stage_2__153_, data_stage_2__152_, data_stage_2__151_, data_stage_2__150_, data_stage_2__149_, data_stage_2__148_, data_stage_2__147_, data_stage_2__146_, data_stage_2__145_, data_stage_2__144_, data_stage_2__143_, data_stage_2__142_, data_stage_2__141_, data_stage_2__140_, data_stage_2__139_, data_stage_2__138_, data_stage_2__137_, data_stage_2__136_, data_stage_2__135_, data_stage_2__134_, data_stage_2__133_, data_stage_2__132_, data_stage_2__131_, data_stage_2__130_, data_stage_2__129_, data_stage_2__128_, data_stage_2__127_, data_stage_2__126_, data_stage_2__125_, data_stage_2__124_, data_stage_2__123_, data_stage_2__122_, data_stage_2__121_, data_stage_2__120_, data_stage_2__119_, data_stage_2__118_, data_stage_2__117_, data_stage_2__116_, data_stage_2__115_, data_stage_2__114_, data_stage_2__113_, data_stage_2__112_, data_stage_2__111_, data_stage_2__110_, data_stage_2__109_, data_stage_2__108_, data_stage_2__107_, data_stage_2__106_, data_stage_2__105_, data_stage_2__104_, data_stage_2__103_, data_stage_2__102_, data_stage_2__101_, data_stage_2__100_, data_stage_2__99_, data_stage_2__98_, data_stage_2__97_, data_stage_2__96_, data_stage_2__95_, data_stage_2__94_, data_stage_2__93_, data_stage_2__92_, data_stage_2__91_, data_stage_2__90_, data_stage_2__89_, data_stage_2__88_, data_stage_2__87_, data_stage_2__86_, data_stage_2__85_, data_stage_2__84_, data_stage_2__83_, data_stage_2__82_, data_stage_2__81_, data_stage_2__80_, data_stage_2__79_, data_stage_2__78_, data_stage_2__77_, data_stage_2__76_, data_stage_2__75_, data_stage_2__74_, data_stage_2__73_, data_stage_2__72_, data_stage_2__71_, data_stage_2__70_, data_stage_2__69_, data_stage_2__68_, data_stage_2__67_, data_stage_2__66_, data_stage_2__65_, data_stage_2__64_, data_stage_2__63_, data_stage_2__62_, data_stage_2__61_, data_stage_2__60_, data_stage_2__59_, data_stage_2__58_, data_stage_2__57_, data_stage_2__56_, data_stage_2__55_, data_stage_2__54_, data_stage_2__53_, data_stage_2__52_, data_stage_2__51_, data_stage_2__50_, data_stage_2__49_, data_stage_2__48_, data_stage_2__47_, data_stage_2__46_, data_stage_2__45_, data_stage_2__44_, data_stage_2__43_, data_stage_2__42_, data_stage_2__41_, data_stage_2__40_, data_stage_2__39_, data_stage_2__38_, data_stage_2__37_, data_stage_2__36_, data_stage_2__35_, data_stage_2__34_, data_stage_2__33_, data_stage_2__32_, data_stage_2__31_, data_stage_2__30_, data_stage_2__29_, data_stage_2__28_, data_stage_2__27_, data_stage_2__26_, data_stage_2__25_, data_stage_2__24_, data_stage_2__23_, data_stage_2__22_, data_stage_2__21_, data_stage_2__20_, data_stage_2__19_, data_stage_2__18_, data_stage_2__17_, data_stage_2__16_, data_stage_2__15_, data_stage_2__14_, data_stage_2__13_, data_stage_2__12_, data_stage_2__11_, data_stage_2__10_, data_stage_2__9_, data_stage_2__8_, data_stage_2__7_, data_stage_2__6_, data_stage_2__5_, data_stage_2__4_, data_stage_2__3_, data_stage_2__2_, data_stage_2__1_, data_stage_2__0_ })
  );


  bsg_swap_width_p128
  mux_stage_1__mux_swap_1__swap_inst
  (
    .data_i({ data_stage_1__511_, data_stage_1__510_, data_stage_1__509_, data_stage_1__508_, data_stage_1__507_, data_stage_1__506_, data_stage_1__505_, data_stage_1__504_, data_stage_1__503_, data_stage_1__502_, data_stage_1__501_, data_stage_1__500_, data_stage_1__499_, data_stage_1__498_, data_stage_1__497_, data_stage_1__496_, data_stage_1__495_, data_stage_1__494_, data_stage_1__493_, data_stage_1__492_, data_stage_1__491_, data_stage_1__490_, data_stage_1__489_, data_stage_1__488_, data_stage_1__487_, data_stage_1__486_, data_stage_1__485_, data_stage_1__484_, data_stage_1__483_, data_stage_1__482_, data_stage_1__481_, data_stage_1__480_, data_stage_1__479_, data_stage_1__478_, data_stage_1__477_, data_stage_1__476_, data_stage_1__475_, data_stage_1__474_, data_stage_1__473_, data_stage_1__472_, data_stage_1__471_, data_stage_1__470_, data_stage_1__469_, data_stage_1__468_, data_stage_1__467_, data_stage_1__466_, data_stage_1__465_, data_stage_1__464_, data_stage_1__463_, data_stage_1__462_, data_stage_1__461_, data_stage_1__460_, data_stage_1__459_, data_stage_1__458_, data_stage_1__457_, data_stage_1__456_, data_stage_1__455_, data_stage_1__454_, data_stage_1__453_, data_stage_1__452_, data_stage_1__451_, data_stage_1__450_, data_stage_1__449_, data_stage_1__448_, data_stage_1__447_, data_stage_1__446_, data_stage_1__445_, data_stage_1__444_, data_stage_1__443_, data_stage_1__442_, data_stage_1__441_, data_stage_1__440_, data_stage_1__439_, data_stage_1__438_, data_stage_1__437_, data_stage_1__436_, data_stage_1__435_, data_stage_1__434_, data_stage_1__433_, data_stage_1__432_, data_stage_1__431_, data_stage_1__430_, data_stage_1__429_, data_stage_1__428_, data_stage_1__427_, data_stage_1__426_, data_stage_1__425_, data_stage_1__424_, data_stage_1__423_, data_stage_1__422_, data_stage_1__421_, data_stage_1__420_, data_stage_1__419_, data_stage_1__418_, data_stage_1__417_, data_stage_1__416_, data_stage_1__415_, data_stage_1__414_, data_stage_1__413_, data_stage_1__412_, data_stage_1__411_, data_stage_1__410_, data_stage_1__409_, data_stage_1__408_, data_stage_1__407_, data_stage_1__406_, data_stage_1__405_, data_stage_1__404_, data_stage_1__403_, data_stage_1__402_, data_stage_1__401_, data_stage_1__400_, data_stage_1__399_, data_stage_1__398_, data_stage_1__397_, data_stage_1__396_, data_stage_1__395_, data_stage_1__394_, data_stage_1__393_, data_stage_1__392_, data_stage_1__391_, data_stage_1__390_, data_stage_1__389_, data_stage_1__388_, data_stage_1__387_, data_stage_1__386_, data_stage_1__385_, data_stage_1__384_, data_stage_1__383_, data_stage_1__382_, data_stage_1__381_, data_stage_1__380_, data_stage_1__379_, data_stage_1__378_, data_stage_1__377_, data_stage_1__376_, data_stage_1__375_, data_stage_1__374_, data_stage_1__373_, data_stage_1__372_, data_stage_1__371_, data_stage_1__370_, data_stage_1__369_, data_stage_1__368_, data_stage_1__367_, data_stage_1__366_, data_stage_1__365_, data_stage_1__364_, data_stage_1__363_, data_stage_1__362_, data_stage_1__361_, data_stage_1__360_, data_stage_1__359_, data_stage_1__358_, data_stage_1__357_, data_stage_1__356_, data_stage_1__355_, data_stage_1__354_, data_stage_1__353_, data_stage_1__352_, data_stage_1__351_, data_stage_1__350_, data_stage_1__349_, data_stage_1__348_, data_stage_1__347_, data_stage_1__346_, data_stage_1__345_, data_stage_1__344_, data_stage_1__343_, data_stage_1__342_, data_stage_1__341_, data_stage_1__340_, data_stage_1__339_, data_stage_1__338_, data_stage_1__337_, data_stage_1__336_, data_stage_1__335_, data_stage_1__334_, data_stage_1__333_, data_stage_1__332_, data_stage_1__331_, data_stage_1__330_, data_stage_1__329_, data_stage_1__328_, data_stage_1__327_, data_stage_1__326_, data_stage_1__325_, data_stage_1__324_, data_stage_1__323_, data_stage_1__322_, data_stage_1__321_, data_stage_1__320_, data_stage_1__319_, data_stage_1__318_, data_stage_1__317_, data_stage_1__316_, data_stage_1__315_, data_stage_1__314_, data_stage_1__313_, data_stage_1__312_, data_stage_1__311_, data_stage_1__310_, data_stage_1__309_, data_stage_1__308_, data_stage_1__307_, data_stage_1__306_, data_stage_1__305_, data_stage_1__304_, data_stage_1__303_, data_stage_1__302_, data_stage_1__301_, data_stage_1__300_, data_stage_1__299_, data_stage_1__298_, data_stage_1__297_, data_stage_1__296_, data_stage_1__295_, data_stage_1__294_, data_stage_1__293_, data_stage_1__292_, data_stage_1__291_, data_stage_1__290_, data_stage_1__289_, data_stage_1__288_, data_stage_1__287_, data_stage_1__286_, data_stage_1__285_, data_stage_1__284_, data_stage_1__283_, data_stage_1__282_, data_stage_1__281_, data_stage_1__280_, data_stage_1__279_, data_stage_1__278_, data_stage_1__277_, data_stage_1__276_, data_stage_1__275_, data_stage_1__274_, data_stage_1__273_, data_stage_1__272_, data_stage_1__271_, data_stage_1__270_, data_stage_1__269_, data_stage_1__268_, data_stage_1__267_, data_stage_1__266_, data_stage_1__265_, data_stage_1__264_, data_stage_1__263_, data_stage_1__262_, data_stage_1__261_, data_stage_1__260_, data_stage_1__259_, data_stage_1__258_, data_stage_1__257_, data_stage_1__256_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__511_, data_stage_2__510_, data_stage_2__509_, data_stage_2__508_, data_stage_2__507_, data_stage_2__506_, data_stage_2__505_, data_stage_2__504_, data_stage_2__503_, data_stage_2__502_, data_stage_2__501_, data_stage_2__500_, data_stage_2__499_, data_stage_2__498_, data_stage_2__497_, data_stage_2__496_, data_stage_2__495_, data_stage_2__494_, data_stage_2__493_, data_stage_2__492_, data_stage_2__491_, data_stage_2__490_, data_stage_2__489_, data_stage_2__488_, data_stage_2__487_, data_stage_2__486_, data_stage_2__485_, data_stage_2__484_, data_stage_2__483_, data_stage_2__482_, data_stage_2__481_, data_stage_2__480_, data_stage_2__479_, data_stage_2__478_, data_stage_2__477_, data_stage_2__476_, data_stage_2__475_, data_stage_2__474_, data_stage_2__473_, data_stage_2__472_, data_stage_2__471_, data_stage_2__470_, data_stage_2__469_, data_stage_2__468_, data_stage_2__467_, data_stage_2__466_, data_stage_2__465_, data_stage_2__464_, data_stage_2__463_, data_stage_2__462_, data_stage_2__461_, data_stage_2__460_, data_stage_2__459_, data_stage_2__458_, data_stage_2__457_, data_stage_2__456_, data_stage_2__455_, data_stage_2__454_, data_stage_2__453_, data_stage_2__452_, data_stage_2__451_, data_stage_2__450_, data_stage_2__449_, data_stage_2__448_, data_stage_2__447_, data_stage_2__446_, data_stage_2__445_, data_stage_2__444_, data_stage_2__443_, data_stage_2__442_, data_stage_2__441_, data_stage_2__440_, data_stage_2__439_, data_stage_2__438_, data_stage_2__437_, data_stage_2__436_, data_stage_2__435_, data_stage_2__434_, data_stage_2__433_, data_stage_2__432_, data_stage_2__431_, data_stage_2__430_, data_stage_2__429_, data_stage_2__428_, data_stage_2__427_, data_stage_2__426_, data_stage_2__425_, data_stage_2__424_, data_stage_2__423_, data_stage_2__422_, data_stage_2__421_, data_stage_2__420_, data_stage_2__419_, data_stage_2__418_, data_stage_2__417_, data_stage_2__416_, data_stage_2__415_, data_stage_2__414_, data_stage_2__413_, data_stage_2__412_, data_stage_2__411_, data_stage_2__410_, data_stage_2__409_, data_stage_2__408_, data_stage_2__407_, data_stage_2__406_, data_stage_2__405_, data_stage_2__404_, data_stage_2__403_, data_stage_2__402_, data_stage_2__401_, data_stage_2__400_, data_stage_2__399_, data_stage_2__398_, data_stage_2__397_, data_stage_2__396_, data_stage_2__395_, data_stage_2__394_, data_stage_2__393_, data_stage_2__392_, data_stage_2__391_, data_stage_2__390_, data_stage_2__389_, data_stage_2__388_, data_stage_2__387_, data_stage_2__386_, data_stage_2__385_, data_stage_2__384_, data_stage_2__383_, data_stage_2__382_, data_stage_2__381_, data_stage_2__380_, data_stage_2__379_, data_stage_2__378_, data_stage_2__377_, data_stage_2__376_, data_stage_2__375_, data_stage_2__374_, data_stage_2__373_, data_stage_2__372_, data_stage_2__371_, data_stage_2__370_, data_stage_2__369_, data_stage_2__368_, data_stage_2__367_, data_stage_2__366_, data_stage_2__365_, data_stage_2__364_, data_stage_2__363_, data_stage_2__362_, data_stage_2__361_, data_stage_2__360_, data_stage_2__359_, data_stage_2__358_, data_stage_2__357_, data_stage_2__356_, data_stage_2__355_, data_stage_2__354_, data_stage_2__353_, data_stage_2__352_, data_stage_2__351_, data_stage_2__350_, data_stage_2__349_, data_stage_2__348_, data_stage_2__347_, data_stage_2__346_, data_stage_2__345_, data_stage_2__344_, data_stage_2__343_, data_stage_2__342_, data_stage_2__341_, data_stage_2__340_, data_stage_2__339_, data_stage_2__338_, data_stage_2__337_, data_stage_2__336_, data_stage_2__335_, data_stage_2__334_, data_stage_2__333_, data_stage_2__332_, data_stage_2__331_, data_stage_2__330_, data_stage_2__329_, data_stage_2__328_, data_stage_2__327_, data_stage_2__326_, data_stage_2__325_, data_stage_2__324_, data_stage_2__323_, data_stage_2__322_, data_stage_2__321_, data_stage_2__320_, data_stage_2__319_, data_stage_2__318_, data_stage_2__317_, data_stage_2__316_, data_stage_2__315_, data_stage_2__314_, data_stage_2__313_, data_stage_2__312_, data_stage_2__311_, data_stage_2__310_, data_stage_2__309_, data_stage_2__308_, data_stage_2__307_, data_stage_2__306_, data_stage_2__305_, data_stage_2__304_, data_stage_2__303_, data_stage_2__302_, data_stage_2__301_, data_stage_2__300_, data_stage_2__299_, data_stage_2__298_, data_stage_2__297_, data_stage_2__296_, data_stage_2__295_, data_stage_2__294_, data_stage_2__293_, data_stage_2__292_, data_stage_2__291_, data_stage_2__290_, data_stage_2__289_, data_stage_2__288_, data_stage_2__287_, data_stage_2__286_, data_stage_2__285_, data_stage_2__284_, data_stage_2__283_, data_stage_2__282_, data_stage_2__281_, data_stage_2__280_, data_stage_2__279_, data_stage_2__278_, data_stage_2__277_, data_stage_2__276_, data_stage_2__275_, data_stage_2__274_, data_stage_2__273_, data_stage_2__272_, data_stage_2__271_, data_stage_2__270_, data_stage_2__269_, data_stage_2__268_, data_stage_2__267_, data_stage_2__266_, data_stage_2__265_, data_stage_2__264_, data_stage_2__263_, data_stage_2__262_, data_stage_2__261_, data_stage_2__260_, data_stage_2__259_, data_stage_2__258_, data_stage_2__257_, data_stage_2__256_ })
  );


  bsg_swap_width_p256
  mux_stage_2__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_2__511_, data_stage_2__510_, data_stage_2__509_, data_stage_2__508_, data_stage_2__507_, data_stage_2__506_, data_stage_2__505_, data_stage_2__504_, data_stage_2__503_, data_stage_2__502_, data_stage_2__501_, data_stage_2__500_, data_stage_2__499_, data_stage_2__498_, data_stage_2__497_, data_stage_2__496_, data_stage_2__495_, data_stage_2__494_, data_stage_2__493_, data_stage_2__492_, data_stage_2__491_, data_stage_2__490_, data_stage_2__489_, data_stage_2__488_, data_stage_2__487_, data_stage_2__486_, data_stage_2__485_, data_stage_2__484_, data_stage_2__483_, data_stage_2__482_, data_stage_2__481_, data_stage_2__480_, data_stage_2__479_, data_stage_2__478_, data_stage_2__477_, data_stage_2__476_, data_stage_2__475_, data_stage_2__474_, data_stage_2__473_, data_stage_2__472_, data_stage_2__471_, data_stage_2__470_, data_stage_2__469_, data_stage_2__468_, data_stage_2__467_, data_stage_2__466_, data_stage_2__465_, data_stage_2__464_, data_stage_2__463_, data_stage_2__462_, data_stage_2__461_, data_stage_2__460_, data_stage_2__459_, data_stage_2__458_, data_stage_2__457_, data_stage_2__456_, data_stage_2__455_, data_stage_2__454_, data_stage_2__453_, data_stage_2__452_, data_stage_2__451_, data_stage_2__450_, data_stage_2__449_, data_stage_2__448_, data_stage_2__447_, data_stage_2__446_, data_stage_2__445_, data_stage_2__444_, data_stage_2__443_, data_stage_2__442_, data_stage_2__441_, data_stage_2__440_, data_stage_2__439_, data_stage_2__438_, data_stage_2__437_, data_stage_2__436_, data_stage_2__435_, data_stage_2__434_, data_stage_2__433_, data_stage_2__432_, data_stage_2__431_, data_stage_2__430_, data_stage_2__429_, data_stage_2__428_, data_stage_2__427_, data_stage_2__426_, data_stage_2__425_, data_stage_2__424_, data_stage_2__423_, data_stage_2__422_, data_stage_2__421_, data_stage_2__420_, data_stage_2__419_, data_stage_2__418_, data_stage_2__417_, data_stage_2__416_, data_stage_2__415_, data_stage_2__414_, data_stage_2__413_, data_stage_2__412_, data_stage_2__411_, data_stage_2__410_, data_stage_2__409_, data_stage_2__408_, data_stage_2__407_, data_stage_2__406_, data_stage_2__405_, data_stage_2__404_, data_stage_2__403_, data_stage_2__402_, data_stage_2__401_, data_stage_2__400_, data_stage_2__399_, data_stage_2__398_, data_stage_2__397_, data_stage_2__396_, data_stage_2__395_, data_stage_2__394_, data_stage_2__393_, data_stage_2__392_, data_stage_2__391_, data_stage_2__390_, data_stage_2__389_, data_stage_2__388_, data_stage_2__387_, data_stage_2__386_, data_stage_2__385_, data_stage_2__384_, data_stage_2__383_, data_stage_2__382_, data_stage_2__381_, data_stage_2__380_, data_stage_2__379_, data_stage_2__378_, data_stage_2__377_, data_stage_2__376_, data_stage_2__375_, data_stage_2__374_, data_stage_2__373_, data_stage_2__372_, data_stage_2__371_, data_stage_2__370_, data_stage_2__369_, data_stage_2__368_, data_stage_2__367_, data_stage_2__366_, data_stage_2__365_, data_stage_2__364_, data_stage_2__363_, data_stage_2__362_, data_stage_2__361_, data_stage_2__360_, data_stage_2__359_, data_stage_2__358_, data_stage_2__357_, data_stage_2__356_, data_stage_2__355_, data_stage_2__354_, data_stage_2__353_, data_stage_2__352_, data_stage_2__351_, data_stage_2__350_, data_stage_2__349_, data_stage_2__348_, data_stage_2__347_, data_stage_2__346_, data_stage_2__345_, data_stage_2__344_, data_stage_2__343_, data_stage_2__342_, data_stage_2__341_, data_stage_2__340_, data_stage_2__339_, data_stage_2__338_, data_stage_2__337_, data_stage_2__336_, data_stage_2__335_, data_stage_2__334_, data_stage_2__333_, data_stage_2__332_, data_stage_2__331_, data_stage_2__330_, data_stage_2__329_, data_stage_2__328_, data_stage_2__327_, data_stage_2__326_, data_stage_2__325_, data_stage_2__324_, data_stage_2__323_, data_stage_2__322_, data_stage_2__321_, data_stage_2__320_, data_stage_2__319_, data_stage_2__318_, data_stage_2__317_, data_stage_2__316_, data_stage_2__315_, data_stage_2__314_, data_stage_2__313_, data_stage_2__312_, data_stage_2__311_, data_stage_2__310_, data_stage_2__309_, data_stage_2__308_, data_stage_2__307_, data_stage_2__306_, data_stage_2__305_, data_stage_2__304_, data_stage_2__303_, data_stage_2__302_, data_stage_2__301_, data_stage_2__300_, data_stage_2__299_, data_stage_2__298_, data_stage_2__297_, data_stage_2__296_, data_stage_2__295_, data_stage_2__294_, data_stage_2__293_, data_stage_2__292_, data_stage_2__291_, data_stage_2__290_, data_stage_2__289_, data_stage_2__288_, data_stage_2__287_, data_stage_2__286_, data_stage_2__285_, data_stage_2__284_, data_stage_2__283_, data_stage_2__282_, data_stage_2__281_, data_stage_2__280_, data_stage_2__279_, data_stage_2__278_, data_stage_2__277_, data_stage_2__276_, data_stage_2__275_, data_stage_2__274_, data_stage_2__273_, data_stage_2__272_, data_stage_2__271_, data_stage_2__270_, data_stage_2__269_, data_stage_2__268_, data_stage_2__267_, data_stage_2__266_, data_stage_2__265_, data_stage_2__264_, data_stage_2__263_, data_stage_2__262_, data_stage_2__261_, data_stage_2__260_, data_stage_2__259_, data_stage_2__258_, data_stage_2__257_, data_stage_2__256_, data_stage_2__255_, data_stage_2__254_, data_stage_2__253_, data_stage_2__252_, data_stage_2__251_, data_stage_2__250_, data_stage_2__249_, data_stage_2__248_, data_stage_2__247_, data_stage_2__246_, data_stage_2__245_, data_stage_2__244_, data_stage_2__243_, data_stage_2__242_, data_stage_2__241_, data_stage_2__240_, data_stage_2__239_, data_stage_2__238_, data_stage_2__237_, data_stage_2__236_, data_stage_2__235_, data_stage_2__234_, data_stage_2__233_, data_stage_2__232_, data_stage_2__231_, data_stage_2__230_, data_stage_2__229_, data_stage_2__228_, data_stage_2__227_, data_stage_2__226_, data_stage_2__225_, data_stage_2__224_, data_stage_2__223_, data_stage_2__222_, data_stage_2__221_, data_stage_2__220_, data_stage_2__219_, data_stage_2__218_, data_stage_2__217_, data_stage_2__216_, data_stage_2__215_, data_stage_2__214_, data_stage_2__213_, data_stage_2__212_, data_stage_2__211_, data_stage_2__210_, data_stage_2__209_, data_stage_2__208_, data_stage_2__207_, data_stage_2__206_, data_stage_2__205_, data_stage_2__204_, data_stage_2__203_, data_stage_2__202_, data_stage_2__201_, data_stage_2__200_, data_stage_2__199_, data_stage_2__198_, data_stage_2__197_, data_stage_2__196_, data_stage_2__195_, data_stage_2__194_, data_stage_2__193_, data_stage_2__192_, data_stage_2__191_, data_stage_2__190_, data_stage_2__189_, data_stage_2__188_, data_stage_2__187_, data_stage_2__186_, data_stage_2__185_, data_stage_2__184_, data_stage_2__183_, data_stage_2__182_, data_stage_2__181_, data_stage_2__180_, data_stage_2__179_, data_stage_2__178_, data_stage_2__177_, data_stage_2__176_, data_stage_2__175_, data_stage_2__174_, data_stage_2__173_, data_stage_2__172_, data_stage_2__171_, data_stage_2__170_, data_stage_2__169_, data_stage_2__168_, data_stage_2__167_, data_stage_2__166_, data_stage_2__165_, data_stage_2__164_, data_stage_2__163_, data_stage_2__162_, data_stage_2__161_, data_stage_2__160_, data_stage_2__159_, data_stage_2__158_, data_stage_2__157_, data_stage_2__156_, data_stage_2__155_, data_stage_2__154_, data_stage_2__153_, data_stage_2__152_, data_stage_2__151_, data_stage_2__150_, data_stage_2__149_, data_stage_2__148_, data_stage_2__147_, data_stage_2__146_, data_stage_2__145_, data_stage_2__144_, data_stage_2__143_, data_stage_2__142_, data_stage_2__141_, data_stage_2__140_, data_stage_2__139_, data_stage_2__138_, data_stage_2__137_, data_stage_2__136_, data_stage_2__135_, data_stage_2__134_, data_stage_2__133_, data_stage_2__132_, data_stage_2__131_, data_stage_2__130_, data_stage_2__129_, data_stage_2__128_, data_stage_2__127_, data_stage_2__126_, data_stage_2__125_, data_stage_2__124_, data_stage_2__123_, data_stage_2__122_, data_stage_2__121_, data_stage_2__120_, data_stage_2__119_, data_stage_2__118_, data_stage_2__117_, data_stage_2__116_, data_stage_2__115_, data_stage_2__114_, data_stage_2__113_, data_stage_2__112_, data_stage_2__111_, data_stage_2__110_, data_stage_2__109_, data_stage_2__108_, data_stage_2__107_, data_stage_2__106_, data_stage_2__105_, data_stage_2__104_, data_stage_2__103_, data_stage_2__102_, data_stage_2__101_, data_stage_2__100_, data_stage_2__99_, data_stage_2__98_, data_stage_2__97_, data_stage_2__96_, data_stage_2__95_, data_stage_2__94_, data_stage_2__93_, data_stage_2__92_, data_stage_2__91_, data_stage_2__90_, data_stage_2__89_, data_stage_2__88_, data_stage_2__87_, data_stage_2__86_, data_stage_2__85_, data_stage_2__84_, data_stage_2__83_, data_stage_2__82_, data_stage_2__81_, data_stage_2__80_, data_stage_2__79_, data_stage_2__78_, data_stage_2__77_, data_stage_2__76_, data_stage_2__75_, data_stage_2__74_, data_stage_2__73_, data_stage_2__72_, data_stage_2__71_, data_stage_2__70_, data_stage_2__69_, data_stage_2__68_, data_stage_2__67_, data_stage_2__66_, data_stage_2__65_, data_stage_2__64_, data_stage_2__63_, data_stage_2__62_, data_stage_2__61_, data_stage_2__60_, data_stage_2__59_, data_stage_2__58_, data_stage_2__57_, data_stage_2__56_, data_stage_2__55_, data_stage_2__54_, data_stage_2__53_, data_stage_2__52_, data_stage_2__51_, data_stage_2__50_, data_stage_2__49_, data_stage_2__48_, data_stage_2__47_, data_stage_2__46_, data_stage_2__45_, data_stage_2__44_, data_stage_2__43_, data_stage_2__42_, data_stage_2__41_, data_stage_2__40_, data_stage_2__39_, data_stage_2__38_, data_stage_2__37_, data_stage_2__36_, data_stage_2__35_, data_stage_2__34_, data_stage_2__33_, data_stage_2__32_, data_stage_2__31_, data_stage_2__30_, data_stage_2__29_, data_stage_2__28_, data_stage_2__27_, data_stage_2__26_, data_stage_2__25_, data_stage_2__24_, data_stage_2__23_, data_stage_2__22_, data_stage_2__21_, data_stage_2__20_, data_stage_2__19_, data_stage_2__18_, data_stage_2__17_, data_stage_2__16_, data_stage_2__15_, data_stage_2__14_, data_stage_2__13_, data_stage_2__12_, data_stage_2__11_, data_stage_2__10_, data_stage_2__9_, data_stage_2__8_, data_stage_2__7_, data_stage_2__6_, data_stage_2__5_, data_stage_2__4_, data_stage_2__3_, data_stage_2__2_, data_stage_2__1_, data_stage_2__0_ }),
    .swap_i(sel_i[2]),
    .data_o(data_o)
  );


endmodule



module bsg_decode_num_out_p8
(
  i,
  o
);

  input [2:0] i;
  output [7:0] o;
  wire [7:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_lru_pseudo_tree_decode_ways_p8
(
  way_id_i,
  data_o,
  mask_o
);

  input [2:0] way_id_i;
  output [6:0] data_o;
  output [6:0] mask_o;
  wire [6:0] data_o,mask_o;
  wire N0,N1,N2;
  assign mask_o[0] = 1'b1;
  assign data_o[0] = 1'b1 & N0;
  assign N0 = ~way_id_i[2];
  assign mask_o[1] = 1'b1 & N0;
  assign data_o[1] = mask_o[1] & N1;
  assign N1 = ~way_id_i[1];
  assign mask_o[2] = 1'b1 & way_id_i[2];
  assign data_o[2] = mask_o[2] & N1;
  assign mask_o[3] = mask_o[1] & N1;
  assign data_o[3] = mask_o[3] & N2;
  assign N2 = ~way_id_i[0];
  assign mask_o[4] = mask_o[1] & way_id_i[1];
  assign data_o[4] = mask_o[4] & N2;
  assign mask_o[5] = mask_o[2] & N1;
  assign data_o[5] = mask_o[5] & N2;
  assign mask_o[6] = mask_o[2] & way_id_i[1];
  assign data_o[6] = mask_o[6] & N2;

endmodule



module icache_eaddr_width_p64_paddr_width_p22_data_width_p64_instr_width_p32_num_cce_p1_num_lce_p2_ways_p8_sets_p64
(
  clk_i,
  reset_i,
  id_i,
  pc_gen_icache_vaddr_i,
  pc_gen_icache_vaddr_v_i,
  pc_gen_icache_vaddr_ready_o,
  icache_pc_gen_data_o,
  icache_pc_gen_data_v_o,
  icache_pc_gen_data_ready_i,
  itlb_icache_data_resp_i,
  itlb_icache_data_resp_v_i,
  itlb_icache_data_resp_ready_o,
  cache_miss_o,
  poison_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i
);

  input [0:0] id_i;
  input [63:0] pc_gen_icache_vaddr_i;
  output [95:0] icache_pc_gen_data_o;
  input [9:0] itlb_icache_data_resp_i;
  output [96:0] lce_req_o;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  input [35:0] lce_cmd_i;
  input [517:0] lce_data_cmd_i;
  output [517:0] lce_data_cmd_o;
  input clk_i;
  input reset_i;
  input pc_gen_icache_vaddr_v_i;
  input icache_pc_gen_data_ready_i;
  input itlb_icache_data_resp_v_i;
  input poison_i;
  input lce_req_ready_i;
  input lce_resp_ready_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_v_i;
  input lce_data_cmd_ready_i;
  output pc_gen_icache_vaddr_ready_o;
  output icache_pc_gen_data_v_o;
  output itlb_icache_data_resp_ready_o;
  output cache_miss_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_ready_o;
  output lce_data_cmd_ready_o;
  output lce_data_cmd_v_o;
  wire [96:0] lce_req_o;
  wire [25:0] lce_resp_o;
  wire [536:0] lce_data_resp_o;
  wire [517:0] lce_data_cmd_o;
  wire pc_gen_icache_vaddr_ready_o,icache_pc_gen_data_v_o,cache_miss_o,lce_req_v_o,
  lce_resp_v_o,lce_data_resp_v_o,lce_cmd_ready_o,lce_data_cmd_ready_o,
  lce_data_cmd_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,tl_we,N16,N17,N18,N19,
  n_0_net_,tag_mem_w_li,tag_mem_v_li,n_1_net_,n_2_net_,n_3_net_,n_4_net_,n_5_net_,
  n_6_net_,n_7_net_,n_8_net_,tv_we,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,
  N32,N33,N34,N35,N36,N37,hit,miss_v,n_9_net_,metadata_mem_w_li,metadata_mem_v_li,
  n_10_net__7_,n_10_net__6_,n_10_net__5_,n_10_net__4_,n_10_net__3_,n_10_net__2_,
  n_10_net__1_,n_10_net__0_,invalid_exist,N38,data_mem_pkt_v_lo,data_mem_pkt_yumi_li,
  tag_mem_pkt_v_lo,tag_mem_pkt_yumi_li,metadata_mem_pkt_v_lo,
  metadata_mem_pkt_yumi_li,n_11_net__2_,n_11_net__1_,n_11_net__0_,N39,N40,N41,N42,N43,N44,N45,N46,N47,
  N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,
  N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,
  N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98;
  wire [95:0] tag_mem_data_li,tag_mem_w_mask_li,tag_mem_data_lo;
  wire [5:0] tag_mem_addr_li,metadata_mem_addr_li;
  wire [511:0] data_mem_bank_data_li,data_mem_bank_data_lo,data_mem_data_li;
  wire [71:0] data_mem_bank_addr_li;
  wire [7:0] data_mem_bank_w_li,data_mem_bank_v_li,hit_v,lce_tag_mem_way_one_hot;
  wire [2:0] hit_index,lru_encode,way_invalid_index,lru_way_li;
  wire [6:0] metadata_mem_data_li,metadata_mem_mask_li,metadata_mem_data_lo,
  lru_decode_data_lo,lru_decode_mask_lo;
  wire [521:0] data_mem_pkt;
  wire [22:0] tag_mem_pkt;
  wire [9:0] metadata_mem_pkt;
  wire [63:0] ld_data_way_picked;
  reg [11:0] vaddr_tl_r;
  reg itlb_icache_data_resp_ready_o,v_tv_r;
  reg [63:0] eaddr_tl_r;
  reg [15:0] state_tv_r;
  reg [511:0] ld_data_tv_r;
  reg [21:0] addr_tv_r;
  reg [95:0] icache_pc_gen_data_o;
  reg [79:0] tag_tv_r;
  reg [2:0] data_mem_pkt_way_r;

  bsg_mem_1rw_sync_mask_write_bit_width_p96_els_p64
  tag_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(tag_mem_data_li),
    .addr_i(tag_mem_addr_li),
    .v_i(n_0_net_),
    .w_mask_i(tag_mem_w_mask_li),
    .w_i(tag_mem_w_li),
    .data_o(tag_mem_data_lo)
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_banks_0__data_mem_bank
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_1_net_),
    .w_i(data_mem_bank_w_li[0]),
    .addr_i(data_mem_bank_addr_li[8:0]),
    .data_i(data_mem_bank_data_li[63:0]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_bank_data_lo[63:0])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_banks_1__data_mem_bank
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_2_net_),
    .w_i(data_mem_bank_w_li[1]),
    .addr_i(data_mem_bank_addr_li[17:9]),
    .data_i(data_mem_bank_data_li[127:64]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_bank_data_lo[127:64])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_banks_2__data_mem_bank
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_3_net_),
    .w_i(data_mem_bank_w_li[2]),
    .addr_i(data_mem_bank_addr_li[26:18]),
    .data_i(data_mem_bank_data_li[191:128]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_bank_data_lo[191:128])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_banks_3__data_mem_bank
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_4_net_),
    .w_i(data_mem_bank_w_li[3]),
    .addr_i(data_mem_bank_addr_li[35:27]),
    .data_i(data_mem_bank_data_li[255:192]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_bank_data_lo[255:192])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_banks_4__data_mem_bank
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_5_net_),
    .w_i(data_mem_bank_w_li[4]),
    .addr_i(data_mem_bank_addr_li[44:36]),
    .data_i(data_mem_bank_data_li[319:256]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_bank_data_lo[319:256])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_banks_5__data_mem_bank
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_6_net_),
    .w_i(data_mem_bank_w_li[5]),
    .addr_i(data_mem_bank_addr_li[53:45]),
    .data_i(data_mem_bank_data_li[383:320]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_bank_data_lo[383:320])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_banks_6__data_mem_bank
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_7_net_),
    .w_i(data_mem_bank_w_li[6]),
    .addr_i(data_mem_bank_addr_li[62:54]),
    .data_i(data_mem_bank_data_li[447:384]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_bank_data_lo[447:384])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_banks_7__data_mem_bank
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_8_net_),
    .w_i(data_mem_bank_w_li[7]),
    .addr_i(data_mem_bank_addr_li[71:63]),
    .data_i(data_mem_bank_data_li[511:448]),
    .write_mask_i({ 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 }),
    .data_o(data_mem_bank_data_lo[511:448])
  );

  assign N30 = tag_tv_r[9:0] == addr_tv_r[21:12];
  assign N31 = tag_tv_r[19:10] == addr_tv_r[21:12];
  assign N32 = tag_tv_r[29:20] == addr_tv_r[21:12];
  assign N33 = tag_tv_r[39:30] == addr_tv_r[21:12];
  assign N34 = tag_tv_r[49:40] == addr_tv_r[21:12];
  assign N35 = tag_tv_r[59:50] == addr_tv_r[21:12];
  assign N36 = tag_tv_r[69:60] == addr_tv_r[21:12];
  assign N37 = tag_tv_r[79:70] == addr_tv_r[21:12];

  bsg_priority_encode_width_p8_lo_to_hi_p1
  pe_load_hit
  (
    .i(hit_v),
    .addr_o(hit_index),
    .v_o(hit)
  );


  bsg_mem_1rw_sync_mask_write_bit_width_p7_els_p64
  metadata_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(metadata_mem_data_li),
    .addr_i(metadata_mem_addr_li),
    .v_i(n_9_net_),
    .w_mask_i(metadata_mem_mask_li),
    .w_i(metadata_mem_w_li),
    .data_o(metadata_mem_data_lo)
  );


  bsg_lru_pseudo_tree_encode_ways_p8
  lru_encoder
  (
    .lru_i(metadata_mem_data_lo),
    .way_id_o(lru_encode)
  );


  bsg_priority_encode_width_p8_lo_to_hi_p1
  pe_invalid
  (
    .i({ n_10_net__7_, n_10_net__6_, n_10_net__5_, n_10_net__4_, n_10_net__3_, n_10_net__2_, n_10_net__1_, n_10_net__0_ }),
    .addr_o(way_invalid_index),
    .v_o(invalid_exist)
  );


  bp_fe_lce_data_width_p64_paddr_width_p22_lce_data_width_p512_sets_p64_ways_p8_num_cce_p1_num_lce_p2
  lce
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .id_i(id_i[0]),
    .ready_o(pc_gen_icache_vaddr_ready_o),
    .cache_miss_o(cache_miss_o),
    .miss_i(miss_v),
    .miss_addr_i(addr_tv_r),
    .data_mem_data_i(data_mem_data_li),
    .data_mem_pkt_o(data_mem_pkt),
    .data_mem_pkt_v_o(data_mem_pkt_v_lo),
    .data_mem_pkt_yumi_i(data_mem_pkt_yumi_li),
    .tag_mem_pkt_o(tag_mem_pkt),
    .tag_mem_pkt_v_o(tag_mem_pkt_v_lo),
    .tag_mem_pkt_yumi_i(tag_mem_pkt_yumi_li),
    .metadata_mem_pkt_v_o(metadata_mem_pkt_v_lo),
    .metadata_mem_pkt_o(metadata_mem_pkt),
    .lru_way_i(lru_way_li),
    .metadata_mem_pkt_yumi_i(metadata_mem_pkt_yumi_li),
    .lce_req_o(lce_req_o),
    .lce_req_v_o(lce_req_v_o),
    .lce_req_ready_i(lce_req_ready_i),
    .lce_resp_o(lce_resp_o),
    .lce_resp_v_o(lce_resp_v_o),
    .lce_resp_ready_i(lce_resp_ready_i),
    .lce_data_resp_o(lce_data_resp_o),
    .lce_data_resp_v_o(lce_data_resp_v_o),
    .lce_data_resp_ready_i(lce_data_resp_ready_i),
    .lce_cmd_i(lce_cmd_i),
    .lce_cmd_v_i(lce_cmd_v_i),
    .lce_cmd_ready_o(lce_cmd_ready_o),
    .lce_data_cmd_i(lce_data_cmd_i),
    .lce_data_cmd_v_i(lce_data_cmd_v_i),
    .lce_data_cmd_ready_o(lce_data_cmd_ready_o),
    .lce_data_cmd_o(lce_data_cmd_o),
    .lce_data_cmd_v_o(lce_data_cmd_v_o),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_i)
  );


  bsg_mux_width_p64_els_p8
  data_set_select_mux
  (
    .data_i(ld_data_tv_r),
    .sel_i({ n_11_net__2_, n_11_net__1_, n_11_net__0_ }),
    .data_o(ld_data_way_picked)
  );


  bsg_mux_butterfly_width_p64_els_p8
  write_mux_butterfly
  (
    .data_i(data_mem_pkt[511:0]),
    .sel_i(data_mem_pkt[515:513]),
    .data_o(data_mem_bank_data_li)
  );


  bsg_decode_num_out_p8
  lce_tag_mem_way_decode
  (
    .i(tag_mem_pkt[16:14]),
    .o(lce_tag_mem_way_one_hot)
  );

  assign N56 = N54 & N55;
  assign N57 = tag_mem_pkt[1] | N55;
  assign N59 = N54 | tag_mem_pkt[0];
  assign N61 = tag_mem_pkt[1] & tag_mem_pkt[0];

  bsg_lru_pseudo_tree_decode_ways_p8
  lru_decode
  (
    .way_id_i(hit_index),
    .data_o(lru_decode_data_lo),
    .mask_o(lru_decode_mask_lo)
  );


  bsg_mux_butterfly_width_p64_els_p8
  read_mux_butterfly
  (
    .data_i(data_mem_bank_data_lo),
    .sel_i(data_mem_pkt_way_r),
    .data_o(data_mem_data_li)
  );

  assign N65 = state_tv_r[14] | state_tv_r[15];
  assign N66 = state_tv_r[12] | state_tv_r[13];
  assign N67 = state_tv_r[10] | state_tv_r[11];
  assign N68 = state_tv_r[8] | state_tv_r[9];
  assign N69 = state_tv_r[6] | state_tv_r[7];
  assign N70 = state_tv_r[4] | state_tv_r[5];
  assign N71 = state_tv_r[2] | state_tv_r[3];
  assign N72 = state_tv_r[0] | state_tv_r[1];
  assign N73 = state_tv_r[14] | state_tv_r[15];
  assign N74 = state_tv_r[12] | state_tv_r[13];
  assign N75 = state_tv_r[10] | state_tv_r[11];
  assign N76 = state_tv_r[8] | state_tv_r[9];
  assign N77 = state_tv_r[6] | state_tv_r[7];
  assign N78 = state_tv_r[4] | state_tv_r[5];
  assign N79 = state_tv_r[2] | state_tv_r[3];
  assign N80 = state_tv_r[0] | state_tv_r[1];
  assign N18 = (N0)? 1'b0 :
               (N1)? tl_we : 1'b0;
  assign N0 = N17;
  assign N1 = N16;
  assign N19 = (N0)? 1'b0 :
               (N1)? tl_we : 1'b0;
  assign N22 = (N2)? 1'b0 :
               (N3)? tv_we : 1'b0;
  assign N2 = N21;
  assign N3 = N20;
  assign { N29, N28, N27, N26, N25, N24, N23 } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                 (N3)? { tv_we, tv_we, tv_we, tv_we, tv_we, tv_we, tv_we } : 1'b0;
  assign lru_way_li = (N4)? way_invalid_index :
                      (N5)? lru_encode : 1'b0;
  assign N4 = invalid_exist;
  assign N5 = N38;
  assign icache_pc_gen_data_o[95:64] = (N6)? ld_data_way_picked[63:32] :
                                       (N7)? ld_data_way_picked[31:0] : 1'b0;
  assign N6 = N40;
  assign N7 = N39;
  assign data_mem_bank_v_li = (N8)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } :
                              (N9)? { data_mem_pkt_yumi_li, data_mem_pkt_yumi_li, data_mem_pkt_yumi_li, data_mem_pkt_yumi_li, data_mem_pkt_yumi_li, data_mem_pkt_yumi_li, data_mem_pkt_yumi_li, data_mem_pkt_yumi_li } : 1'b0;
  assign N8 = tl_we;
  assign N9 = N41;
  assign data_mem_bank_addr_li[8:0] = (N8)? pc_gen_icache_vaddr_i[11:3] :
                                      (N9)? data_mem_pkt[521:513] : 1'b0;
  assign data_mem_bank_addr_li[17:9] = (N8)? pc_gen_icache_vaddr_i[11:3] :
                                       (N9)? { data_mem_pkt[521:514], N42 } : 1'b0;
  assign data_mem_bank_addr_li[26:18] = (N8)? pc_gen_icache_vaddr_i[11:3] :
                                        (N9)? { data_mem_pkt[521:515], N43, data_mem_pkt[513:513] } : 1'b0;
  assign data_mem_bank_addr_li[35:27] = (N8)? pc_gen_icache_vaddr_i[11:3] :
                                        (N9)? { data_mem_pkt[521:515], N44, N45 } : 1'b0;
  assign data_mem_bank_addr_li[44:36] = (N8)? pc_gen_icache_vaddr_i[11:3] :
                                        (N9)? { data_mem_pkt[521:516], N46, data_mem_pkt[514:513] } : 1'b0;
  assign data_mem_bank_addr_li[53:45] = (N8)? pc_gen_icache_vaddr_i[11:3] :
                                        (N9)? { data_mem_pkt[521:516], N47, data_mem_pkt[514:514], N48 } : 1'b0;
  assign data_mem_bank_addr_li[62:54] = (N8)? pc_gen_icache_vaddr_i[11:3] :
                                        (N9)? { data_mem_pkt[521:516], N49, N50, data_mem_pkt[513:513] } : 1'b0;
  assign data_mem_bank_addr_li[71:63] = (N8)? pc_gen_icache_vaddr_i[11:3] :
                                        (N9)? { data_mem_pkt[521:516], N51, N52, N53 } : 1'b0;
  assign tag_mem_addr_li = (N8)? pc_gen_icache_vaddr_i[11:6] :
                           (N9)? tag_mem_pkt[22:17] : 1'b0;
  assign tag_mem_w_mask_li = (N10)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } :
                             (N11)? { lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                             (N12)? { lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0] } :
                             (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = N56;
  assign N11 = N58;
  assign N12 = N60;
  assign N13 = N61;
  assign tag_mem_data_li = (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                           (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                           (N12)? { tag_mem_pkt[13:2], tag_mem_pkt[13:2], tag_mem_pkt[13:2], tag_mem_pkt[13:2], tag_mem_pkt[13:2], tag_mem_pkt[13:2], tag_mem_pkt[13:2], tag_mem_pkt[13:2] } :
                           (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign metadata_mem_w_li = (N14)? N63 :
                             (N15)? metadata_mem_pkt_yumi_li : 1'b0;
  assign N14 = v_tv_r;
  assign N15 = N62;
  assign metadata_mem_addr_li = (N14)? addr_tv_r[11:6] :
                                (N15)? metadata_mem_pkt[9:4] : 1'b0;
  assign metadata_mem_data_li = (N14)? lru_decode_data_lo :
                                (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign metadata_mem_mask_li = (N14)? lru_decode_mask_lo :
                                (N15)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign tl_we = N81 & N82;
  assign N81 = pc_gen_icache_vaddr_v_i & pc_gen_icache_vaddr_ready_o;
  assign N82 = ~poison_i;
  assign N16 = ~reset_i;
  assign N17 = reset_i;
  assign n_0_net_ = N83 & tag_mem_v_li;
  assign N83 = ~reset_i;
  assign n_1_net_ = N84 & data_mem_bank_v_li[0];
  assign N84 = ~reset_i;
  assign n_2_net_ = N85 & data_mem_bank_v_li[1];
  assign N85 = ~reset_i;
  assign n_3_net_ = N86 & data_mem_bank_v_li[2];
  assign N86 = ~reset_i;
  assign n_4_net_ = N87 & data_mem_bank_v_li[3];
  assign N87 = ~reset_i;
  assign n_5_net_ = N88 & data_mem_bank_v_li[4];
  assign N88 = ~reset_i;
  assign n_6_net_ = N89 & data_mem_bank_v_li[5];
  assign N89 = ~reset_i;
  assign n_7_net_ = N90 & data_mem_bank_v_li[6];
  assign N90 = ~reset_i;
  assign n_8_net_ = N91 & data_mem_bank_v_li[7];
  assign N91 = ~reset_i;
  assign tv_we = N92 & itlb_icache_data_resp_v_i;
  assign N92 = itlb_icache_data_resp_ready_o & N82;
  assign N20 = ~reset_i;
  assign N21 = reset_i;
  assign hit_v[0] = N30 & N72;
  assign hit_v[1] = N31 & N71;
  assign hit_v[2] = N32 & N70;
  assign hit_v[3] = N33 & N69;
  assign hit_v[4] = N34 & N68;
  assign hit_v[5] = N35 & N67;
  assign hit_v[6] = N36 & N66;
  assign hit_v[7] = N37 & N65;
  assign miss_v = N93 & v_tv_r;
  assign N93 = ~hit;
  assign n_9_net_ = N94 & metadata_mem_v_li;
  assign N94 = ~reset_i;
  assign n_10_net__7_ = ~N73;
  assign n_10_net__6_ = ~N74;
  assign n_10_net__5_ = ~N75;
  assign n_10_net__4_ = ~N76;
  assign n_10_net__3_ = ~N77;
  assign n_10_net__2_ = ~N78;
  assign n_10_net__1_ = ~N79;
  assign n_10_net__0_ = ~N80;
  assign N38 = ~invalid_exist;
  assign icache_pc_gen_data_v_o = N96 & N97;
  assign N96 = v_tv_r & N95;
  assign N95 = ~miss_v;
  assign N97 = ~reset_i;
  assign n_11_net__2_ = hit_index[2] ^ addr_tv_r[5];
  assign n_11_net__1_ = hit_index[1] ^ addr_tv_r[4];
  assign n_11_net__0_ = hit_index[0] ^ addr_tv_r[3];
  assign N39 = ~addr_tv_r[2];
  assign N40 = addr_tv_r[2];
  assign N41 = ~tl_we;
  assign data_mem_bank_w_li[7] = data_mem_pkt_yumi_li & data_mem_pkt[512];
  assign data_mem_bank_w_li[6] = data_mem_pkt_yumi_li & data_mem_pkt[512];
  assign data_mem_bank_w_li[5] = data_mem_pkt_yumi_li & data_mem_pkt[512];
  assign data_mem_bank_w_li[4] = data_mem_pkt_yumi_li & data_mem_pkt[512];
  assign data_mem_bank_w_li[3] = data_mem_pkt_yumi_li & data_mem_pkt[512];
  assign data_mem_bank_w_li[2] = data_mem_pkt_yumi_li & data_mem_pkt[512];
  assign data_mem_bank_w_li[1] = data_mem_pkt_yumi_li & data_mem_pkt[512];
  assign data_mem_bank_w_li[0] = data_mem_pkt_yumi_li & data_mem_pkt[512];
  assign N42 = ~data_mem_pkt[513];
  assign N43 = ~data_mem_pkt[514];
  assign N44 = ~data_mem_pkt[514];
  assign N45 = ~data_mem_pkt[513];
  assign N46 = ~data_mem_pkt[515];
  assign N47 = ~data_mem_pkt[515];
  assign N48 = ~data_mem_pkt[513];
  assign N49 = ~data_mem_pkt[515];
  assign N50 = ~data_mem_pkt[514];
  assign N51 = ~data_mem_pkt[515];
  assign N52 = ~data_mem_pkt[514];
  assign N53 = ~data_mem_pkt[513];
  assign tag_mem_v_li = tl_we | tag_mem_pkt_yumi_li;
  assign tag_mem_w_li = N41 & tag_mem_pkt_v_lo;
  assign N54 = ~tag_mem_pkt[1];
  assign N55 = ~tag_mem_pkt[0];
  assign N58 = ~N57;
  assign N60 = ~N59;
  assign metadata_mem_v_li = v_tv_r | metadata_mem_pkt_yumi_li;
  assign N62 = ~v_tv_r;
  assign N63 = ~miss_v;
  assign N64 = data_mem_pkt_yumi_li & N98;
  assign N98 = ~data_mem_pkt[512];
  assign data_mem_pkt_yumi_li = data_mem_pkt_v_lo & N41;
  assign tag_mem_pkt_yumi_li = tag_mem_pkt_v_lo & N41;
  assign metadata_mem_pkt_yumi_li = N62 & metadata_mem_pkt_v_lo;

  always @(posedge clk_i) begin
    if(N19) begin
      { vaddr_tl_r[11:0] } <= { pc_gen_icache_vaddr_i[11:0] };
      { eaddr_tl_r[63:0] } <= { pc_gen_icache_vaddr_i[63:0] };
    end
    if(1'b1) begin
      itlb_icache_data_resp_ready_o <= N18;
      v_tv_r <= N22;
    end
    if(N28) begin
      { state_tv_r[15:0] } <= { tag_mem_data_lo[95:94], tag_mem_data_lo[83:82], tag_mem_data_lo[71:70], tag_mem_data_lo[59:58], tag_mem_data_lo[47:46], tag_mem_data_lo[35:34], tag_mem_data_lo[23:22], tag_mem_data_lo[11:10] };
      { ld_data_tv_r[16:0] } <= { data_mem_bank_data_lo[16:0] };
      { addr_tv_r[5:5] } <= { vaddr_tl_r[5:5] };
      { tag_tv_r[79:14] } <= { tag_mem_data_lo[93:84], tag_mem_data_lo[81:72], tag_mem_data_lo[69:60], tag_mem_data_lo[57:48], tag_mem_data_lo[45:36], tag_mem_data_lo[33:24], tag_mem_data_lo[21:16] };
    end
    if(N23) begin
      { ld_data_tv_r[511:413] } <= { data_mem_bank_data_lo[511:413] };
      { addr_tv_r[0:0] } <= { vaddr_tl_r[0:0] };
    end
    if(N24) begin
      { ld_data_tv_r[412:314] } <= { data_mem_bank_data_lo[412:314] };
      { addr_tv_r[1:1] } <= { vaddr_tl_r[1:1] };
    end
    if(N25) begin
      { ld_data_tv_r[313:215] } <= { data_mem_bank_data_lo[313:215] };
      { addr_tv_r[2:2] } <= { vaddr_tl_r[2:2] };
    end
    if(N26) begin
      { ld_data_tv_r[214:116] } <= { data_mem_bank_data_lo[214:116] };
      { addr_tv_r[3:3] } <= { vaddr_tl_r[3:3] };
    end
    if(N27) begin
      { ld_data_tv_r[115:17] } <= { data_mem_bank_data_lo[115:17] };
      { addr_tv_r[4:4] } <= { vaddr_tl_r[4:4] };
    end
    if(N29) begin
      { addr_tv_r[21:6] } <= { itlb_icache_data_resp_i[9:0], vaddr_tl_r[11:6] };
      { icache_pc_gen_data_o[63:0] } <= { eaddr_tl_r[63:0] };
      { tag_tv_r[13:0] } <= { tag_mem_data_lo[15:12], tag_mem_data_lo[9:0] };
    end
    if(N64) begin
      { data_mem_pkt_way_r[2:0] } <= { data_mem_pkt[515:513] };
    end
  end


endmodule



module itlb_vaddr_width_p39_paddr_width_p22_eaddr_width_p64_tag_width_p10_btb_indx_width_p9_bht_indx_width_p5_ras_addr_width_p22_asid_width_p10_ppn_start_bit_p12
(
  clk_i,
  reset_i,
  fe_itlb_i,
  fe_itlb_v_i,
  fe_itlb_ready_o,
  pc_gen_itlb_i,
  pc_gen_itlb_v_i,
  pc_gen_itlb_ready_o,
  itlb_icache_o,
  itlb_icache_data_resp_v_o,
  itlb_icache_data_resp_ready_i,
  itlb_fe_o,
  itlb_fe_v_o,
  itlb_fe_ready_i
);

  input [108:0] fe_itlb_i;
  input [63:0] pc_gen_itlb_i;
  output [9:0] itlb_icache_o;
  output [133:0] itlb_fe_o;
  input clk_i;
  input reset_i;
  input fe_itlb_v_i;
  input pc_gen_itlb_v_i;
  input itlb_icache_data_resp_ready_i;
  input itlb_fe_ready_i;
  output fe_itlb_ready_o;
  output pc_gen_itlb_ready_o;
  output itlb_icache_data_resp_v_o;
  output itlb_fe_v_o;
  wire [133:0] itlb_fe_o;
  wire fe_itlb_ready_o,pc_gen_itlb_ready_o,itlb_icache_data_resp_v_o,itlb_fe_v_o;
  reg [9:0] itlb_icache_o;
  assign pc_gen_itlb_ready_o = 1'b1;
  assign itlb_icache_data_resp_v_o = 1'b1;
  assign fe_itlb_ready_o = 1'b0;
  assign itlb_fe_v_o = 1'b0;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { itlb_icache_o[9:0] } <= { pc_gen_itlb_i[21:12] };
    end
  end


endmodule



module bp_fe_top_39_22_1_2_8_64_64_9_5_22_10_80000124
(
  clk_i,
  reset_i,
  icache_id_i,
  fe_cmd_i,
  fe_cmd_v_i,
  fe_cmd_ready_o,
  fe_queue_o,
  fe_queue_v_o,
  fe_queue_ready_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i
);

  input [0:0] icache_id_i;
  input [108:0] fe_cmd_i;
  output [133:0] fe_queue_o;
  output [96:0] lce_req_o;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  input [35:0] lce_cmd_i;
  input [517:0] lce_data_cmd_i;
  output [517:0] lce_data_cmd_o;
  input clk_i;
  input reset_i;
  input fe_cmd_v_i;
  input fe_queue_ready_i;
  input lce_req_ready_i;
  input lce_resp_ready_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_v_i;
  input lce_data_cmd_ready_i;
  output fe_cmd_ready_o;
  output fe_queue_v_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_ready_o;
  output lce_data_cmd_ready_o;
  output lce_data_cmd_v_o;
  wire [133:0] fe_queue_o,itlb_fe_queue;
  wire [96:0] lce_req_o;
  wire [25:0] lce_resp_o;
  wire [536:0] lce_data_resp_o;
  wire [517:0] lce_data_cmd_o;
  wire fe_cmd_ready_o,fe_queue_v_o,lce_req_v_o,lce_resp_v_o,lce_data_resp_v_o,
  lce_cmd_ready_o,lce_data_cmd_ready_o,lce_data_cmd_v_o,N0,N1,pc_gen_queue_scan_instr__68_,
  pc_gen_queue_scan_instr__67_,pc_gen_queue_scan_instr__66_,
  pc_gen_queue_scan_instr__65_,pc_gen_queue_scan_instr__64_,pc_gen_queue_scan_instr__63_,
  pc_gen_queue_scan_instr__62_,pc_gen_queue_scan_instr__61_,pc_gen_queue_scan_instr__60_,
  pc_gen_queue_scan_instr__59_,pc_gen_queue_scan_instr__58_,pc_gen_queue_scan_instr__57_,
  pc_gen_queue_scan_instr__56_,pc_gen_queue_scan_instr__55_,
  pc_gen_queue_scan_instr__54_,pc_gen_queue_scan_instr__53_,pc_gen_queue_scan_instr__52_,
  pc_gen_queue_scan_instr__51_,pc_gen_queue_scan_instr__50_,pc_gen_queue_scan_instr__49_,
  pc_gen_queue_scan_instr__48_,pc_gen_queue_scan_instr__47_,pc_gen_queue_scan_instr__46_,
  pc_gen_queue_scan_instr__45_,pc_gen_queue_scan_instr__44_,
  pc_gen_queue_scan_instr__43_,pc_gen_queue_scan_instr__42_,pc_gen_queue_scan_instr__41_,
  pc_gen_queue_scan_instr__40_,pc_gen_queue_scan_instr__39_,pc_gen_queue_scan_instr__38_,
  pc_gen_queue_scan_instr__37_,pc_gen_queue_scan_instr__36_,pc_gen_queue_scan_instr__35_,
  pc_gen_queue_scan_instr__34_,pc_gen_queue_scan_instr__33_,
  pc_gen_queue_scan_instr__32_,pc_gen_queue_scan_instr__31_,pc_gen_queue_scan_instr__30_,
  pc_gen_queue_scan_instr__29_,pc_gen_queue_scan_instr__28_,pc_gen_queue_scan_instr__27_,
  pc_gen_queue_scan_instr__26_,pc_gen_queue_scan_instr__25_,pc_gen_queue_scan_instr__24_,
  pc_gen_queue_scan_instr__23_,pc_gen_queue_scan_instr__22_,
  pc_gen_queue_scan_instr__21_,pc_gen_queue_scan_instr__20_,pc_gen_queue_scan_instr__19_,
  pc_gen_queue_scan_instr__18_,pc_gen_queue_scan_instr__17_,pc_gen_queue_scan_instr__16_,
  pc_gen_queue_scan_instr__15_,pc_gen_queue_scan_instr__14_,pc_gen_queue_scan_instr__13_,
  pc_gen_queue_scan_instr__12_,pc_gen_queue_scan_instr__11_,
  pc_gen_queue_scan_instr__10_,pc_gen_queue_scan_instr__9_,pc_gen_queue_scan_instr__8_,
  pc_gen_queue_scan_instr__7_,pc_gen_queue_scan_instr__6_,pc_gen_queue_scan_instr__5_,
  pc_gen_queue_scan_instr__4_,pc_gen_queue_scan_instr__3_,pc_gen_queue_scan_instr__2_,
  pc_gen_queue_scan_instr__1_,pc_gen_queue_scan_instr__0_,fe_pc_gen_branch_metadata_fwd__35_,
  fe_pc_gen_branch_metadata_fwd__34_,fe_pc_gen_branch_metadata_fwd__33_,
  fe_pc_gen_branch_metadata_fwd__32_,fe_pc_gen_branch_metadata_fwd__31_,
  fe_pc_gen_branch_metadata_fwd__30_,fe_pc_gen_branch_metadata_fwd__29_,
  fe_pc_gen_branch_metadata_fwd__28_,fe_pc_gen_branch_metadata_fwd__27_,fe_pc_gen_branch_metadata_fwd__26_,
  fe_pc_gen_branch_metadata_fwd__25_,fe_pc_gen_branch_metadata_fwd__24_,
  fe_pc_gen_branch_metadata_fwd__23_,fe_pc_gen_branch_metadata_fwd__22_,
  fe_pc_gen_branch_metadata_fwd__21_,fe_pc_gen_branch_metadata_fwd__20_,fe_pc_gen_branch_metadata_fwd__19_,
  fe_pc_gen_branch_metadata_fwd__18_,fe_pc_gen_branch_metadata_fwd__17_,
  fe_pc_gen_branch_metadata_fwd__16_,fe_pc_gen_branch_metadata_fwd__15_,
  fe_pc_gen_branch_metadata_fwd__14_,fe_pc_gen_branch_metadata_fwd__13_,
  fe_pc_gen_branch_metadata_fwd__12_,fe_pc_gen_branch_metadata_fwd__11_,fe_pc_gen_branch_metadata_fwd__10_,
  fe_pc_gen_branch_metadata_fwd__9_,fe_pc_gen_branch_metadata_fwd__8_,
  fe_pc_gen_branch_metadata_fwd__7_,fe_pc_gen_branch_metadata_fwd__6_,
  fe_pc_gen_branch_metadata_fwd__5_,fe_pc_gen_branch_metadata_fwd__4_,fe_pc_gen_branch_metadata_fwd__3_,
  fe_pc_gen_branch_metadata_fwd__2_,fe_pc_gen_branch_metadata_fwd__1_,
  fe_pc_gen_branch_metadata_fwd__0_,fe_pc_gen_pc_redirect_valid_,N2,N3,cache_miss,poison,
  pc_gen_icache_v,pc_gen_icache_ready,icache_pc_gen_v,icache_pc_gen_ready,pc_gen_itlb_v,
  pc_gen_itlb_ready,itlb_icache_data_resp_v,itlb_icache_data_resp_ready,fe_itlb_ready,
  itlb_fe_v,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,
  N24,N25,N26,N27,N28;
  wire [63:0] pc_gen_icache,pc_gen_itlb;
  wire [95:0] icache_pc_gen;
  wire [9:0] itlb_icache;

  bp_fe_pc_gen_39_22_64_9_5_22_32_10_80000124_1
  bp_fe_pc_gen_1
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(1'b1),
    .pc_gen_icache_o(pc_gen_icache),
    .pc_gen_icache_v_o(pc_gen_icache_v),
    .pc_gen_icache_ready_i(pc_gen_icache_ready),
    .icache_pc_gen_i(icache_pc_gen),
    .icache_pc_gen_v_i(icache_pc_gen_v),
    .icache_pc_gen_ready_o(icache_pc_gen_ready),
    .icache_miss_i(cache_miss),
    .pc_gen_itlb_o(pc_gen_itlb),
    .pc_gen_itlb_v_o(pc_gen_itlb_v),
    .pc_gen_itlb_ready_i(pc_gen_itlb_ready),
    .pc_gen_fe_o({ fe_queue_o[133:133], pc_gen_queue_scan_instr__68_, pc_gen_queue_scan_instr__67_, pc_gen_queue_scan_instr__66_, pc_gen_queue_scan_instr__65_, pc_gen_queue_scan_instr__64_, pc_gen_queue_scan_instr__63_, pc_gen_queue_scan_instr__62_, pc_gen_queue_scan_instr__61_, pc_gen_queue_scan_instr__60_, pc_gen_queue_scan_instr__59_, pc_gen_queue_scan_instr__58_, pc_gen_queue_scan_instr__57_, pc_gen_queue_scan_instr__56_, pc_gen_queue_scan_instr__55_, pc_gen_queue_scan_instr__54_, pc_gen_queue_scan_instr__53_, pc_gen_queue_scan_instr__52_, pc_gen_queue_scan_instr__51_, pc_gen_queue_scan_instr__50_, pc_gen_queue_scan_instr__49_, pc_gen_queue_scan_instr__48_, pc_gen_queue_scan_instr__47_, pc_gen_queue_scan_instr__46_, pc_gen_queue_scan_instr__45_, pc_gen_queue_scan_instr__44_, pc_gen_queue_scan_instr__43_, pc_gen_queue_scan_instr__42_, pc_gen_queue_scan_instr__41_, pc_gen_queue_scan_instr__40_, pc_gen_queue_scan_instr__39_, pc_gen_queue_scan_instr__38_, pc_gen_queue_scan_instr__37_, pc_gen_queue_scan_instr__36_, pc_gen_queue_scan_instr__35_, pc_gen_queue_scan_instr__34_, pc_gen_queue_scan_instr__33_, pc_gen_queue_scan_instr__32_, pc_gen_queue_scan_instr__31_, pc_gen_queue_scan_instr__30_, pc_gen_queue_scan_instr__29_, pc_gen_queue_scan_instr__28_, pc_gen_queue_scan_instr__27_, pc_gen_queue_scan_instr__26_, pc_gen_queue_scan_instr__25_, pc_gen_queue_scan_instr__24_, pc_gen_queue_scan_instr__23_, pc_gen_queue_scan_instr__22_, pc_gen_queue_scan_instr__21_, pc_gen_queue_scan_instr__20_, pc_gen_queue_scan_instr__19_, pc_gen_queue_scan_instr__18_, pc_gen_queue_scan_instr__17_, pc_gen_queue_scan_instr__16_, pc_gen_queue_scan_instr__15_, pc_gen_queue_scan_instr__14_, pc_gen_queue_scan_instr__13_, pc_gen_queue_scan_instr__12_, pc_gen_queue_scan_instr__11_, pc_gen_queue_scan_instr__10_, pc_gen_queue_scan_instr__9_, pc_gen_queue_scan_instr__8_, pc_gen_queue_scan_instr__7_, pc_gen_queue_scan_instr__6_, pc_gen_queue_scan_instr__5_, pc_gen_queue_scan_instr__4_, pc_gen_queue_scan_instr__3_, pc_gen_queue_scan_instr__2_, pc_gen_queue_scan_instr__1_, pc_gen_queue_scan_instr__0_, fe_queue_o[132:0] }),
    .pc_gen_fe_v_o(fe_queue_v_o),
    .pc_gen_fe_ready_i(fe_queue_ready_i),
    .fe_pc_gen_i({ fe_cmd_i[105:42], fe_pc_gen_branch_metadata_fwd__35_, fe_pc_gen_branch_metadata_fwd__34_, fe_pc_gen_branch_metadata_fwd__33_, fe_pc_gen_branch_metadata_fwd__32_, fe_pc_gen_branch_metadata_fwd__31_, fe_pc_gen_branch_metadata_fwd__30_, fe_pc_gen_branch_metadata_fwd__29_, fe_pc_gen_branch_metadata_fwd__28_, fe_pc_gen_branch_metadata_fwd__27_, fe_pc_gen_branch_metadata_fwd__26_, fe_pc_gen_branch_metadata_fwd__25_, fe_pc_gen_branch_metadata_fwd__24_, fe_pc_gen_branch_metadata_fwd__23_, fe_pc_gen_branch_metadata_fwd__22_, fe_pc_gen_branch_metadata_fwd__21_, fe_pc_gen_branch_metadata_fwd__20_, fe_pc_gen_branch_metadata_fwd__19_, fe_pc_gen_branch_metadata_fwd__18_, fe_pc_gen_branch_metadata_fwd__17_, fe_pc_gen_branch_metadata_fwd__16_, fe_pc_gen_branch_metadata_fwd__15_, fe_pc_gen_branch_metadata_fwd__14_, fe_pc_gen_branch_metadata_fwd__13_, fe_pc_gen_branch_metadata_fwd__12_, fe_pc_gen_branch_metadata_fwd__11_, fe_pc_gen_branch_metadata_fwd__10_, fe_pc_gen_branch_metadata_fwd__9_, fe_pc_gen_branch_metadata_fwd__8_, fe_pc_gen_branch_metadata_fwd__7_, fe_pc_gen_branch_metadata_fwd__6_, fe_pc_gen_branch_metadata_fwd__5_, fe_pc_gen_branch_metadata_fwd__4_, fe_pc_gen_branch_metadata_fwd__3_, fe_pc_gen_branch_metadata_fwd__2_, fe_pc_gen_branch_metadata_fwd__1_, fe_pc_gen_branch_metadata_fwd__0_, fe_pc_gen_pc_redirect_valid_, N7 }),
    .fe_pc_gen_v_i(fe_cmd_v_i),
    .fe_pc_gen_ready_o(fe_cmd_ready_o)
  );


  icache_eaddr_width_p64_paddr_width_p22_data_width_p64_instr_width_p32_num_cce_p1_num_lce_p2_ways_p8_sets_p64
  icache_1
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .id_i(icache_id_i[0]),
    .pc_gen_icache_vaddr_i(pc_gen_icache),
    .pc_gen_icache_vaddr_v_i(pc_gen_icache_v),
    .pc_gen_icache_vaddr_ready_o(pc_gen_icache_ready),
    .icache_pc_gen_data_o(icache_pc_gen),
    .icache_pc_gen_data_v_o(icache_pc_gen_v),
    .icache_pc_gen_data_ready_i(icache_pc_gen_ready),
    .itlb_icache_data_resp_i(itlb_icache),
    .itlb_icache_data_resp_v_i(itlb_icache_data_resp_v),
    .itlb_icache_data_resp_ready_o(itlb_icache_data_resp_ready),
    .cache_miss_o(cache_miss),
    .poison_i(poison),
    .lce_req_o(lce_req_o),
    .lce_req_v_o(lce_req_v_o),
    .lce_req_ready_i(lce_req_ready_i),
    .lce_resp_o(lce_resp_o),
    .lce_resp_v_o(lce_resp_v_o),
    .lce_resp_ready_i(lce_resp_ready_i),
    .lce_data_resp_o(lce_data_resp_o),
    .lce_data_resp_v_o(lce_data_resp_v_o),
    .lce_data_resp_ready_i(lce_data_resp_ready_i),
    .lce_cmd_i(lce_cmd_i),
    .lce_cmd_v_i(lce_cmd_v_i),
    .lce_cmd_ready_o(lce_cmd_ready_o),
    .lce_data_cmd_i(lce_data_cmd_i),
    .lce_data_cmd_v_i(lce_data_cmd_v_i),
    .lce_data_cmd_ready_o(lce_data_cmd_ready_o),
    .lce_data_cmd_o(lce_data_cmd_o),
    .lce_data_cmd_v_o(lce_data_cmd_v_o),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_i)
  );


  itlb_vaddr_width_p39_paddr_width_p22_eaddr_width_p64_tag_width_p10_btb_indx_width_p9_bht_indx_width_p5_ras_addr_width_p22_asid_width_p10_ppn_start_bit_p12
  itlb_1
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .fe_itlb_i(fe_cmd_i),
    .fe_itlb_v_i(fe_cmd_v_i),
    .fe_itlb_ready_o(fe_itlb_ready),
    .pc_gen_itlb_i(pc_gen_itlb),
    .pc_gen_itlb_v_i(pc_gen_itlb_v),
    .pc_gen_itlb_ready_o(pc_gen_itlb_ready),
    .itlb_icache_o(itlb_icache),
    .itlb_icache_data_resp_v_o(itlb_icache_data_resp_v),
    .itlb_icache_data_resp_ready_i(itlb_icache_data_resp_ready),
    .itlb_fe_o(itlb_fe_queue),
    .itlb_fe_v_o(itlb_fe_v),
    .itlb_fe_ready_i(fe_queue_ready_i)
  );

  assign N4 = ~fe_cmd_i[108];
  assign N5 = fe_cmd_i[107] | N4;
  assign N6 = fe_cmd_i[106] | N5;
  assign N7 = ~N6;
  assign N8 = ~fe_cmd_i[106];
  assign N9 = fe_cmd_i[107] | fe_cmd_i[108];
  assign N10 = N8 | N9;
  assign N11 = ~N10;
  assign N12 = ~fe_cmd_i[41];
  assign N13 = fe_cmd_i[40] | N12;
  assign N14 = fe_cmd_i[39] | N13;
  assign N15 = ~N14;
  assign N16 = ~fe_cmd_i[107];
  assign N17 = ~fe_cmd_i[106];
  assign N18 = N16 | fe_cmd_i[108];
  assign N19 = N17 | N18;
  assign N20 = ~N19;
  assign N21 = ~fe_cmd_i[106];
  assign N22 = fe_cmd_i[107] | fe_cmd_i[108];
  assign N23 = N21 | N22;
  assign N24 = ~N23;
  assign N25 = ~fe_cmd_i[108];
  assign N26 = fe_cmd_i[107] | N25;
  assign N27 = fe_cmd_i[106] | N26;
  assign N28 = ~N27;
  assign { fe_pc_gen_branch_metadata_fwd__35_, fe_pc_gen_branch_metadata_fwd__34_, fe_pc_gen_branch_metadata_fwd__33_, fe_pc_gen_branch_metadata_fwd__32_, fe_pc_gen_branch_metadata_fwd__31_, fe_pc_gen_branch_metadata_fwd__30_, fe_pc_gen_branch_metadata_fwd__29_, fe_pc_gen_branch_metadata_fwd__28_, fe_pc_gen_branch_metadata_fwd__27_, fe_pc_gen_branch_metadata_fwd__26_, fe_pc_gen_branch_metadata_fwd__25_, fe_pc_gen_branch_metadata_fwd__24_, fe_pc_gen_branch_metadata_fwd__23_, fe_pc_gen_branch_metadata_fwd__22_, fe_pc_gen_branch_metadata_fwd__21_, fe_pc_gen_branch_metadata_fwd__20_, fe_pc_gen_branch_metadata_fwd__19_, fe_pc_gen_branch_metadata_fwd__18_, fe_pc_gen_branch_metadata_fwd__17_, fe_pc_gen_branch_metadata_fwd__16_, fe_pc_gen_branch_metadata_fwd__15_, fe_pc_gen_branch_metadata_fwd__14_, fe_pc_gen_branch_metadata_fwd__13_, fe_pc_gen_branch_metadata_fwd__12_, fe_pc_gen_branch_metadata_fwd__11_, fe_pc_gen_branch_metadata_fwd__10_, fe_pc_gen_branch_metadata_fwd__9_, fe_pc_gen_branch_metadata_fwd__8_, fe_pc_gen_branch_metadata_fwd__7_, fe_pc_gen_branch_metadata_fwd__6_, fe_pc_gen_branch_metadata_fwd__5_, fe_pc_gen_branch_metadata_fwd__4_, fe_pc_gen_branch_metadata_fwd__3_, fe_pc_gen_branch_metadata_fwd__2_, fe_pc_gen_branch_metadata_fwd__1_, fe_pc_gen_branch_metadata_fwd__0_ } = (N0)? fe_cmd_i[41:6] :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N1)? fe_cmd_i[38:3] :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N28;
  assign N1 = N24;
  assign fe_pc_gen_pc_redirect_valid_ = N11 & N15;
  assign N2 = N24 | N28;
  assign N3 = ~N2;
  assign poison = cache_miss & N20;

endmodule



module bsg_circular_ptr_slots_p16_max_add_p1
(
  clk,
  reset_i,
  add_i,
  o
);

  input [0:0] add_i;
  output [3:0] o;
  input clk;
  input reset_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9;
  wire [3:0] genblk1_genblk1_ptr_r_p1;
  reg [3:0] o;
  assign genblk1_genblk1_ptr_r_p1 = o + 1'b1;
  assign { N6, N5, N4, N3 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0 } :
                              (N1)? genblk1_genblk1_ptr_r_p1 : 1'b0;
  assign N0 = reset_i;
  assign N1 = N2;
  assign N2 = ~reset_i;
  assign N7 = ~add_i[0];
  assign N8 = N7 & N2;
  assign N9 = ~N8;

  always @(posedge clk) begin
    if(N9) begin
      { o[3:0] } <= { N6, N5, N4, N3 };
    end
  end


endmodule



module bsg_circular_ptr_slots_p16_max_add_p15
(
  clk,
  reset_i,
  add_i,
  o
);

  input [3:0] add_i;
  output [3:0] o;
  input clk;
  input reset_i;
  wire N0,N1,N2,N3,N4,N5,N6;
  wire [3:0] ptr_n;
  reg [3:0] o;
  assign ptr_n = o + add_i;
  assign { N6, N5, N4, N3 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0 } :
                              (N1)? ptr_n : 1'b0;
  assign N0 = reset_i;
  assign N1 = N2;
  assign N2 = ~reset_i;

  always @(posedge clk) begin
    if(1'b1) begin
      { o[3:0] } <= { N6, N5, N4, N3 };
    end
  end


endmodule



module bsg_mem_p134
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [2:0] w_addr_i;
  input [133:0] w_data_i;
  input [2:0] r_addr_i;
  output [133:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [133:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53;
  reg [1071:0] mem;
  assign r_data_o[133] = (N17)? mem[133] :
                         (N19)? mem[267] :
                         (N21)? mem[401] :
                         (N23)? mem[535] :
                         (N18)? mem[669] :
                         (N20)? mem[803] :
                         (N22)? mem[937] :
                         (N24)? mem[1071] : 1'b0;
  assign r_data_o[132] = (N17)? mem[132] :
                         (N19)? mem[266] :
                         (N21)? mem[400] :
                         (N23)? mem[534] :
                         (N18)? mem[668] :
                         (N20)? mem[802] :
                         (N22)? mem[936] :
                         (N24)? mem[1070] : 1'b0;
  assign r_data_o[131] = (N17)? mem[131] :
                         (N19)? mem[265] :
                         (N21)? mem[399] :
                         (N23)? mem[533] :
                         (N18)? mem[667] :
                         (N20)? mem[801] :
                         (N22)? mem[935] :
                         (N24)? mem[1069] : 1'b0;
  assign r_data_o[130] = (N17)? mem[130] :
                         (N19)? mem[264] :
                         (N21)? mem[398] :
                         (N23)? mem[532] :
                         (N18)? mem[666] :
                         (N20)? mem[800] :
                         (N22)? mem[934] :
                         (N24)? mem[1068] : 1'b0;
  assign r_data_o[129] = (N17)? mem[129] :
                         (N19)? mem[263] :
                         (N21)? mem[397] :
                         (N23)? mem[531] :
                         (N18)? mem[665] :
                         (N20)? mem[799] :
                         (N22)? mem[933] :
                         (N24)? mem[1067] : 1'b0;
  assign r_data_o[128] = (N17)? mem[128] :
                         (N19)? mem[262] :
                         (N21)? mem[396] :
                         (N23)? mem[530] :
                         (N18)? mem[664] :
                         (N20)? mem[798] :
                         (N22)? mem[932] :
                         (N24)? mem[1066] : 1'b0;
  assign r_data_o[127] = (N17)? mem[127] :
                         (N19)? mem[261] :
                         (N21)? mem[395] :
                         (N23)? mem[529] :
                         (N18)? mem[663] :
                         (N20)? mem[797] :
                         (N22)? mem[931] :
                         (N24)? mem[1065] : 1'b0;
  assign r_data_o[126] = (N17)? mem[126] :
                         (N19)? mem[260] :
                         (N21)? mem[394] :
                         (N23)? mem[528] :
                         (N18)? mem[662] :
                         (N20)? mem[796] :
                         (N22)? mem[930] :
                         (N24)? mem[1064] : 1'b0;
  assign r_data_o[125] = (N17)? mem[125] :
                         (N19)? mem[259] :
                         (N21)? mem[393] :
                         (N23)? mem[527] :
                         (N18)? mem[661] :
                         (N20)? mem[795] :
                         (N22)? mem[929] :
                         (N24)? mem[1063] : 1'b0;
  assign r_data_o[124] = (N17)? mem[124] :
                         (N19)? mem[258] :
                         (N21)? mem[392] :
                         (N23)? mem[526] :
                         (N18)? mem[660] :
                         (N20)? mem[794] :
                         (N22)? mem[928] :
                         (N24)? mem[1062] : 1'b0;
  assign r_data_o[123] = (N17)? mem[123] :
                         (N19)? mem[257] :
                         (N21)? mem[391] :
                         (N23)? mem[525] :
                         (N18)? mem[659] :
                         (N20)? mem[793] :
                         (N22)? mem[927] :
                         (N24)? mem[1061] : 1'b0;
  assign r_data_o[122] = (N17)? mem[122] :
                         (N19)? mem[256] :
                         (N21)? mem[390] :
                         (N23)? mem[524] :
                         (N18)? mem[658] :
                         (N20)? mem[792] :
                         (N22)? mem[926] :
                         (N24)? mem[1060] : 1'b0;
  assign r_data_o[121] = (N17)? mem[121] :
                         (N19)? mem[255] :
                         (N21)? mem[389] :
                         (N23)? mem[523] :
                         (N18)? mem[657] :
                         (N20)? mem[791] :
                         (N22)? mem[925] :
                         (N24)? mem[1059] : 1'b0;
  assign r_data_o[120] = (N17)? mem[120] :
                         (N19)? mem[254] :
                         (N21)? mem[388] :
                         (N23)? mem[522] :
                         (N18)? mem[656] :
                         (N20)? mem[790] :
                         (N22)? mem[924] :
                         (N24)? mem[1058] : 1'b0;
  assign r_data_o[119] = (N17)? mem[119] :
                         (N19)? mem[253] :
                         (N21)? mem[387] :
                         (N23)? mem[521] :
                         (N18)? mem[655] :
                         (N20)? mem[789] :
                         (N22)? mem[923] :
                         (N24)? mem[1057] : 1'b0;
  assign r_data_o[118] = (N17)? mem[118] :
                         (N19)? mem[252] :
                         (N21)? mem[386] :
                         (N23)? mem[520] :
                         (N18)? mem[654] :
                         (N20)? mem[788] :
                         (N22)? mem[922] :
                         (N24)? mem[1056] : 1'b0;
  assign r_data_o[117] = (N17)? mem[117] :
                         (N19)? mem[251] :
                         (N21)? mem[385] :
                         (N23)? mem[519] :
                         (N18)? mem[653] :
                         (N20)? mem[787] :
                         (N22)? mem[921] :
                         (N24)? mem[1055] : 1'b0;
  assign r_data_o[116] = (N17)? mem[116] :
                         (N19)? mem[250] :
                         (N21)? mem[384] :
                         (N23)? mem[518] :
                         (N18)? mem[652] :
                         (N20)? mem[786] :
                         (N22)? mem[920] :
                         (N24)? mem[1054] : 1'b0;
  assign r_data_o[115] = (N17)? mem[115] :
                         (N19)? mem[249] :
                         (N21)? mem[383] :
                         (N23)? mem[517] :
                         (N18)? mem[651] :
                         (N20)? mem[785] :
                         (N22)? mem[919] :
                         (N24)? mem[1053] : 1'b0;
  assign r_data_o[114] = (N17)? mem[114] :
                         (N19)? mem[248] :
                         (N21)? mem[382] :
                         (N23)? mem[516] :
                         (N18)? mem[650] :
                         (N20)? mem[784] :
                         (N22)? mem[918] :
                         (N24)? mem[1052] : 1'b0;
  assign r_data_o[113] = (N17)? mem[113] :
                         (N19)? mem[247] :
                         (N21)? mem[381] :
                         (N23)? mem[515] :
                         (N18)? mem[649] :
                         (N20)? mem[783] :
                         (N22)? mem[917] :
                         (N24)? mem[1051] : 1'b0;
  assign r_data_o[112] = (N17)? mem[112] :
                         (N19)? mem[246] :
                         (N21)? mem[380] :
                         (N23)? mem[514] :
                         (N18)? mem[648] :
                         (N20)? mem[782] :
                         (N22)? mem[916] :
                         (N24)? mem[1050] : 1'b0;
  assign r_data_o[111] = (N17)? mem[111] :
                         (N19)? mem[245] :
                         (N21)? mem[379] :
                         (N23)? mem[513] :
                         (N18)? mem[647] :
                         (N20)? mem[781] :
                         (N22)? mem[915] :
                         (N24)? mem[1049] : 1'b0;
  assign r_data_o[110] = (N17)? mem[110] :
                         (N19)? mem[244] :
                         (N21)? mem[378] :
                         (N23)? mem[512] :
                         (N18)? mem[646] :
                         (N20)? mem[780] :
                         (N22)? mem[914] :
                         (N24)? mem[1048] : 1'b0;
  assign r_data_o[109] = (N17)? mem[109] :
                         (N19)? mem[243] :
                         (N21)? mem[377] :
                         (N23)? mem[511] :
                         (N18)? mem[645] :
                         (N20)? mem[779] :
                         (N22)? mem[913] :
                         (N24)? mem[1047] : 1'b0;
  assign r_data_o[108] = (N17)? mem[108] :
                         (N19)? mem[242] :
                         (N21)? mem[376] :
                         (N23)? mem[510] :
                         (N18)? mem[644] :
                         (N20)? mem[778] :
                         (N22)? mem[912] :
                         (N24)? mem[1046] : 1'b0;
  assign r_data_o[107] = (N17)? mem[107] :
                         (N19)? mem[241] :
                         (N21)? mem[375] :
                         (N23)? mem[509] :
                         (N18)? mem[643] :
                         (N20)? mem[777] :
                         (N22)? mem[911] :
                         (N24)? mem[1045] : 1'b0;
  assign r_data_o[106] = (N17)? mem[106] :
                         (N19)? mem[240] :
                         (N21)? mem[374] :
                         (N23)? mem[508] :
                         (N18)? mem[642] :
                         (N20)? mem[776] :
                         (N22)? mem[910] :
                         (N24)? mem[1044] : 1'b0;
  assign r_data_o[105] = (N17)? mem[105] :
                         (N19)? mem[239] :
                         (N21)? mem[373] :
                         (N23)? mem[507] :
                         (N18)? mem[641] :
                         (N20)? mem[775] :
                         (N22)? mem[909] :
                         (N24)? mem[1043] : 1'b0;
  assign r_data_o[104] = (N17)? mem[104] :
                         (N19)? mem[238] :
                         (N21)? mem[372] :
                         (N23)? mem[506] :
                         (N18)? mem[640] :
                         (N20)? mem[774] :
                         (N22)? mem[908] :
                         (N24)? mem[1042] : 1'b0;
  assign r_data_o[103] = (N17)? mem[103] :
                         (N19)? mem[237] :
                         (N21)? mem[371] :
                         (N23)? mem[505] :
                         (N18)? mem[639] :
                         (N20)? mem[773] :
                         (N22)? mem[907] :
                         (N24)? mem[1041] : 1'b0;
  assign r_data_o[102] = (N17)? mem[102] :
                         (N19)? mem[236] :
                         (N21)? mem[370] :
                         (N23)? mem[504] :
                         (N18)? mem[638] :
                         (N20)? mem[772] :
                         (N22)? mem[906] :
                         (N24)? mem[1040] : 1'b0;
  assign r_data_o[101] = (N17)? mem[101] :
                         (N19)? mem[235] :
                         (N21)? mem[369] :
                         (N23)? mem[503] :
                         (N18)? mem[637] :
                         (N20)? mem[771] :
                         (N22)? mem[905] :
                         (N24)? mem[1039] : 1'b0;
  assign r_data_o[100] = (N17)? mem[100] :
                         (N19)? mem[234] :
                         (N21)? mem[368] :
                         (N23)? mem[502] :
                         (N18)? mem[636] :
                         (N20)? mem[770] :
                         (N22)? mem[904] :
                         (N24)? mem[1038] : 1'b0;
  assign r_data_o[99] = (N17)? mem[99] :
                        (N19)? mem[233] :
                        (N21)? mem[367] :
                        (N23)? mem[501] :
                        (N18)? mem[635] :
                        (N20)? mem[769] :
                        (N22)? mem[903] :
                        (N24)? mem[1037] : 1'b0;
  assign r_data_o[98] = (N17)? mem[98] :
                        (N19)? mem[232] :
                        (N21)? mem[366] :
                        (N23)? mem[500] :
                        (N18)? mem[634] :
                        (N20)? mem[768] :
                        (N22)? mem[902] :
                        (N24)? mem[1036] : 1'b0;
  assign r_data_o[97] = (N17)? mem[97] :
                        (N19)? mem[231] :
                        (N21)? mem[365] :
                        (N23)? mem[499] :
                        (N18)? mem[633] :
                        (N20)? mem[767] :
                        (N22)? mem[901] :
                        (N24)? mem[1035] : 1'b0;
  assign r_data_o[96] = (N17)? mem[96] :
                        (N19)? mem[230] :
                        (N21)? mem[364] :
                        (N23)? mem[498] :
                        (N18)? mem[632] :
                        (N20)? mem[766] :
                        (N22)? mem[900] :
                        (N24)? mem[1034] : 1'b0;
  assign r_data_o[95] = (N17)? mem[95] :
                        (N19)? mem[229] :
                        (N21)? mem[363] :
                        (N23)? mem[497] :
                        (N18)? mem[631] :
                        (N20)? mem[765] :
                        (N22)? mem[899] :
                        (N24)? mem[1033] : 1'b0;
  assign r_data_o[94] = (N17)? mem[94] :
                        (N19)? mem[228] :
                        (N21)? mem[362] :
                        (N23)? mem[496] :
                        (N18)? mem[630] :
                        (N20)? mem[764] :
                        (N22)? mem[898] :
                        (N24)? mem[1032] : 1'b0;
  assign r_data_o[93] = (N17)? mem[93] :
                        (N19)? mem[227] :
                        (N21)? mem[361] :
                        (N23)? mem[495] :
                        (N18)? mem[629] :
                        (N20)? mem[763] :
                        (N22)? mem[897] :
                        (N24)? mem[1031] : 1'b0;
  assign r_data_o[92] = (N17)? mem[92] :
                        (N19)? mem[226] :
                        (N21)? mem[360] :
                        (N23)? mem[494] :
                        (N18)? mem[628] :
                        (N20)? mem[762] :
                        (N22)? mem[896] :
                        (N24)? mem[1030] : 1'b0;
  assign r_data_o[91] = (N17)? mem[91] :
                        (N19)? mem[225] :
                        (N21)? mem[359] :
                        (N23)? mem[493] :
                        (N18)? mem[627] :
                        (N20)? mem[761] :
                        (N22)? mem[895] :
                        (N24)? mem[1029] : 1'b0;
  assign r_data_o[90] = (N17)? mem[90] :
                        (N19)? mem[224] :
                        (N21)? mem[358] :
                        (N23)? mem[492] :
                        (N18)? mem[626] :
                        (N20)? mem[760] :
                        (N22)? mem[894] :
                        (N24)? mem[1028] : 1'b0;
  assign r_data_o[89] = (N17)? mem[89] :
                        (N19)? mem[223] :
                        (N21)? mem[357] :
                        (N23)? mem[491] :
                        (N18)? mem[625] :
                        (N20)? mem[759] :
                        (N22)? mem[893] :
                        (N24)? mem[1027] : 1'b0;
  assign r_data_o[88] = (N17)? mem[88] :
                        (N19)? mem[222] :
                        (N21)? mem[356] :
                        (N23)? mem[490] :
                        (N18)? mem[624] :
                        (N20)? mem[758] :
                        (N22)? mem[892] :
                        (N24)? mem[1026] : 1'b0;
  assign r_data_o[87] = (N17)? mem[87] :
                        (N19)? mem[221] :
                        (N21)? mem[355] :
                        (N23)? mem[489] :
                        (N18)? mem[623] :
                        (N20)? mem[757] :
                        (N22)? mem[891] :
                        (N24)? mem[1025] : 1'b0;
  assign r_data_o[86] = (N17)? mem[86] :
                        (N19)? mem[220] :
                        (N21)? mem[354] :
                        (N23)? mem[488] :
                        (N18)? mem[622] :
                        (N20)? mem[756] :
                        (N22)? mem[890] :
                        (N24)? mem[1024] : 1'b0;
  assign r_data_o[85] = (N17)? mem[85] :
                        (N19)? mem[219] :
                        (N21)? mem[353] :
                        (N23)? mem[487] :
                        (N18)? mem[621] :
                        (N20)? mem[755] :
                        (N22)? mem[889] :
                        (N24)? mem[1023] : 1'b0;
  assign r_data_o[84] = (N17)? mem[84] :
                        (N19)? mem[218] :
                        (N21)? mem[352] :
                        (N23)? mem[486] :
                        (N18)? mem[620] :
                        (N20)? mem[754] :
                        (N22)? mem[888] :
                        (N24)? mem[1022] : 1'b0;
  assign r_data_o[83] = (N17)? mem[83] :
                        (N19)? mem[217] :
                        (N21)? mem[351] :
                        (N23)? mem[485] :
                        (N18)? mem[619] :
                        (N20)? mem[753] :
                        (N22)? mem[887] :
                        (N24)? mem[1021] : 1'b0;
  assign r_data_o[82] = (N17)? mem[82] :
                        (N19)? mem[216] :
                        (N21)? mem[350] :
                        (N23)? mem[484] :
                        (N18)? mem[618] :
                        (N20)? mem[752] :
                        (N22)? mem[886] :
                        (N24)? mem[1020] : 1'b0;
  assign r_data_o[81] = (N17)? mem[81] :
                        (N19)? mem[215] :
                        (N21)? mem[349] :
                        (N23)? mem[483] :
                        (N18)? mem[617] :
                        (N20)? mem[751] :
                        (N22)? mem[885] :
                        (N24)? mem[1019] : 1'b0;
  assign r_data_o[80] = (N17)? mem[80] :
                        (N19)? mem[214] :
                        (N21)? mem[348] :
                        (N23)? mem[482] :
                        (N18)? mem[616] :
                        (N20)? mem[750] :
                        (N22)? mem[884] :
                        (N24)? mem[1018] : 1'b0;
  assign r_data_o[79] = (N17)? mem[79] :
                        (N19)? mem[213] :
                        (N21)? mem[347] :
                        (N23)? mem[481] :
                        (N18)? mem[615] :
                        (N20)? mem[749] :
                        (N22)? mem[883] :
                        (N24)? mem[1017] : 1'b0;
  assign r_data_o[78] = (N17)? mem[78] :
                        (N19)? mem[212] :
                        (N21)? mem[346] :
                        (N23)? mem[480] :
                        (N18)? mem[614] :
                        (N20)? mem[748] :
                        (N22)? mem[882] :
                        (N24)? mem[1016] : 1'b0;
  assign r_data_o[77] = (N17)? mem[77] :
                        (N19)? mem[211] :
                        (N21)? mem[345] :
                        (N23)? mem[479] :
                        (N18)? mem[613] :
                        (N20)? mem[747] :
                        (N22)? mem[881] :
                        (N24)? mem[1015] : 1'b0;
  assign r_data_o[76] = (N17)? mem[76] :
                        (N19)? mem[210] :
                        (N21)? mem[344] :
                        (N23)? mem[478] :
                        (N18)? mem[612] :
                        (N20)? mem[746] :
                        (N22)? mem[880] :
                        (N24)? mem[1014] : 1'b0;
  assign r_data_o[75] = (N17)? mem[75] :
                        (N19)? mem[209] :
                        (N21)? mem[343] :
                        (N23)? mem[477] :
                        (N18)? mem[611] :
                        (N20)? mem[745] :
                        (N22)? mem[879] :
                        (N24)? mem[1013] : 1'b0;
  assign r_data_o[74] = (N17)? mem[74] :
                        (N19)? mem[208] :
                        (N21)? mem[342] :
                        (N23)? mem[476] :
                        (N18)? mem[610] :
                        (N20)? mem[744] :
                        (N22)? mem[878] :
                        (N24)? mem[1012] : 1'b0;
  assign r_data_o[73] = (N17)? mem[73] :
                        (N19)? mem[207] :
                        (N21)? mem[341] :
                        (N23)? mem[475] :
                        (N18)? mem[609] :
                        (N20)? mem[743] :
                        (N22)? mem[877] :
                        (N24)? mem[1011] : 1'b0;
  assign r_data_o[72] = (N17)? mem[72] :
                        (N19)? mem[206] :
                        (N21)? mem[340] :
                        (N23)? mem[474] :
                        (N18)? mem[608] :
                        (N20)? mem[742] :
                        (N22)? mem[876] :
                        (N24)? mem[1010] : 1'b0;
  assign r_data_o[71] = (N17)? mem[71] :
                        (N19)? mem[205] :
                        (N21)? mem[339] :
                        (N23)? mem[473] :
                        (N18)? mem[607] :
                        (N20)? mem[741] :
                        (N22)? mem[875] :
                        (N24)? mem[1009] : 1'b0;
  assign r_data_o[70] = (N17)? mem[70] :
                        (N19)? mem[204] :
                        (N21)? mem[338] :
                        (N23)? mem[472] :
                        (N18)? mem[606] :
                        (N20)? mem[740] :
                        (N22)? mem[874] :
                        (N24)? mem[1008] : 1'b0;
  assign r_data_o[69] = (N17)? mem[69] :
                        (N19)? mem[203] :
                        (N21)? mem[337] :
                        (N23)? mem[471] :
                        (N18)? mem[605] :
                        (N20)? mem[739] :
                        (N22)? mem[873] :
                        (N24)? mem[1007] : 1'b0;
  assign r_data_o[68] = (N17)? mem[68] :
                        (N19)? mem[202] :
                        (N21)? mem[336] :
                        (N23)? mem[470] :
                        (N18)? mem[604] :
                        (N20)? mem[738] :
                        (N22)? mem[872] :
                        (N24)? mem[1006] : 1'b0;
  assign r_data_o[67] = (N17)? mem[67] :
                        (N19)? mem[201] :
                        (N21)? mem[335] :
                        (N23)? mem[469] :
                        (N18)? mem[603] :
                        (N20)? mem[737] :
                        (N22)? mem[871] :
                        (N24)? mem[1005] : 1'b0;
  assign r_data_o[66] = (N17)? mem[66] :
                        (N19)? mem[200] :
                        (N21)? mem[334] :
                        (N23)? mem[468] :
                        (N18)? mem[602] :
                        (N20)? mem[736] :
                        (N22)? mem[870] :
                        (N24)? mem[1004] : 1'b0;
  assign r_data_o[65] = (N17)? mem[65] :
                        (N19)? mem[199] :
                        (N21)? mem[333] :
                        (N23)? mem[467] :
                        (N18)? mem[601] :
                        (N20)? mem[735] :
                        (N22)? mem[869] :
                        (N24)? mem[1003] : 1'b0;
  assign r_data_o[64] = (N17)? mem[64] :
                        (N19)? mem[198] :
                        (N21)? mem[332] :
                        (N23)? mem[466] :
                        (N18)? mem[600] :
                        (N20)? mem[734] :
                        (N22)? mem[868] :
                        (N24)? mem[1002] : 1'b0;
  assign r_data_o[63] = (N17)? mem[63] :
                        (N19)? mem[197] :
                        (N21)? mem[331] :
                        (N23)? mem[465] :
                        (N18)? mem[599] :
                        (N20)? mem[733] :
                        (N22)? mem[867] :
                        (N24)? mem[1001] : 1'b0;
  assign r_data_o[62] = (N17)? mem[62] :
                        (N19)? mem[196] :
                        (N21)? mem[330] :
                        (N23)? mem[464] :
                        (N18)? mem[598] :
                        (N20)? mem[732] :
                        (N22)? mem[866] :
                        (N24)? mem[1000] : 1'b0;
  assign r_data_o[61] = (N17)? mem[61] :
                        (N19)? mem[195] :
                        (N21)? mem[329] :
                        (N23)? mem[463] :
                        (N18)? mem[597] :
                        (N20)? mem[731] :
                        (N22)? mem[865] :
                        (N24)? mem[999] : 1'b0;
  assign r_data_o[60] = (N17)? mem[60] :
                        (N19)? mem[194] :
                        (N21)? mem[328] :
                        (N23)? mem[462] :
                        (N18)? mem[596] :
                        (N20)? mem[730] :
                        (N22)? mem[864] :
                        (N24)? mem[998] : 1'b0;
  assign r_data_o[59] = (N17)? mem[59] :
                        (N19)? mem[193] :
                        (N21)? mem[327] :
                        (N23)? mem[461] :
                        (N18)? mem[595] :
                        (N20)? mem[729] :
                        (N22)? mem[863] :
                        (N24)? mem[997] : 1'b0;
  assign r_data_o[58] = (N17)? mem[58] :
                        (N19)? mem[192] :
                        (N21)? mem[326] :
                        (N23)? mem[460] :
                        (N18)? mem[594] :
                        (N20)? mem[728] :
                        (N22)? mem[862] :
                        (N24)? mem[996] : 1'b0;
  assign r_data_o[57] = (N17)? mem[57] :
                        (N19)? mem[191] :
                        (N21)? mem[325] :
                        (N23)? mem[459] :
                        (N18)? mem[593] :
                        (N20)? mem[727] :
                        (N22)? mem[861] :
                        (N24)? mem[995] : 1'b0;
  assign r_data_o[56] = (N17)? mem[56] :
                        (N19)? mem[190] :
                        (N21)? mem[324] :
                        (N23)? mem[458] :
                        (N18)? mem[592] :
                        (N20)? mem[726] :
                        (N22)? mem[860] :
                        (N24)? mem[994] : 1'b0;
  assign r_data_o[55] = (N17)? mem[55] :
                        (N19)? mem[189] :
                        (N21)? mem[323] :
                        (N23)? mem[457] :
                        (N18)? mem[591] :
                        (N20)? mem[725] :
                        (N22)? mem[859] :
                        (N24)? mem[993] : 1'b0;
  assign r_data_o[54] = (N17)? mem[54] :
                        (N19)? mem[188] :
                        (N21)? mem[322] :
                        (N23)? mem[456] :
                        (N18)? mem[590] :
                        (N20)? mem[724] :
                        (N22)? mem[858] :
                        (N24)? mem[992] : 1'b0;
  assign r_data_o[53] = (N17)? mem[53] :
                        (N19)? mem[187] :
                        (N21)? mem[321] :
                        (N23)? mem[455] :
                        (N18)? mem[589] :
                        (N20)? mem[723] :
                        (N22)? mem[857] :
                        (N24)? mem[991] : 1'b0;
  assign r_data_o[52] = (N17)? mem[52] :
                        (N19)? mem[186] :
                        (N21)? mem[320] :
                        (N23)? mem[454] :
                        (N18)? mem[588] :
                        (N20)? mem[722] :
                        (N22)? mem[856] :
                        (N24)? mem[990] : 1'b0;
  assign r_data_o[51] = (N17)? mem[51] :
                        (N19)? mem[185] :
                        (N21)? mem[319] :
                        (N23)? mem[453] :
                        (N18)? mem[587] :
                        (N20)? mem[721] :
                        (N22)? mem[855] :
                        (N24)? mem[989] : 1'b0;
  assign r_data_o[50] = (N17)? mem[50] :
                        (N19)? mem[184] :
                        (N21)? mem[318] :
                        (N23)? mem[452] :
                        (N18)? mem[586] :
                        (N20)? mem[720] :
                        (N22)? mem[854] :
                        (N24)? mem[988] : 1'b0;
  assign r_data_o[49] = (N17)? mem[49] :
                        (N19)? mem[183] :
                        (N21)? mem[317] :
                        (N23)? mem[451] :
                        (N18)? mem[585] :
                        (N20)? mem[719] :
                        (N22)? mem[853] :
                        (N24)? mem[987] : 1'b0;
  assign r_data_o[48] = (N17)? mem[48] :
                        (N19)? mem[182] :
                        (N21)? mem[316] :
                        (N23)? mem[450] :
                        (N18)? mem[584] :
                        (N20)? mem[718] :
                        (N22)? mem[852] :
                        (N24)? mem[986] : 1'b0;
  assign r_data_o[47] = (N17)? mem[47] :
                        (N19)? mem[181] :
                        (N21)? mem[315] :
                        (N23)? mem[449] :
                        (N18)? mem[583] :
                        (N20)? mem[717] :
                        (N22)? mem[851] :
                        (N24)? mem[985] : 1'b0;
  assign r_data_o[46] = (N17)? mem[46] :
                        (N19)? mem[180] :
                        (N21)? mem[314] :
                        (N23)? mem[448] :
                        (N18)? mem[582] :
                        (N20)? mem[716] :
                        (N22)? mem[850] :
                        (N24)? mem[984] : 1'b0;
  assign r_data_o[45] = (N17)? mem[45] :
                        (N19)? mem[179] :
                        (N21)? mem[313] :
                        (N23)? mem[447] :
                        (N18)? mem[581] :
                        (N20)? mem[715] :
                        (N22)? mem[849] :
                        (N24)? mem[983] : 1'b0;
  assign r_data_o[44] = (N17)? mem[44] :
                        (N19)? mem[178] :
                        (N21)? mem[312] :
                        (N23)? mem[446] :
                        (N18)? mem[580] :
                        (N20)? mem[714] :
                        (N22)? mem[848] :
                        (N24)? mem[982] : 1'b0;
  assign r_data_o[43] = (N17)? mem[43] :
                        (N19)? mem[177] :
                        (N21)? mem[311] :
                        (N23)? mem[445] :
                        (N18)? mem[579] :
                        (N20)? mem[713] :
                        (N22)? mem[847] :
                        (N24)? mem[981] : 1'b0;
  assign r_data_o[42] = (N17)? mem[42] :
                        (N19)? mem[176] :
                        (N21)? mem[310] :
                        (N23)? mem[444] :
                        (N18)? mem[578] :
                        (N20)? mem[712] :
                        (N22)? mem[846] :
                        (N24)? mem[980] : 1'b0;
  assign r_data_o[41] = (N17)? mem[41] :
                        (N19)? mem[175] :
                        (N21)? mem[309] :
                        (N23)? mem[443] :
                        (N18)? mem[577] :
                        (N20)? mem[711] :
                        (N22)? mem[845] :
                        (N24)? mem[979] : 1'b0;
  assign r_data_o[40] = (N17)? mem[40] :
                        (N19)? mem[174] :
                        (N21)? mem[308] :
                        (N23)? mem[442] :
                        (N18)? mem[576] :
                        (N20)? mem[710] :
                        (N22)? mem[844] :
                        (N24)? mem[978] : 1'b0;
  assign r_data_o[39] = (N17)? mem[39] :
                        (N19)? mem[173] :
                        (N21)? mem[307] :
                        (N23)? mem[441] :
                        (N18)? mem[575] :
                        (N20)? mem[709] :
                        (N22)? mem[843] :
                        (N24)? mem[977] : 1'b0;
  assign r_data_o[38] = (N17)? mem[38] :
                        (N19)? mem[172] :
                        (N21)? mem[306] :
                        (N23)? mem[440] :
                        (N18)? mem[574] :
                        (N20)? mem[708] :
                        (N22)? mem[842] :
                        (N24)? mem[976] : 1'b0;
  assign r_data_o[37] = (N17)? mem[37] :
                        (N19)? mem[171] :
                        (N21)? mem[305] :
                        (N23)? mem[439] :
                        (N18)? mem[573] :
                        (N20)? mem[707] :
                        (N22)? mem[841] :
                        (N24)? mem[975] : 1'b0;
  assign r_data_o[36] = (N17)? mem[36] :
                        (N19)? mem[170] :
                        (N21)? mem[304] :
                        (N23)? mem[438] :
                        (N18)? mem[572] :
                        (N20)? mem[706] :
                        (N22)? mem[840] :
                        (N24)? mem[974] : 1'b0;
  assign r_data_o[35] = (N17)? mem[35] :
                        (N19)? mem[169] :
                        (N21)? mem[303] :
                        (N23)? mem[437] :
                        (N18)? mem[571] :
                        (N20)? mem[705] :
                        (N22)? mem[839] :
                        (N24)? mem[973] : 1'b0;
  assign r_data_o[34] = (N17)? mem[34] :
                        (N19)? mem[168] :
                        (N21)? mem[302] :
                        (N23)? mem[436] :
                        (N18)? mem[570] :
                        (N20)? mem[704] :
                        (N22)? mem[838] :
                        (N24)? mem[972] : 1'b0;
  assign r_data_o[33] = (N17)? mem[33] :
                        (N19)? mem[167] :
                        (N21)? mem[301] :
                        (N23)? mem[435] :
                        (N18)? mem[569] :
                        (N20)? mem[703] :
                        (N22)? mem[837] :
                        (N24)? mem[971] : 1'b0;
  assign r_data_o[32] = (N17)? mem[32] :
                        (N19)? mem[166] :
                        (N21)? mem[300] :
                        (N23)? mem[434] :
                        (N18)? mem[568] :
                        (N20)? mem[702] :
                        (N22)? mem[836] :
                        (N24)? mem[970] : 1'b0;
  assign r_data_o[31] = (N17)? mem[31] :
                        (N19)? mem[165] :
                        (N21)? mem[299] :
                        (N23)? mem[433] :
                        (N18)? mem[567] :
                        (N20)? mem[701] :
                        (N22)? mem[835] :
                        (N24)? mem[969] : 1'b0;
  assign r_data_o[30] = (N17)? mem[30] :
                        (N19)? mem[164] :
                        (N21)? mem[298] :
                        (N23)? mem[432] :
                        (N18)? mem[566] :
                        (N20)? mem[700] :
                        (N22)? mem[834] :
                        (N24)? mem[968] : 1'b0;
  assign r_data_o[29] = (N17)? mem[29] :
                        (N19)? mem[163] :
                        (N21)? mem[297] :
                        (N23)? mem[431] :
                        (N18)? mem[565] :
                        (N20)? mem[699] :
                        (N22)? mem[833] :
                        (N24)? mem[967] : 1'b0;
  assign r_data_o[28] = (N17)? mem[28] :
                        (N19)? mem[162] :
                        (N21)? mem[296] :
                        (N23)? mem[430] :
                        (N18)? mem[564] :
                        (N20)? mem[698] :
                        (N22)? mem[832] :
                        (N24)? mem[966] : 1'b0;
  assign r_data_o[27] = (N17)? mem[27] :
                        (N19)? mem[161] :
                        (N21)? mem[295] :
                        (N23)? mem[429] :
                        (N18)? mem[563] :
                        (N20)? mem[697] :
                        (N22)? mem[831] :
                        (N24)? mem[965] : 1'b0;
  assign r_data_o[26] = (N17)? mem[26] :
                        (N19)? mem[160] :
                        (N21)? mem[294] :
                        (N23)? mem[428] :
                        (N18)? mem[562] :
                        (N20)? mem[696] :
                        (N22)? mem[830] :
                        (N24)? mem[964] : 1'b0;
  assign r_data_o[25] = (N17)? mem[25] :
                        (N19)? mem[159] :
                        (N21)? mem[293] :
                        (N23)? mem[427] :
                        (N18)? mem[561] :
                        (N20)? mem[695] :
                        (N22)? mem[829] :
                        (N24)? mem[963] : 1'b0;
  assign r_data_o[24] = (N17)? mem[24] :
                        (N19)? mem[158] :
                        (N21)? mem[292] :
                        (N23)? mem[426] :
                        (N18)? mem[560] :
                        (N20)? mem[694] :
                        (N22)? mem[828] :
                        (N24)? mem[962] : 1'b0;
  assign r_data_o[23] = (N17)? mem[23] :
                        (N19)? mem[157] :
                        (N21)? mem[291] :
                        (N23)? mem[425] :
                        (N18)? mem[559] :
                        (N20)? mem[693] :
                        (N22)? mem[827] :
                        (N24)? mem[961] : 1'b0;
  assign r_data_o[22] = (N17)? mem[22] :
                        (N19)? mem[156] :
                        (N21)? mem[290] :
                        (N23)? mem[424] :
                        (N18)? mem[558] :
                        (N20)? mem[692] :
                        (N22)? mem[826] :
                        (N24)? mem[960] : 1'b0;
  assign r_data_o[21] = (N17)? mem[21] :
                        (N19)? mem[155] :
                        (N21)? mem[289] :
                        (N23)? mem[423] :
                        (N18)? mem[557] :
                        (N20)? mem[691] :
                        (N22)? mem[825] :
                        (N24)? mem[959] : 1'b0;
  assign r_data_o[20] = (N17)? mem[20] :
                        (N19)? mem[154] :
                        (N21)? mem[288] :
                        (N23)? mem[422] :
                        (N18)? mem[556] :
                        (N20)? mem[690] :
                        (N22)? mem[824] :
                        (N24)? mem[958] : 1'b0;
  assign r_data_o[19] = (N17)? mem[19] :
                        (N19)? mem[153] :
                        (N21)? mem[287] :
                        (N23)? mem[421] :
                        (N18)? mem[555] :
                        (N20)? mem[689] :
                        (N22)? mem[823] :
                        (N24)? mem[957] : 1'b0;
  assign r_data_o[18] = (N17)? mem[18] :
                        (N19)? mem[152] :
                        (N21)? mem[286] :
                        (N23)? mem[420] :
                        (N18)? mem[554] :
                        (N20)? mem[688] :
                        (N22)? mem[822] :
                        (N24)? mem[956] : 1'b0;
  assign r_data_o[17] = (N17)? mem[17] :
                        (N19)? mem[151] :
                        (N21)? mem[285] :
                        (N23)? mem[419] :
                        (N18)? mem[553] :
                        (N20)? mem[687] :
                        (N22)? mem[821] :
                        (N24)? mem[955] : 1'b0;
  assign r_data_o[16] = (N17)? mem[16] :
                        (N19)? mem[150] :
                        (N21)? mem[284] :
                        (N23)? mem[418] :
                        (N18)? mem[552] :
                        (N20)? mem[686] :
                        (N22)? mem[820] :
                        (N24)? mem[954] : 1'b0;
  assign r_data_o[15] = (N17)? mem[15] :
                        (N19)? mem[149] :
                        (N21)? mem[283] :
                        (N23)? mem[417] :
                        (N18)? mem[551] :
                        (N20)? mem[685] :
                        (N22)? mem[819] :
                        (N24)? mem[953] : 1'b0;
  assign r_data_o[14] = (N17)? mem[14] :
                        (N19)? mem[148] :
                        (N21)? mem[282] :
                        (N23)? mem[416] :
                        (N18)? mem[550] :
                        (N20)? mem[684] :
                        (N22)? mem[818] :
                        (N24)? mem[952] : 1'b0;
  assign r_data_o[13] = (N17)? mem[13] :
                        (N19)? mem[147] :
                        (N21)? mem[281] :
                        (N23)? mem[415] :
                        (N18)? mem[549] :
                        (N20)? mem[683] :
                        (N22)? mem[817] :
                        (N24)? mem[951] : 1'b0;
  assign r_data_o[12] = (N17)? mem[12] :
                        (N19)? mem[146] :
                        (N21)? mem[280] :
                        (N23)? mem[414] :
                        (N18)? mem[548] :
                        (N20)? mem[682] :
                        (N22)? mem[816] :
                        (N24)? mem[950] : 1'b0;
  assign r_data_o[11] = (N17)? mem[11] :
                        (N19)? mem[145] :
                        (N21)? mem[279] :
                        (N23)? mem[413] :
                        (N18)? mem[547] :
                        (N20)? mem[681] :
                        (N22)? mem[815] :
                        (N24)? mem[949] : 1'b0;
  assign r_data_o[10] = (N17)? mem[10] :
                        (N19)? mem[144] :
                        (N21)? mem[278] :
                        (N23)? mem[412] :
                        (N18)? mem[546] :
                        (N20)? mem[680] :
                        (N22)? mem[814] :
                        (N24)? mem[948] : 1'b0;
  assign r_data_o[9] = (N17)? mem[9] :
                       (N19)? mem[143] :
                       (N21)? mem[277] :
                       (N23)? mem[411] :
                       (N18)? mem[545] :
                       (N20)? mem[679] :
                       (N22)? mem[813] :
                       (N24)? mem[947] : 1'b0;
  assign r_data_o[8] = (N17)? mem[8] :
                       (N19)? mem[142] :
                       (N21)? mem[276] :
                       (N23)? mem[410] :
                       (N18)? mem[544] :
                       (N20)? mem[678] :
                       (N22)? mem[812] :
                       (N24)? mem[946] : 1'b0;
  assign r_data_o[7] = (N17)? mem[7] :
                       (N19)? mem[141] :
                       (N21)? mem[275] :
                       (N23)? mem[409] :
                       (N18)? mem[543] :
                       (N20)? mem[677] :
                       (N22)? mem[811] :
                       (N24)? mem[945] : 1'b0;
  assign r_data_o[6] = (N17)? mem[6] :
                       (N19)? mem[140] :
                       (N21)? mem[274] :
                       (N23)? mem[408] :
                       (N18)? mem[542] :
                       (N20)? mem[676] :
                       (N22)? mem[810] :
                       (N24)? mem[944] : 1'b0;
  assign r_data_o[5] = (N17)? mem[5] :
                       (N19)? mem[139] :
                       (N21)? mem[273] :
                       (N23)? mem[407] :
                       (N18)? mem[541] :
                       (N20)? mem[675] :
                       (N22)? mem[809] :
                       (N24)? mem[943] : 1'b0;
  assign r_data_o[4] = (N17)? mem[4] :
                       (N19)? mem[138] :
                       (N21)? mem[272] :
                       (N23)? mem[406] :
                       (N18)? mem[540] :
                       (N20)? mem[674] :
                       (N22)? mem[808] :
                       (N24)? mem[942] : 1'b0;
  assign r_data_o[3] = (N17)? mem[3] :
                       (N19)? mem[137] :
                       (N21)? mem[271] :
                       (N23)? mem[405] :
                       (N18)? mem[539] :
                       (N20)? mem[673] :
                       (N22)? mem[807] :
                       (N24)? mem[941] : 1'b0;
  assign r_data_o[2] = (N17)? mem[2] :
                       (N19)? mem[136] :
                       (N21)? mem[270] :
                       (N23)? mem[404] :
                       (N18)? mem[538] :
                       (N20)? mem[672] :
                       (N22)? mem[806] :
                       (N24)? mem[940] : 1'b0;
  assign r_data_o[1] = (N17)? mem[1] :
                       (N19)? mem[135] :
                       (N21)? mem[269] :
                       (N23)? mem[403] :
                       (N18)? mem[537] :
                       (N20)? mem[671] :
                       (N22)? mem[805] :
                       (N24)? mem[939] : 1'b0;
  assign r_data_o[0] = (N17)? mem[0] :
                       (N19)? mem[134] :
                       (N21)? mem[268] :
                       (N23)? mem[402] :
                       (N18)? mem[536] :
                       (N20)? mem[670] :
                       (N22)? mem[804] :
                       (N24)? mem[938] : 1'b0;
  assign N50 = w_addr_i[0] & w_addr_i[1];
  assign N33 = N50 & w_addr_i[2];
  assign N51 = N0 & w_addr_i[1];
  assign N0 = ~w_addr_i[0];
  assign N32 = N51 & w_addr_i[2];
  assign N52 = w_addr_i[0] & N1;
  assign N1 = ~w_addr_i[1];
  assign N31 = N52 & w_addr_i[2];
  assign N53 = N2 & N3;
  assign N2 = ~w_addr_i[0];
  assign N3 = ~w_addr_i[1];
  assign N30 = N53 & w_addr_i[2];
  assign N29 = N50 & N4;
  assign N4 = ~w_addr_i[2];
  assign N28 = N51 & N5;
  assign N5 = ~w_addr_i[2];
  assign N27 = N52 & N6;
  assign N6 = ~w_addr_i[2];
  assign N26 = N53 & N7;
  assign N7 = ~w_addr_i[2];
  assign { N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34 } = (N8)? { N33, N33, N32, N32, N31, N31, N30, N30, N29, N29, N28, N28, N27, N27, N26, N26 } :
                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N25;
  assign N10 = ~r_addr_i[0];
  assign N11 = ~r_addr_i[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r_addr_i[1];
  assign N14 = r_addr_i[0] & N11;
  assign N15 = r_addr_i[0] & r_addr_i[1];
  assign N16 = ~r_addr_i[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r_addr_i[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r_addr_i[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r_addr_i[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r_addr_i[2];
  assign N25 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N48) begin
      { mem[1071:973], mem[938:938] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N49) begin
      { mem[972:939] } <= { w_data_i[34:1] };
    end
    if(N46) begin
      { mem[937:839], mem[804:804] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N47) begin
      { mem[838:805] } <= { w_data_i[34:1] };
    end
    if(N44) begin
      { mem[803:705], mem[670:670] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N45) begin
      { mem[704:671] } <= { w_data_i[34:1] };
    end
    if(N42) begin
      { mem[669:571], mem[536:536] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N43) begin
      { mem[570:537] } <= { w_data_i[34:1] };
    end
    if(N40) begin
      { mem[535:437], mem[402:402] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N41) begin
      { mem[436:403] } <= { w_data_i[34:1] };
    end
    if(N38) begin
      { mem[401:303], mem[268:268] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N39) begin
      { mem[302:269] } <= { w_data_i[34:1] };
    end
    if(N36) begin
      { mem[267:169], mem[134:134] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N37) begin
      { mem[168:135] } <= { w_data_i[34:1] };
    end
    if(N34) begin
      { mem[133:35], mem[0:0] } <= { w_data_i[133:35], w_data_i[0:0] };
    end
    if(N35) begin
      { mem[34:1] } <= { w_data_i[34:1] };
    end
  end


endmodule



module bsg_mem_1r1w_width_p134_els_p8
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [2:0] w_addr_i;
  input [133:0] w_data_i;
  input [2:0] r_addr_i;
  output [133:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [133:0] r_data_o;

  bsg_mem_p134
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_fifo_1r1w_rolly_width_p134_els_p8_ready_THEN_valid_p1
(
  clk_i,
  reset_i,
  clr_v_i,
  ckpt_v_i,
  roll_v_i,
  data_i,
  v_i,
  ready_o,
  data_o,
  v_o,
  yumi_i
);

  input [133:0] data_i;
  output [133:0] data_o;
  input clk_i;
  input reset_i;
  input clr_v_i;
  input ckpt_v_i;
  input roll_v_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [133:0] data_o;
  wire ready_o,v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,empty,N23,N24,full,N25,N26,N27,N28,N29,N30,N31,N32,N33;
  wire [3:0] cptr_r,rptr_r,rptr_jmp,wptr_r,wptr_jmp;
  assign N21 = rptr_r[2:0] == wptr_r[2:0];
  assign N0 = rptr_r[3] ^ wptr_r[3];
  assign N22 = ~N0;
  assign N23 = cptr_r[2:0] == wptr_r[2:0];
  assign N24 = cptr_r[3] ^ wptr_r[3];

  bsg_circular_ptr_slots_p16_max_add_p1
  cptr_circ_ptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(ckpt_v_i),
    .o(cptr_r)
  );


  bsg_circular_ptr_slots_p16_max_add_p15
  wptr_circ_ptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(wptr_jmp),
    .o(wptr_r)
  );


  bsg_circular_ptr_slots_p16_max_add_p15
  rptr_circ_ptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(rptr_jmp),
    .o(rptr_r)
  );


  bsg_mem_1r1w_width_p134_els_p8
  fifo_mem
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(v_i),
    .w_addr_i(wptr_r[2:0]),
    .w_data_i(data_i),
    .r_v_i(yumi_i),
    .r_addr_i(rptr_r[2:0]),
    .r_data_o(data_o)
  );

  assign { N18, N17, N16, N15 } = rptr_r - wptr_r;
  assign { N9, N8, N7, N6 } = cptr_r - rptr_r;
  assign rptr_jmp = (N1)? { N9, N8, N7, N6 } :
                    (N11)? { 1'b0, 1'b0, 1'b0, 1'b1 } :
                    (N5)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = roll_v_i;
  assign wptr_jmp = (N2)? { N18, N17, N16, N15 } :
                    (N20)? { 1'b0, 1'b0, 1'b0, 1'b1 } :
                    (N14)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2 = clr_v_i;
  assign N3 = yumi_i;
  assign N4 = N3 | roll_v_i;
  assign N5 = ~N4;
  assign N10 = ~roll_v_i;
  assign N11 = N3 & N10;
  assign N12 = v_i;
  assign N13 = N12 | clr_v_i;
  assign N14 = ~N13;
  assign N19 = ~clr_v_i;
  assign N20 = N12 & N19;
  assign empty = N21 & N22;
  assign full = N23 & N24;
  assign ready_o = N27 & N28;
  assign N27 = N25 & N26;
  assign N25 = ~reset_i;
  assign N26 = ~clr_v_i;
  assign N28 = ~full;
  assign v_o = N32 & N33;
  assign N32 = N30 & N31;
  assign N30 = N29 & N26;
  assign N29 = ~reset_i;
  assign N31 = ~roll_v_i;
  assign N33 = ~empty;

endmodule



module bsg_circular_ptr_slots_p2_max_add_p1
(
  clk,
  reset_i,
  add_i,
  o
);

  input [0:0] add_i;
  output [0:0] o;
  input clk;
  input reset_i;
  wire N0,N1,N2,N3,N4,N5,N6;
  wire [0:0] genblk1_genblk1_ptr_r_p1;
  reg [0:0] o;
  assign genblk1_genblk1_ptr_r_p1[0] = o[0] ^ 1'b1;
  assign N3 = (N0)? 1'b0 :
              (N1)? genblk1_genblk1_ptr_r_p1[0] : 1'b0;
  assign N0 = reset_i;
  assign N1 = N2;
  assign N2 = ~reset_i;
  assign N4 = ~add_i[0];
  assign N5 = N4 & N2;
  assign N6 = ~N5;

  always @(posedge clk) begin
    if(N6) begin
      { o[0:0] } <= { N3 };
    end
  end


endmodule



module bsg_fifo_tracker_els_p2
(
  clk_i,
  reset_i,
  enq_i,
  deq_i,
  wptr_r_o,
  rptr_r_o,
  full_o,
  empty_o
);

  output [0:0] wptr_r_o;
  output [0:0] rptr_r_o;
  input clk_i;
  input reset_i;
  input enq_i;
  input deq_i;
  output full_o;
  output empty_o;
  wire [0:0] wptr_r_o,rptr_r_o;
  wire full_o,empty_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,equal_ptrs;
  reg deq_r,enq_r;

  bsg_circular_ptr_slots_p2_max_add_p1
  rptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(deq_i),
    .o(rptr_r_o[0])
  );


  bsg_circular_ptr_slots_p2_max_add_p1
  wptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(enq_i),
    .o(wptr_r_o[0])
  );

  assign N0 = rptr_r_o[0] ^ wptr_r_o[0];
  assign equal_ptrs = ~N0;
  assign N6 = (N1)? 1'b1 :
              (N10)? 1'b1 :
              (N5)? 1'b0 : 1'b0;
  assign N1 = N3;
  assign N7 = (N1)? 1'b0 :
              (N10)? enq_i : 1'b0;
  assign N8 = (N1)? 1'b1 :
              (N10)? deq_i : 1'b0;
  assign N2 = enq_i | deq_i;
  assign N3 = reset_i;
  assign N4 = N2 | N3;
  assign N5 = ~N4;
  assign N9 = ~N3;
  assign N10 = N2 & N9;
  assign empty_o = equal_ptrs & deq_r;
  assign full_o = equal_ptrs & enq_r;

  always @(posedge clk_i) begin
    if(N6) begin
      deq_r <= N8;
      enq_r <= N7;
    end
  end


endmodule



module bsg_mem_p109
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [108:0] w_data_i;
  input [0:0] r_addr_i;
  output [108:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [108:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10;
  reg [217:0] mem;
  assign r_data_o[108] = (N3)? mem[108] :
                         (N0)? mem[217] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[107] = (N3)? mem[107] :
                         (N0)? mem[216] : 1'b0;
  assign r_data_o[106] = (N3)? mem[106] :
                         (N0)? mem[215] : 1'b0;
  assign r_data_o[105] = (N3)? mem[105] :
                         (N0)? mem[214] : 1'b0;
  assign r_data_o[104] = (N3)? mem[104] :
                         (N0)? mem[213] : 1'b0;
  assign r_data_o[103] = (N3)? mem[103] :
                         (N0)? mem[212] : 1'b0;
  assign r_data_o[102] = (N3)? mem[102] :
                         (N0)? mem[211] : 1'b0;
  assign r_data_o[101] = (N3)? mem[101] :
                         (N0)? mem[210] : 1'b0;
  assign r_data_o[100] = (N3)? mem[100] :
                         (N0)? mem[209] : 1'b0;
  assign r_data_o[99] = (N3)? mem[99] :
                        (N0)? mem[208] : 1'b0;
  assign r_data_o[98] = (N3)? mem[98] :
                        (N0)? mem[207] : 1'b0;
  assign r_data_o[97] = (N3)? mem[97] :
                        (N0)? mem[206] : 1'b0;
  assign r_data_o[96] = (N3)? mem[96] :
                        (N0)? mem[205] : 1'b0;
  assign r_data_o[95] = (N3)? mem[95] :
                        (N0)? mem[204] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] :
                        (N0)? mem[203] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] :
                        (N0)? mem[202] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] :
                        (N0)? mem[201] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] :
                        (N0)? mem[200] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] :
                        (N0)? mem[199] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] :
                        (N0)? mem[198] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] :
                        (N0)? mem[197] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] :
                        (N0)? mem[196] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] :
                        (N0)? mem[195] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] :
                        (N0)? mem[194] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] :
                        (N0)? mem[193] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] :
                        (N0)? mem[192] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] :
                        (N0)? mem[191] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] :
                        (N0)? mem[190] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] :
                        (N0)? mem[189] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] :
                        (N0)? mem[188] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] :
                        (N0)? mem[187] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] :
                        (N0)? mem[186] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] :
                        (N0)? mem[185] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] :
                        (N0)? mem[184] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] :
                        (N0)? mem[183] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] :
                        (N0)? mem[182] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] :
                        (N0)? mem[181] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] :
                        (N0)? mem[180] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] :
                        (N0)? mem[179] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] :
                        (N0)? mem[178] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] :
                        (N0)? mem[177] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] :
                        (N0)? mem[176] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] :
                        (N0)? mem[175] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] :
                        (N0)? mem[174] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] :
                        (N0)? mem[173] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] :
                        (N0)? mem[172] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] :
                        (N0)? mem[171] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] :
                        (N0)? mem[170] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] :
                        (N0)? mem[169] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] :
                        (N0)? mem[168] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] :
                        (N0)? mem[167] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] :
                        (N0)? mem[166] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] :
                        (N0)? mem[165] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] :
                        (N0)? mem[164] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] :
                        (N0)? mem[163] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] :
                        (N0)? mem[162] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] :
                        (N0)? mem[161] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] :
                        (N0)? mem[160] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] :
                        (N0)? mem[159] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] :
                        (N0)? mem[158] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] :
                        (N0)? mem[157] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] :
                        (N0)? mem[156] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] :
                        (N0)? mem[155] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] :
                        (N0)? mem[154] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] :
                        (N0)? mem[153] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] :
                        (N0)? mem[152] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] :
                        (N0)? mem[151] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] :
                        (N0)? mem[150] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] :
                        (N0)? mem[149] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] :
                        (N0)? mem[148] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] :
                        (N0)? mem[147] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] :
                        (N0)? mem[146] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] :
                        (N0)? mem[145] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] :
                        (N0)? mem[144] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] :
                        (N0)? mem[143] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] :
                        (N0)? mem[142] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] :
                        (N0)? mem[141] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] :
                        (N0)? mem[140] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] :
                        (N0)? mem[139] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] :
                        (N0)? mem[138] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] :
                        (N0)? mem[137] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] :
                        (N0)? mem[136] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] :
                        (N0)? mem[135] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] :
                        (N0)? mem[134] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] :
                        (N0)? mem[133] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] :
                        (N0)? mem[132] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] :
                        (N0)? mem[131] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] :
                        (N0)? mem[130] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] :
                        (N0)? mem[129] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] :
                        (N0)? mem[128] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] :
                        (N0)? mem[127] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] :
                        (N0)? mem[126] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] :
                        (N0)? mem[125] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] :
                        (N0)? mem[124] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] :
                        (N0)? mem[123] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] :
                        (N0)? mem[122] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] :
                        (N0)? mem[121] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] :
                        (N0)? mem[120] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] :
                        (N0)? mem[119] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] :
                       (N0)? mem[118] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] :
                       (N0)? mem[117] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] :
                       (N0)? mem[116] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] :
                       (N0)? mem[115] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] :
                       (N0)? mem[114] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] :
                       (N0)? mem[113] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] :
                       (N0)? mem[112] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] :
                       (N0)? mem[111] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] :
                       (N0)? mem[110] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] :
                       (N0)? mem[109] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], N5, N5 } :
                               (N2)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N9) begin
      { mem[217:119], mem[109:109] } <= { w_data_i[108:10], w_data_i[0:0] };
    end
    if(N10) begin
      { mem[118:110] } <= { w_data_i[9:1] };
    end
    if(N7) begin
      { mem[108:10], mem[0:0] } <= { w_data_i[108:10], w_data_i[0:0] };
    end
    if(N8) begin
      { mem[9:1] } <= { w_data_i[9:1] };
    end
  end


endmodule



module bsg_mem_1r1w_width_p109_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [108:0] w_data_i;
  input [0:0] r_addr_i;
  output [108:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [108:0] r_data_o;

  bsg_mem_p109
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_fifo_1r1w_small_width_p109_els_p2_ready_THEN_valid_p1
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [108:0] data_i;
  output [108:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [108:0] data_o;
  wire ready_o,v_o,full,empty;
  wire [0:0] wptr_r,rptr_r;

  bsg_fifo_tracker_els_p2
  ft
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .enq_i(v_i),
    .deq_i(yumi_i),
    .wptr_r_o(wptr_r[0]),
    .rptr_r_o(rptr_r[0]),
    .full_o(full),
    .empty_o(empty)
  );


  bsg_mem_1r1w_width_p109_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(v_i),
    .w_addr_i(wptr_r[0]),
    .w_data_i(data_i),
    .r_v_i(v_o),
    .r_addr_i(rptr_r[0]),
    .r_data_o(data_o)
  );

  assign ready_o = ~full;
  assign v_o = ~empty;

endmodule



module bsg_dff_reset_en_64_80000124
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [63:0] data_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69;
  reg [63:0] data_o;
  assign N3 = (N0)? 1'b1 :
              (N69)? 1'b1 :
              (N2)? 1'b0 : 1'b0;
  assign N0 = reset_i;
  assign { N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } :
                                                                                                                                                                                                                                                                                                                                        (N69)? data_i : 1'b0;
  assign N1 = en_i | reset_i;
  assign N2 = ~N1;
  assign N68 = ~reset_i;
  assign N69 = en_i & N68;

  always @(posedge clk_i) begin
    if(N3) begin
      { data_o[63:0] } <= { N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4 };
    end
  end


endmodule



module bsg_mux_width_p64_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [127:0] data_i;
  input [0:0] sel_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1;
  assign data_o[63] = (N1)? data_i[63] :
                      (N0)? data_i[127] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[62] = (N1)? data_i[62] :
                      (N0)? data_i[126] : 1'b0;
  assign data_o[61] = (N1)? data_i[61] :
                      (N0)? data_i[125] : 1'b0;
  assign data_o[60] = (N1)? data_i[60] :
                      (N0)? data_i[124] : 1'b0;
  assign data_o[59] = (N1)? data_i[59] :
                      (N0)? data_i[123] : 1'b0;
  assign data_o[58] = (N1)? data_i[58] :
                      (N0)? data_i[122] : 1'b0;
  assign data_o[57] = (N1)? data_i[57] :
                      (N0)? data_i[121] : 1'b0;
  assign data_o[56] = (N1)? data_i[56] :
                      (N0)? data_i[120] : 1'b0;
  assign data_o[55] = (N1)? data_i[55] :
                      (N0)? data_i[119] : 1'b0;
  assign data_o[54] = (N1)? data_i[54] :
                      (N0)? data_i[118] : 1'b0;
  assign data_o[53] = (N1)? data_i[53] :
                      (N0)? data_i[117] : 1'b0;
  assign data_o[52] = (N1)? data_i[52] :
                      (N0)? data_i[116] : 1'b0;
  assign data_o[51] = (N1)? data_i[51] :
                      (N0)? data_i[115] : 1'b0;
  assign data_o[50] = (N1)? data_i[50] :
                      (N0)? data_i[114] : 1'b0;
  assign data_o[49] = (N1)? data_i[49] :
                      (N0)? data_i[113] : 1'b0;
  assign data_o[48] = (N1)? data_i[48] :
                      (N0)? data_i[112] : 1'b0;
  assign data_o[47] = (N1)? data_i[47] :
                      (N0)? data_i[111] : 1'b0;
  assign data_o[46] = (N1)? data_i[46] :
                      (N0)? data_i[110] : 1'b0;
  assign data_o[45] = (N1)? data_i[45] :
                      (N0)? data_i[109] : 1'b0;
  assign data_o[44] = (N1)? data_i[44] :
                      (N0)? data_i[108] : 1'b0;
  assign data_o[43] = (N1)? data_i[43] :
                      (N0)? data_i[107] : 1'b0;
  assign data_o[42] = (N1)? data_i[42] :
                      (N0)? data_i[106] : 1'b0;
  assign data_o[41] = (N1)? data_i[41] :
                      (N0)? data_i[105] : 1'b0;
  assign data_o[40] = (N1)? data_i[40] :
                      (N0)? data_i[104] : 1'b0;
  assign data_o[39] = (N1)? data_i[39] :
                      (N0)? data_i[103] : 1'b0;
  assign data_o[38] = (N1)? data_i[38] :
                      (N0)? data_i[102] : 1'b0;
  assign data_o[37] = (N1)? data_i[37] :
                      (N0)? data_i[101] : 1'b0;
  assign data_o[36] = (N1)? data_i[36] :
                      (N0)? data_i[100] : 1'b0;
  assign data_o[35] = (N1)? data_i[35] :
                      (N0)? data_i[99] : 1'b0;
  assign data_o[34] = (N1)? data_i[34] :
                      (N0)? data_i[98] : 1'b0;
  assign data_o[33] = (N1)? data_i[33] :
                      (N0)? data_i[97] : 1'b0;
  assign data_o[32] = (N1)? data_i[32] :
                      (N0)? data_i[96] : 1'b0;
  assign data_o[31] = (N1)? data_i[31] :
                      (N0)? data_i[95] : 1'b0;
  assign data_o[30] = (N1)? data_i[30] :
                      (N0)? data_i[94] : 1'b0;
  assign data_o[29] = (N1)? data_i[29] :
                      (N0)? data_i[93] : 1'b0;
  assign data_o[28] = (N1)? data_i[28] :
                      (N0)? data_i[92] : 1'b0;
  assign data_o[27] = (N1)? data_i[27] :
                      (N0)? data_i[91] : 1'b0;
  assign data_o[26] = (N1)? data_i[26] :
                      (N0)? data_i[90] : 1'b0;
  assign data_o[25] = (N1)? data_i[25] :
                      (N0)? data_i[89] : 1'b0;
  assign data_o[24] = (N1)? data_i[24] :
                      (N0)? data_i[88] : 1'b0;
  assign data_o[23] = (N1)? data_i[23] :
                      (N0)? data_i[87] : 1'b0;
  assign data_o[22] = (N1)? data_i[22] :
                      (N0)? data_i[86] : 1'b0;
  assign data_o[21] = (N1)? data_i[21] :
                      (N0)? data_i[85] : 1'b0;
  assign data_o[20] = (N1)? data_i[20] :
                      (N0)? data_i[84] : 1'b0;
  assign data_o[19] = (N1)? data_i[19] :
                      (N0)? data_i[83] : 1'b0;
  assign data_o[18] = (N1)? data_i[18] :
                      (N0)? data_i[82] : 1'b0;
  assign data_o[17] = (N1)? data_i[17] :
                      (N0)? data_i[81] : 1'b0;
  assign data_o[16] = (N1)? data_i[16] :
                      (N0)? data_i[80] : 1'b0;
  assign data_o[15] = (N1)? data_i[15] :
                      (N0)? data_i[79] : 1'b0;
  assign data_o[14] = (N1)? data_i[14] :
                      (N0)? data_i[78] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] :
                      (N0)? data_i[77] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] :
                      (N0)? data_i[76] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] :
                      (N0)? data_i[75] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] :
                      (N0)? data_i[74] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] :
                     (N0)? data_i[73] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] :
                     (N0)? data_i[72] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] :
                     (N0)? data_i[71] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] :
                     (N0)? data_i[70] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] :
                     (N0)? data_i[69] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] :
                     (N0)? data_i[68] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] :
                     (N0)? data_i[67] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] :
                     (N0)? data_i[66] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] :
                     (N0)? data_i[65] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] :
                     (N0)? data_i[64] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_dff_reset_en_width_p1
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire N0,N1,N2,N3,N4,N5,N6;
  reg [0:0] data_o;
  assign N3 = (N0)? 1'b1 :
              (N6)? 1'b1 :
              (N2)? 1'b0 : 1'b0;
  assign N0 = reset_i;
  assign N4 = (N0)? 1'b0 :
              (N6)? data_i[0] : 1'b0;
  assign N1 = en_i | reset_i;
  assign N2 = ~N1;
  assign N5 = ~reset_i;
  assign N6 = en_i & N5;

  always @(posedge clk_i) begin
    if(N3) begin
      { data_o[0:0] } <= { N4 };
    end
  end


endmodule



module bsg_dff_en_width_p64
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [63:0] data_i;
  output [63:0] data_o;
  input clk_i;
  input en_i;
  reg [63:0] data_o;

  always @(posedge clk_i) begin
    if(en_i) begin
      { data_o[63:0] } <= { data_i[63:0] };
    end
  end


endmodule



module bp_be_director_vaddr_width_p39_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36
(
  clk_i,
  reset_i,
  calc_status_i,
  expected_npc_o,
  fe_cmd_o,
  fe_cmd_v_o,
  fe_cmd_ready_i,
  chk_flush_fe_o,
  chk_dequeue_fe_o,
  chk_roll_fe_o,
  mtvec_i,
  mtvec_w_v_i,
  mtvec_o,
  mepc_i,
  mepc_w_v_i,
  mepc_o
);

  input [306:0] calc_status_i;
  output [63:0] expected_npc_o;
  output [108:0] fe_cmd_o;
  input [63:0] mtvec_i;
  output [63:0] mtvec_o;
  input [63:0] mepc_i;
  output [63:0] mepc_o;
  input clk_i;
  input reset_i;
  input fe_cmd_ready_i;
  input mtvec_w_v_i;
  input mepc_w_v_i;
  output fe_cmd_v_o;
  output chk_flush_fe_o;
  output chk_dequeue_fe_o;
  output chk_roll_fe_o;
  wire [63:0] expected_npc_o,mtvec_o,mepc_o,npc_n,ret_mux_o,roll_mux_o,br_mux_o,npc_plus4,
  mepc_mux_lo;
  wire [108:0] fe_cmd_o;
  wire fe_cmd_v_o,chk_flush_fe_o,chk_dequeue_fe_o,chk_roll_fe_o,N0,N1,N2,
  npc_mismatch_v,npc_w_v,n_1_net_,btaken_v,redirect_pending,attaboy_pending,n_10_net_,N3,N4,N5,
  N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26;
  assign fe_cmd_o[107] = 1'b0;
  assign chk_roll_fe_o = calc_status_i[3];

  bsg_dff_reset_en_64_80000124
  npc
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(npc_w_v),
    .data_i(npc_n),
    .data_o(expected_npc_o)
  );


  bsg_mux_width_p64_els_p2
  exception_mux
  (
    .data_i({ ret_mux_o, roll_mux_o }),
    .sel_i(n_1_net_),
    .data_o(npc_n)
  );


  bsg_mux_width_p64_els_p2
  roll_mux
  (
    .data_i({ calc_status_i[67:4], br_mux_o }),
    .sel_i(calc_status_i[3]),
    .data_o(roll_mux_o)
  );


  bsg_mux_width_p64_els_p2
  br_mux
  (
    .data_i({ calc_status_i[290:227], npc_plus4 }),
    .sel_i(btaken_v),
    .data_o(br_mux_o)
  );


  bsg_mux_width_p64_els_p2
  ret_mux
  (
    .data_i({ mepc_o, mtvec_o }),
    .sel_i(calc_status_i[1]),
    .data_o(ret_mux_o)
  );

  assign npc_mismatch_v = expected_npc_o != calc_status_i[187:124];

  bsg_dff_reset_en_width_p1
  redirect_pending_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(calc_status_i[188]),
    .data_i(npc_mismatch_v),
    .data_o(redirect_pending)
  );


  bsg_dff_reset_en_width_p1
  attaboy_pending_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(calc_status_i[188]),
    .data_i(calc_status_i[190]),
    .data_o(attaboy_pending)
  );


  bsg_dff_en_width_p64
  mtvec_csr_reg
  (
    .clk_i(clk_i),
    .data_i(mtvec_i),
    .en_i(mtvec_w_v_i),
    .data_o(mtvec_o)
  );


  bsg_dff_en_width_p64
  mepc_csr_reg
  (
    .clk_i(clk_i),
    .data_i(mepc_mux_lo),
    .en_i(n_10_net_),
    .data_o(mepc_o)
  );


  bsg_mux_width_p64_els_p2
  mepc_mux
  (
    .data_i({ calc_status_i[67:4], mepc_i }),
    .sel_i(calc_status_i[2]),
    .data_o(mepc_mux_lo)
  );

  assign N12 = ~fe_cmd_o[106];
  assign N13 = N12 | fe_cmd_o[108];
  assign N14 = ~N13;
  assign npc_plus4 = expected_npc_o + { 1'b1, 1'b0, 1'b0 };
  assign N8 = ~N7;
  assign { fe_cmd_o[108:108], fe_cmd_o[105:0] } = (N0)? { 1'b0, expected_npc_o, 1'b1, 1'b0, 1'b0, calc_status_i[226:191], N8, 1'b0, 1'b0 } :
                                                  (N1)? { 1'b1, calc_status_i[187:124], calc_status_i[226:191], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                  (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N3;
  assign N1 = N4;
  assign fe_cmd_o[106] = (N0)? 1'b1 :
                         (N11)? 1'b0 :
                         (N2)? 1'b0 : 1'b0;
  assign N2 = 1'b0;
  assign fe_cmd_v_o = (N0)? N9 :
                      (N1)? N10 :
                      (N6)? 1'b0 : 1'b0;
  assign npc_w_v = N18 | calc_status_i[1];
  assign N18 = N17 | calc_status_i[2];
  assign N17 = N16 | calc_status_i[3];
  assign N16 = calc_status_i[188] & N15;
  assign N15 = ~npc_mismatch_v;
  assign n_1_net_ = calc_status_i[2] | calc_status_i[1];
  assign btaken_v = calc_status_i[291] & calc_status_i[189];
  assign n_10_net_ = mepc_w_v_i | calc_status_i[2];
  assign chk_dequeue_fe_o = N19 & calc_status_i[0];
  assign N19 = ~calc_status_i[3];
  assign chk_flush_fe_o = fe_cmd_v_o & N14;
  assign N3 = calc_status_i[188] & npc_mismatch_v;
  assign N4 = N21 & attaboy_pending;
  assign N21 = calc_status_i[188] & N20;
  assign N20 = ~npc_mismatch_v;
  assign N5 = N4 | N3;
  assign N6 = ~N5;
  assign N7 = calc_status_i[190];
  assign N9 = N23 & N24;
  assign N23 = fe_cmd_ready_i & N22;
  assign N22 = ~calc_status_i[3];
  assign N24 = ~redirect_pending;
  assign N10 = N26 & N24;
  assign N26 = fe_cmd_ready_i & N25;
  assign N25 = ~calc_status_i[3];
  assign N11 = ~N3;

endmodule



module bp_be_detector_vaddr_width_p39_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36_load_to_use_forwarding_p1
(
  clk_i,
  reset_i,
  calc_status_i,
  expected_npc_i,
  mmu_cmd_ready_i,
  chk_dispatch_v_o,
  chk_roll_o,
  chk_poison_isd_o,
  chk_poison_ex1_o,
  chk_poison_ex2_o,
  chk_poison_ex3_o
);

  input [306:0] calc_status_i;
  input [63:0] expected_npc_i;
  input clk_i;
  input reset_i;
  input mmu_cmd_ready_i;
  output chk_dispatch_v_o;
  output chk_roll_o;
  output chk_poison_isd_o;
  output chk_poison_ex1_o;
  output chk_poison_ex2_o;
  output chk_poison_ex3_o;
  wire chk_dispatch_v_o,chk_roll_o,chk_poison_isd_o,chk_poison_ex1_o,chk_poison_ex2_o,
  chk_poison_ex3_o,N0,N1,N2,N3,N4,N5,stall_haz_v,data_haz_v,struct_haz_v,N6,
  mispredict_v,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,
  N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,
  N46,N47,N48,N49,N50,N51,N52;
  wire [2:0] rs1_match_vector,rs2_match_vector,frs1_data_haz_v,frs2_data_haz_v;
  wire [1:0] irs1_data_haz_v,irs2_data_haz_v;
  assign chk_roll_o = calc_status_i[3];
  assign N0 = calc_status_i[303:299] == calc_status_i[73:69];
  assign N1 = calc_status_i[296:292] == calc_status_i[73:69];
  assign N2 = calc_status_i[303:299] == calc_status_i[84:80];
  assign N3 = calc_status_i[296:292] == calc_status_i[84:80];
  assign N4 = calc_status_i[303:299] == calc_status_i[95:91];
  assign N5 = calc_status_i[296:292] == calc_status_i[95:91];
  assign N6 = calc_status_i[187:124] != expected_npc_i;
  assign N7 = calc_status_i[302] | calc_status_i[303];
  assign N8 = calc_status_i[301] | N7;
  assign N9 = calc_status_i[300] | N8;
  assign N10 = calc_status_i[299] | N9;
  assign N11 = calc_status_i[295] | calc_status_i[296];
  assign N12 = calc_status_i[294] | N11;
  assign N13 = calc_status_i[293] | N12;
  assign N14 = calc_status_i[292] | N13;
  assign rs1_match_vector[0] = N10 & N0;
  assign rs2_match_vector[0] = N14 & N1;
  assign rs1_match_vector[1] = N10 & N2;
  assign rs2_match_vector[1] = N14 & N3;
  assign rs1_match_vector[2] = N10 & N4;
  assign rs2_match_vector[2] = N14 & N5;
  assign irs1_data_haz_v[0] = N15 & N16;
  assign N15 = calc_status_i[305] & rs1_match_vector[0];
  assign N16 = calc_status_i[78] | calc_status_i[77];
  assign irs2_data_haz_v[0] = N17 & N18;
  assign N17 = calc_status_i[298] & rs2_match_vector[0];
  assign N18 = calc_status_i[78] | calc_status_i[77];
  assign frs1_data_haz_v[0] = N19 & N20;
  assign N19 = calc_status_i[304] & rs1_match_vector[0];
  assign N20 = calc_status_i[76] | calc_status_i[75];
  assign frs2_data_haz_v[0] = N21 & N22;
  assign N21 = calc_status_i[297] & rs2_match_vector[0];
  assign N22 = calc_status_i[76] | calc_status_i[75];
  assign irs1_data_haz_v[1] = N23 & calc_status_i[88];
  assign N23 = calc_status_i[305] & rs1_match_vector[1];
  assign irs2_data_haz_v[1] = N24 & calc_status_i[88];
  assign N24 = calc_status_i[298] & rs2_match_vector[1];
  assign frs1_data_haz_v[1] = N25 & N26;
  assign N25 = calc_status_i[304] & rs1_match_vector[1];
  assign N26 = calc_status_i[87] | calc_status_i[86];
  assign frs2_data_haz_v[1] = N27 & N28;
  assign N27 = calc_status_i[297] & rs2_match_vector[1];
  assign N28 = calc_status_i[87] | calc_status_i[86];
  assign frs1_data_haz_v[2] = N29 & calc_status_i[97];
  assign N29 = calc_status_i[304] & rs1_match_vector[2];
  assign frs2_data_haz_v[2] = N30 & calc_status_i[97];
  assign N30 = calc_status_i[297] & rs2_match_vector[2];
  assign stall_haz_v = N32 | calc_status_i[107];
  assign N32 = N31 | calc_status_i[96];
  assign N31 = calc_status_i[74] | calc_status_i[85];
  assign data_haz_v = N39 | N41;
  assign N39 = N36 | N38;
  assign N36 = N34 | N35;
  assign N34 = stall_haz_v | N33;
  assign N33 = irs1_data_haz_v[1] | irs1_data_haz_v[0];
  assign N35 = irs2_data_haz_v[1] | irs2_data_haz_v[0];
  assign N38 = N37 | frs1_data_haz_v[0];
  assign N37 = frs1_data_haz_v[2] | frs1_data_haz_v[1];
  assign N41 = N40 | frs2_data_haz_v[0];
  assign N40 = frs2_data_haz_v[2] | frs2_data_haz_v[1];
  assign struct_haz_v = ~mmu_cmd_ready_i;
  assign mispredict_v = calc_status_i[188] & N6;
  assign chk_dispatch_v_o = N43 | calc_status_i[3];
  assign N43 = ~N42;
  assign N42 = data_haz_v | struct_haz_v;
  assign chk_poison_isd_o = N45 | calc_status_i[1];
  assign N45 = N44 | calc_status_i[2];
  assign N44 = reset_i | calc_status_i[3];
  assign chk_poison_ex1_o = N48 | calc_status_i[1];
  assign N48 = N47 | calc_status_i[2];
  assign N47 = N46 | calc_status_i[3];
  assign N46 = reset_i | mispredict_v;
  assign chk_poison_ex2_o = N50 | calc_status_i[1];
  assign N50 = N49 | calc_status_i[2];
  assign N49 = reset_i | calc_status_i[3];
  assign chk_poison_ex3_o = N52 | calc_status_i[1];
  assign N52 = N51 | calc_status_i[2];
  assign N51 = reset_i | calc_status_i[3];

endmodule



module bsg_dff_reset_en_width_p8
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [7:0] data_i;
  output [7:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13;
  reg [7:0] data_o;
  assign N3 = (N0)? 1'b1 :
              (N13)? 1'b1 :
              (N2)? 1'b0 : 1'b0;
  assign N0 = reset_i;
  assign { N11, N10, N9, N8, N7, N6, N5, N4 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                (N13)? data_i : 1'b0;
  assign N1 = en_i | reset_i;
  assign N2 = ~N1;
  assign N12 = ~reset_i;
  assign N13 = en_i & N12;

  always @(posedge clk_i) begin
    if(N3) begin
      { data_o[7:0] } <= { N11, N10, N9, N8, N7, N6, N5, N4 };
    end
  end


endmodule



module bp_be_scheduler_vaddr_width_p39_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36
(
  clk_i,
  reset_i,
  fe_queue_i,
  fe_queue_v_i,
  fe_queue_ready_o,
  issue_pkt_o,
  issue_pkt_v_o,
  issue_pkt_ready_i
);

  input [133:0] fe_queue_i;
  output [220:0] issue_pkt_o;
  input clk_i;
  input reset_i;
  input fe_queue_v_i;
  input issue_pkt_ready_i;
  output fe_queue_ready_o;
  output issue_pkt_v_o;
  wire [220:0] issue_pkt_o;
  wire fe_queue_ready_o,issue_pkt_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,
  n_0_net_,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,
  N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,
  N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,
  N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,
  N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,
  N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,
  N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,
  N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,
  N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,
  N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,
  N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,
  N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,
  N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,
  N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,
  N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
  N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,
  N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,
  N302,N303,N304,N305,N306,N307,N308;
  wire [7:0] itag_r,itag_n;
  assign issue_pkt_o[74] = 1'b0;
  assign issue_pkt_o[75] = 1'b0;
  assign issue_pkt_o[212] = fe_queue_i[132];
  assign issue_pkt_o[145] = fe_queue_i[36];
  assign issue_pkt_o[144] = fe_queue_i[35];
  assign issue_pkt_o[143] = fe_queue_i[34];
  assign issue_pkt_o[142] = fe_queue_i[33];
  assign issue_pkt_o[141] = fe_queue_i[32];
  assign issue_pkt_o[140] = fe_queue_i[31];
  assign issue_pkt_o[139] = fe_queue_i[30];
  assign issue_pkt_o[138] = fe_queue_i[29];
  assign issue_pkt_o[137] = fe_queue_i[28];
  assign issue_pkt_o[136] = fe_queue_i[27];
  assign issue_pkt_o[135] = fe_queue_i[26];
  assign issue_pkt_o[134] = fe_queue_i[25];
  assign issue_pkt_o[133] = fe_queue_i[24];
  assign issue_pkt_o[132] = fe_queue_i[23];
  assign issue_pkt_o[131] = fe_queue_i[22];
  assign issue_pkt_o[130] = fe_queue_i[21];
  assign issue_pkt_o[129] = fe_queue_i[20];
  assign issue_pkt_o[128] = fe_queue_i[19];
  assign issue_pkt_o[127] = fe_queue_i[18];
  assign issue_pkt_o[126] = fe_queue_i[17];
  assign issue_pkt_o[125] = fe_queue_i[16];
  assign issue_pkt_o[124] = fe_queue_i[15];
  assign issue_pkt_o[123] = fe_queue_i[14];
  assign issue_pkt_o[122] = fe_queue_i[13];
  assign issue_pkt_o[121] = fe_queue_i[12];
  assign issue_pkt_o[120] = fe_queue_i[11];
  assign issue_pkt_o[119] = fe_queue_i[10];
  assign issue_pkt_o[118] = fe_queue_i[9];
  assign issue_pkt_o[117] = fe_queue_i[8];
  assign issue_pkt_o[116] = fe_queue_i[7];
  assign issue_pkt_o[115] = fe_queue_i[6];
  assign issue_pkt_o[114] = fe_queue_i[5];
  assign issue_pkt_o[113] = fe_queue_i[4];
  assign issue_pkt_o[112] = fe_queue_i[3];
  assign issue_pkt_o[111] = fe_queue_i[2];
  assign issue_pkt_o[110] = fe_queue_i[1];
  assign issue_pkt_o[109] = fe_queue_i[68];
  assign issue_pkt_o[108] = fe_queue_i[67];
  assign issue_pkt_o[107] = fe_queue_i[66];
  assign issue_pkt_o[106] = fe_queue_i[65];
  assign issue_pkt_o[105] = fe_queue_i[64];
  assign issue_pkt_o[104] = fe_queue_i[63];
  assign issue_pkt_o[103] = fe_queue_i[62];
  assign issue_pkt_o[102] = fe_queue_i[61];
  assign issue_pkt_o[101] = fe_queue_i[60];
  assign issue_pkt_o[100] = fe_queue_i[59];
  assign issue_pkt_o[99] = fe_queue_i[58];
  assign issue_pkt_o[98] = fe_queue_i[57];
  assign issue_pkt_o[97] = fe_queue_i[56];
  assign issue_pkt_o[96] = fe_queue_i[55];
  assign issue_pkt_o[95] = fe_queue_i[54];
  assign issue_pkt_o[94] = fe_queue_i[53];
  assign issue_pkt_o[93] = fe_queue_i[52];
  assign issue_pkt_o[92] = fe_queue_i[51];
  assign issue_pkt_o[91] = fe_queue_i[50];
  assign issue_pkt_o[90] = fe_queue_i[49];
  assign issue_pkt_o[89] = fe_queue_i[48];
  assign issue_pkt_o[88] = fe_queue_i[47];
  assign issue_pkt_o[87] = fe_queue_i[46];
  assign issue_pkt_o[86] = fe_queue_i[45];
  assign issue_pkt_o[85] = fe_queue_i[44];
  assign issue_pkt_o[84] = fe_queue_i[43];
  assign issue_pkt_o[83] = fe_queue_i[42];
  assign issue_pkt_o[82] = fe_queue_i[41];
  assign issue_pkt_o[81] = fe_queue_i[40];
  assign issue_pkt_o[80] = fe_queue_i[39];
  assign issue_pkt_o[79] = fe_queue_i[38];
  assign issue_pkt_o[78] = fe_queue_i[37];

  bsg_dff_reset_en_width_p8
  itag_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(n_0_net_),
    .data_i(itag_n),
    .data_o(itag_r)
  );

  assign N15 = fe_queue_i[38] & fe_queue_i[37];
  assign N20 = fe_queue_i[43] | N17;
  assign N21 = N18 | fe_queue_i[40];
  assign N22 = N20 | N21;
  assign N23 = N22 | N19;
  assign N24 = fe_queue_i[43] | fe_queue_i[42];
  assign N25 = N18 | fe_queue_i[40];
  assign N26 = N24 | N25;
  assign N27 = N26 | N19;
  assign N30 = N28 | N17;
  assign N31 = fe_queue_i[41] | N29;
  assign N32 = N30 | N31;
  assign N33 = N32 | N19;
  assign N35 = N28 | N17;
  assign N36 = fe_queue_i[41] | fe_queue_i[40];
  assign N37 = N35 | N36;
  assign N38 = N37 | N19;
  assign N39 = N28 & N17;
  assign N40 = N18 & N29;
  assign N41 = N39 & N40;
  assign N42 = N41 & N19;
  assign N43 = fe_queue_i[43] | fe_queue_i[42];
  assign N44 = N18 | fe_queue_i[40];
  assign N45 = N43 | N44;
  assign N46 = N45 | fe_queue_i[39];
  assign N47 = fe_queue_i[43] | fe_queue_i[42];
  assign N48 = N18 | N29;
  assign N49 = N47 | N48;
  assign N50 = N49 | fe_queue_i[39];
  assign N51 = N28 | N17;
  assign N52 = N18 | fe_queue_i[40];
  assign N53 = N51 | N52;
  assign N54 = N53 | fe_queue_i[39];
  assign N56 = N28 | N17;
  assign N57 = fe_queue_i[41] | fe_queue_i[40];
  assign N58 = N56 | N57;
  assign N59 = N58 | fe_queue_i[39];
  assign N60 = fe_queue_i[43] | N17;
  assign N61 = fe_queue_i[41] | fe_queue_i[40];
  assign N62 = N60 | N61;
  assign N63 = N62 | fe_queue_i[39];
  assign N64 = fe_queue_i[43] | N17;
  assign N65 = N18 | fe_queue_i[40];
  assign N66 = N64 | N65;
  assign N67 = N66 | fe_queue_i[39];
  assign N68 = fe_queue_i[43] | N17;
  assign N69 = N18 | N29;
  assign N70 = N68 | N69;
  assign N71 = N70 | fe_queue_i[39];
  assign N73 = fe_queue_i[43] & fe_queue_i[41];
  assign N74 = N73 & fe_queue_i[39];
  assign N75 = fe_queue_i[43] & fe_queue_i[41];
  assign N76 = N75 & fe_queue_i[40];
  assign N77 = fe_queue_i[41] & fe_queue_i[40];
  assign N78 = N77 & fe_queue_i[39];
  assign N79 = N28 & N18;
  assign N80 = N79 & fe_queue_i[39];
  assign N81 = N17 & N18;
  assign N82 = N81 & fe_queue_i[39];
  assign N83 = N18 & fe_queue_i[40];
  assign N84 = N83 & N19;
  assign N85 = fe_queue_i[43] & N17;
  assign N90 = fe_queue_i[38] & fe_queue_i[37];
  assign N92 = fe_queue_i[43] | N17;
  assign N93 = N18 | fe_queue_i[40];
  assign N94 = N92 | N93;
  assign N95 = N94 | N19;
  assign N96 = fe_queue_i[43] | fe_queue_i[42];
  assign N97 = N18 | fe_queue_i[40];
  assign N98 = N96 | N97;
  assign N99 = N98 | N19;
  assign N101 = N28 | N17;
  assign N102 = fe_queue_i[41] | N29;
  assign N103 = N101 | N102;
  assign N104 = N103 | N19;
  assign N106 = N28 | N17;
  assign N107 = fe_queue_i[41] | fe_queue_i[40];
  assign N108 = N106 | N107;
  assign N109 = N108 | fe_queue_i[39];
  assign N111 = fe_queue_i[43] | N17;
  assign N112 = fe_queue_i[41] | fe_queue_i[40];
  assign N113 = N111 | N112;
  assign N114 = N113 | fe_queue_i[39];
  assign N116 = N28 | N17;
  assign N117 = fe_queue_i[41] | fe_queue_i[40];
  assign N118 = N116 | N117;
  assign N119 = N118 | N19;
  assign N120 = N28 & N17;
  assign N121 = N18 & N29;
  assign N122 = N120 & N121;
  assign N123 = N122 & N19;
  assign N124 = fe_queue_i[43] | fe_queue_i[42];
  assign N125 = N18 | fe_queue_i[40];
  assign N126 = N124 | N125;
  assign N127 = N126 | fe_queue_i[39];
  assign N128 = fe_queue_i[43] | fe_queue_i[42];
  assign N129 = N18 | N29;
  assign N130 = N128 | N129;
  assign N131 = N130 | fe_queue_i[39];
  assign N133 = fe_queue_i[41] & fe_queue_i[40];
  assign N134 = N133 & fe_queue_i[39];
  assign N135 = N28 & N18;
  assign N136 = N135 & fe_queue_i[39];
  assign N137 = N17 & N18;
  assign N138 = N137 & fe_queue_i[39];
  assign N139 = fe_queue_i[43] & fe_queue_i[41];
  assign N140 = fe_queue_i[42] & fe_queue_i[41];
  assign N141 = N140 & N19;
  assign N142 = N18 & fe_queue_i[40];
  assign N143 = N142 & N19;
  assign N144 = fe_queue_i[43] & N17;
  assign N145 = N144 & N19;
  assign itag_n = itag_r + 1'b1;
  assign N87 = (N0)? 1'b0 :
               (N1)? 1'b1 :
               (N2)? 1'b1 :
               (N3)? 1'b0 : 1'b0;
  assign N0 = N34;
  assign N1 = N55;
  assign N2 = N72;
  assign N3 = N86;
  assign { N89, N88 } = (N4)? { N87, N72 } :
                        (N16)? { 1'b0, 1'b0 } : 1'b0;
  assign N4 = N15;
  assign { N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147 } = (N5)? { fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:49], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                                                                                                                                                                                                                                                                              (N6)? { fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[56:49], fe_queue_i[57:57], fe_queue_i[67:58], 1'b0 } :
                                                                                                                                                                                                                                                                                                                                                                                                              (N7)? { fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[44:44], fe_queue_i[67:62], fe_queue_i[48:45], 1'b0 } :
                                                                                                                                                                                                                                                                                                                                                                                                              (N8)? { fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:62], fe_queue_i[48:44] } :
                                                                                                                                                                                                                                                                                                                                                                                                              (N9)? { fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:68], fe_queue_i[68:57] } :
                                                                                                                                                                                                                                                                                                                                                                                                              (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N5 = N100;
  assign N6 = N105;
  assign N7 = N110;
  assign N8 = N115;
  assign N9 = N132;
  assign N10 = N146;
  assign { N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211 } = (N11)? { N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147 } :
                                                                                                                                                                                                                                                                                                                                                                                                              (N91)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = N90;
  assign { issue_pkt_o[220:213], issue_pkt_o[211:149], issue_pkt_o[147:146] } = (N12)? { itag_r, fe_queue_i[131:69], 1'b0, 1'b0 } :
                                                                                (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:132], fe_queue_i[132:92] } : 1'b0;
  assign N12 = N14;
  assign N13 = issue_pkt_o[148];
  assign { issue_pkt_o[77:76], issue_pkt_o[73:0] } = (N12)? { N89, N88, fe_queue_i[56:52], fe_queue_i[61:57], N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211 } :
                                                     (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign fe_queue_ready_o = fe_queue_v_i & issue_pkt_ready_i;
  assign issue_pkt_v_o = fe_queue_v_i & issue_pkt_ready_i;
  assign n_0_net_ = issue_pkt_ready_i & issue_pkt_v_o;
  assign N14 = ~fe_queue_i[133];
  assign issue_pkt_o[148] = fe_queue_i[133];
  assign N16 = ~N15;
  assign N17 = ~fe_queue_i[42];
  assign N18 = ~fe_queue_i[41];
  assign N19 = ~fe_queue_i[39];
  assign N28 = ~fe_queue_i[43];
  assign N29 = ~fe_queue_i[40];
  assign N34 = N277 | N278;
  assign N277 = N275 | N276;
  assign N275 = ~N23;
  assign N276 = ~N27;
  assign N278 = ~N33;
  assign N55 = N284 | N285;
  assign N284 = N282 | N283;
  assign N282 = N280 | N281;
  assign N280 = N279 | N42;
  assign N279 = ~N38;
  assign N281 = ~N46;
  assign N283 = ~N50;
  assign N285 = ~N54;
  assign N72 = N290 | N291;
  assign N290 = N288 | N289;
  assign N288 = N286 | N287;
  assign N286 = ~N59;
  assign N287 = ~N63;
  assign N289 = ~N67;
  assign N291 = ~N71;
  assign N86 = N74 | N296;
  assign N296 = N76 | N295;
  assign N295 = N78 | N294;
  assign N294 = N80 | N293;
  assign N293 = N82 | N292;
  assign N292 = N84 | N85;
  assign N91 = ~N90;
  assign N100 = N297 | N298;
  assign N297 = ~N95;
  assign N298 = ~N99;
  assign N105 = ~N104;
  assign N110 = ~N109;
  assign N115 = ~N114;
  assign N132 = N302 | N303;
  assign N302 = N300 | N301;
  assign N300 = N299 | N123;
  assign N299 = ~N119;
  assign N301 = ~N127;
  assign N303 = ~N131;
  assign N146 = N134 | N308;
  assign N308 = N136 | N307;
  assign N307 = N138 | N306;
  assign N306 = N139 | N305;
  assign N305 = N141 | N304;
  assign N304 = N143 | N145;

endmodule



module bp_be_checker_top_vaddr_width_p39_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36_load_to_use_forwarding_p1
(
  clk_i,
  reset_i,
  fe_cmd_o,
  fe_cmd_v_o,
  fe_cmd_ready_i,
  fe_queue_i,
  fe_queue_v_i,
  fe_queue_ready_o,
  chk_roll_fe_o,
  chk_flush_fe_o,
  chk_dequeue_fe_o,
  issue_pkt_o,
  issue_pkt_v_o,
  issue_pkt_ready_i,
  calc_status_i,
  mmu_cmd_ready_i,
  chk_dispatch_v_o,
  chk_roll_o,
  chk_poison_isd_o,
  chk_poison_ex1_o,
  chk_poison_ex2_o,
  chk_poison_ex3_o,
  mtvec_i,
  mtvec_w_v_i,
  mtvec_o,
  mepc_i,
  mepc_w_v_i,
  mepc_o
);

  output [108:0] fe_cmd_o;
  input [133:0] fe_queue_i;
  output [220:0] issue_pkt_o;
  input [306:0] calc_status_i;
  input [63:0] mtvec_i;
  output [63:0] mtvec_o;
  input [63:0] mepc_i;
  output [63:0] mepc_o;
  input clk_i;
  input reset_i;
  input fe_cmd_ready_i;
  input fe_queue_v_i;
  input issue_pkt_ready_i;
  input mmu_cmd_ready_i;
  input mtvec_w_v_i;
  input mepc_w_v_i;
  output fe_cmd_v_o;
  output fe_queue_ready_o;
  output chk_roll_fe_o;
  output chk_flush_fe_o;
  output chk_dequeue_fe_o;
  output issue_pkt_v_o;
  output chk_dispatch_v_o;
  output chk_roll_o;
  output chk_poison_isd_o;
  output chk_poison_ex1_o;
  output chk_poison_ex2_o;
  output chk_poison_ex3_o;
  wire [108:0] fe_cmd_o;
  wire [220:0] issue_pkt_o;
  wire [63:0] mtvec_o,mepc_o,expected_npc;
  wire fe_cmd_v_o,fe_queue_ready_o,chk_roll_fe_o,chk_flush_fe_o,chk_dequeue_fe_o,
  issue_pkt_v_o,chk_dispatch_v_o,chk_roll_o,chk_poison_isd_o,chk_poison_ex1_o,
  chk_poison_ex2_o,chk_poison_ex3_o;

  bp_be_director_vaddr_width_p39_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36
  director
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .calc_status_i(calc_status_i),
    .expected_npc_o(expected_npc),
    .fe_cmd_o(fe_cmd_o),
    .fe_cmd_v_o(fe_cmd_v_o),
    .fe_cmd_ready_i(fe_cmd_ready_i),
    .chk_flush_fe_o(chk_flush_fe_o),
    .chk_dequeue_fe_o(chk_dequeue_fe_o),
    .chk_roll_fe_o(chk_roll_fe_o),
    .mtvec_i(mtvec_i),
    .mtvec_w_v_i(mtvec_w_v_i),
    .mtvec_o(mtvec_o),
    .mepc_i(mepc_i),
    .mepc_w_v_i(mepc_w_v_i),
    .mepc_o(mepc_o)
  );


  bp_be_detector_vaddr_width_p39_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36_load_to_use_forwarding_p1
  detector
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .calc_status_i(calc_status_i),
    .expected_npc_i(expected_npc),
    .mmu_cmd_ready_i(mmu_cmd_ready_i),
    .chk_dispatch_v_o(chk_dispatch_v_o),
    .chk_roll_o(chk_roll_o),
    .chk_poison_isd_o(chk_poison_isd_o),
    .chk_poison_ex1_o(chk_poison_ex1_o),
    .chk_poison_ex2_o(chk_poison_ex2_o),
    .chk_poison_ex3_o(chk_poison_ex3_o)
  );


  bp_be_scheduler_vaddr_width_p39_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36
  scheduler
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .fe_queue_i(fe_queue_i),
    .fe_queue_v_i(fe_queue_v_i),
    .fe_queue_ready_o(fe_queue_ready_o),
    .issue_pkt_o(issue_pkt_o),
    .issue_pkt_v_o(issue_pkt_v_o),
    .issue_pkt_ready_i(issue_pkt_ready_i)
  );


endmodule



module bsg_mem_2r1w_sync_width_p64_els_p32_read_write_same_addr_p1_harden_p1
(
  clk_i,
  reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r0_v_i,
  r0_addr_i,
  r0_data_o,
  r1_v_i,
  r1_addr_i,
  r1_data_o
);

  input [4:0] w_addr_i;
  input [63:0] w_data_i;
  input [4:0] r0_addr_i;
  output [63:0] r0_data_o;
  input [4:0] r1_addr_i;
  output [63:0] r1_data_o;
  input clk_i;
  input reset_i;
  input w_v_i;
  input r0_v_i;
  input r1_v_i;
  wire [63:0] r0_data_o,r1_data_o;

  hard_mem_1r1w_d32_w64_wrapper
  macro_mem0
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r0_v_i),
    .r_addr_i(r0_addr_i),
    .r_data_o(r0_data_o)
  );


  hard_mem_1r1w_d32_w64_wrapper
  macro_mem1
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r1_v_i),
    .r_addr_i(r1_addr_i),
    .r_data_o(r1_data_o)
  );


endmodule



module bsg_dff_en_width_p5
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [4:0] data_i;
  output [4:0] data_o;
  input clk_i;
  input en_i;
  reg [4:0] data_o;

  always @(posedge clk_i) begin
    if(en_i) begin
      { data_o[4:0] } <= { data_i[4:0] };
    end
  end


endmodule



module bp_be_regfile
(
  clk_i,
  reset_i,
  issue_v_i,
  dispatch_v_i,
  rd_w_v_i,
  rd_addr_i,
  rd_data_i,
  rs1_r_v_i,
  rs1_addr_i,
  rs1_data_o,
  rs2_r_v_i,
  rs2_addr_i,
  rs2_data_o
);

  input [4:0] rd_addr_i;
  input [63:0] rd_data_i;
  input [4:0] rs1_addr_i;
  output [63:0] rs1_data_o;
  input [4:0] rs2_addr_i;
  output [63:0] rs2_data_o;
  input clk_i;
  input reset_i;
  input issue_v_i;
  input dispatch_v_i;
  input rd_w_v_i;
  input rs1_r_v_i;
  input rs2_r_v_i;
  wire [63:0] rs1_data_o,rs2_data_o,rs1_reg_data,rs2_reg_data;
  wire N0,N1,N2,N3,N4,N5,N6,N7,rs1_read_v,rs2_read_v,rs1_issue_v,rs2_issue_v,N8,N9,N10,
  N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;
  wire [4:0] rs1_reread_addr,rs2_reread_addr,rs1_addr_r,rs2_addr_r;

  bsg_mem_2r1w_sync_width_p64_els_p32_read_write_same_addr_p1_harden_p1
  rf
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(rd_w_v_i),
    .w_addr_i(rd_addr_i),
    .w_data_i(rd_data_i),
    .r0_v_i(rs1_read_v),
    .r0_addr_i(rs1_reread_addr),
    .r0_data_o(rs1_reg_data),
    .r1_v_i(rs2_read_v),
    .r1_addr_i(rs2_reread_addr),
    .r1_data_o(rs2_reg_data)
  );


  bsg_dff_en_width_p5
  rs1_addr
  (
    .clk_i(clk_i),
    .data_i(rs1_addr_i),
    .en_i(rs1_issue_v),
    .data_o(rs1_addr_r)
  );


  bsg_dff_en_width_p5
  rs2_addr
  (
    .clk_i(clk_i),
    .data_i(rs2_addr_i),
    .en_i(rs2_issue_v),
    .data_o(rs2_addr_r)
  );

  assign N12 = rs1_addr_r[3] | rs1_addr_r[4];
  assign N13 = rs1_addr_r[2] | N12;
  assign N14 = rs1_addr_r[1] | N13;
  assign N15 = rs1_addr_r[0] | N14;
  assign N16 = ~N15;
  assign N17 = rs2_addr_r[3] | rs2_addr_r[4];
  assign N18 = rs2_addr_r[2] | N17;
  assign N19 = rs2_addr_r[1] | N18;
  assign N20 = rs2_addr_r[0] | N19;
  assign N21 = ~N20;
  assign rs1_reread_addr = (N0)? rs1_addr_i :
                           (N1)? rs1_addr_r : 1'b0;
  assign N0 = N9;
  assign N1 = N8;
  assign rs2_reread_addr = (N2)? rs2_addr_i :
                           (N3)? rs2_addr_r : 1'b0;
  assign N2 = N11;
  assign N3 = N10;
  assign rs1_data_o = (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                      (N5)? rs1_reg_data : 1'b0;
  assign N4 = N16;
  assign N5 = N15;
  assign rs2_data_o = (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                      (N7)? rs2_reg_data : 1'b0;
  assign N6 = N21;
  assign N7 = N20;
  assign rs1_issue_v = issue_v_i & rs1_r_v_i;
  assign rs2_issue_v = issue_v_i & rs2_r_v_i;
  assign rs1_read_v = rs1_issue_v | N22;
  assign N22 = ~dispatch_v_i;
  assign rs2_read_v = rs2_issue_v | N22;
  assign N8 = ~rs1_issue_v;
  assign N9 = rs1_issue_v;
  assign N10 = ~rs2_issue_v;
  assign N11 = rs2_issue_v;

endmodule



module bsg_mem_2r1w_sync_synth_width_p64_els_p32_read_write_same_addr_p1_harden_p0
(
  clk_i,
  reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r0_v_i,
  r0_addr_i,
  r0_data_o,
  r1_v_i,
  r1_addr_i,
  r1_data_o
);

  input [4:0] w_addr_i;
  input [63:0] w_data_i;
  input [4:0] r0_addr_i;
  output [63:0] r0_data_o;
  input [4:0] r1_addr_i;
  output [63:0] r1_data_o;
  input clk_i;
  input reset_i;
  input w_v_i;
  input r0_v_i;
  input r1_v_i;
  wire [63:0] r0_data_o,r1_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221;
  reg [4:0] r0_addr_r,r1_addr_r;
  reg [2047:0] mem;
  assign r0_data_o[63] = (N43)? mem[63] :
                         (N45)? mem[127] :
                         (N47)? mem[191] :
                         (N49)? mem[255] :
                         (N51)? mem[319] :
                         (N53)? mem[383] :
                         (N55)? mem[447] :
                         (N57)? mem[511] :
                         (N59)? mem[575] :
                         (N61)? mem[639] :
                         (N63)? mem[703] :
                         (N65)? mem[767] :
                         (N67)? mem[831] :
                         (N69)? mem[895] :
                         (N71)? mem[959] :
                         (N73)? mem[1023] :
                         (N44)? mem[1087] :
                         (N46)? mem[1151] :
                         (N48)? mem[1215] :
                         (N50)? mem[1279] :
                         (N52)? mem[1343] :
                         (N54)? mem[1407] :
                         (N56)? mem[1471] :
                         (N58)? mem[1535] :
                         (N60)? mem[1599] :
                         (N62)? mem[1663] :
                         (N64)? mem[1727] :
                         (N66)? mem[1791] :
                         (N68)? mem[1855] :
                         (N70)? mem[1919] :
                         (N72)? mem[1983] :
                         (N74)? mem[2047] : 1'b0;
  assign r0_data_o[62] = (N43)? mem[62] :
                         (N45)? mem[126] :
                         (N47)? mem[190] :
                         (N49)? mem[254] :
                         (N51)? mem[318] :
                         (N53)? mem[382] :
                         (N55)? mem[446] :
                         (N57)? mem[510] :
                         (N59)? mem[574] :
                         (N61)? mem[638] :
                         (N63)? mem[702] :
                         (N65)? mem[766] :
                         (N67)? mem[830] :
                         (N69)? mem[894] :
                         (N71)? mem[958] :
                         (N73)? mem[1022] :
                         (N44)? mem[1086] :
                         (N46)? mem[1150] :
                         (N48)? mem[1214] :
                         (N50)? mem[1278] :
                         (N52)? mem[1342] :
                         (N54)? mem[1406] :
                         (N56)? mem[1470] :
                         (N58)? mem[1534] :
                         (N60)? mem[1598] :
                         (N62)? mem[1662] :
                         (N64)? mem[1726] :
                         (N66)? mem[1790] :
                         (N68)? mem[1854] :
                         (N70)? mem[1918] :
                         (N72)? mem[1982] :
                         (N74)? mem[2046] : 1'b0;
  assign r0_data_o[61] = (N43)? mem[61] :
                         (N45)? mem[125] :
                         (N47)? mem[189] :
                         (N49)? mem[253] :
                         (N51)? mem[317] :
                         (N53)? mem[381] :
                         (N55)? mem[445] :
                         (N57)? mem[509] :
                         (N59)? mem[573] :
                         (N61)? mem[637] :
                         (N63)? mem[701] :
                         (N65)? mem[765] :
                         (N67)? mem[829] :
                         (N69)? mem[893] :
                         (N71)? mem[957] :
                         (N73)? mem[1021] :
                         (N44)? mem[1085] :
                         (N46)? mem[1149] :
                         (N48)? mem[1213] :
                         (N50)? mem[1277] :
                         (N52)? mem[1341] :
                         (N54)? mem[1405] :
                         (N56)? mem[1469] :
                         (N58)? mem[1533] :
                         (N60)? mem[1597] :
                         (N62)? mem[1661] :
                         (N64)? mem[1725] :
                         (N66)? mem[1789] :
                         (N68)? mem[1853] :
                         (N70)? mem[1917] :
                         (N72)? mem[1981] :
                         (N74)? mem[2045] : 1'b0;
  assign r0_data_o[60] = (N43)? mem[60] :
                         (N45)? mem[124] :
                         (N47)? mem[188] :
                         (N49)? mem[252] :
                         (N51)? mem[316] :
                         (N53)? mem[380] :
                         (N55)? mem[444] :
                         (N57)? mem[508] :
                         (N59)? mem[572] :
                         (N61)? mem[636] :
                         (N63)? mem[700] :
                         (N65)? mem[764] :
                         (N67)? mem[828] :
                         (N69)? mem[892] :
                         (N71)? mem[956] :
                         (N73)? mem[1020] :
                         (N44)? mem[1084] :
                         (N46)? mem[1148] :
                         (N48)? mem[1212] :
                         (N50)? mem[1276] :
                         (N52)? mem[1340] :
                         (N54)? mem[1404] :
                         (N56)? mem[1468] :
                         (N58)? mem[1532] :
                         (N60)? mem[1596] :
                         (N62)? mem[1660] :
                         (N64)? mem[1724] :
                         (N66)? mem[1788] :
                         (N68)? mem[1852] :
                         (N70)? mem[1916] :
                         (N72)? mem[1980] :
                         (N74)? mem[2044] : 1'b0;
  assign r0_data_o[59] = (N43)? mem[59] :
                         (N45)? mem[123] :
                         (N47)? mem[187] :
                         (N49)? mem[251] :
                         (N51)? mem[315] :
                         (N53)? mem[379] :
                         (N55)? mem[443] :
                         (N57)? mem[507] :
                         (N59)? mem[571] :
                         (N61)? mem[635] :
                         (N63)? mem[699] :
                         (N65)? mem[763] :
                         (N67)? mem[827] :
                         (N69)? mem[891] :
                         (N71)? mem[955] :
                         (N73)? mem[1019] :
                         (N44)? mem[1083] :
                         (N46)? mem[1147] :
                         (N48)? mem[1211] :
                         (N50)? mem[1275] :
                         (N52)? mem[1339] :
                         (N54)? mem[1403] :
                         (N56)? mem[1467] :
                         (N58)? mem[1531] :
                         (N60)? mem[1595] :
                         (N62)? mem[1659] :
                         (N64)? mem[1723] :
                         (N66)? mem[1787] :
                         (N68)? mem[1851] :
                         (N70)? mem[1915] :
                         (N72)? mem[1979] :
                         (N74)? mem[2043] : 1'b0;
  assign r0_data_o[58] = (N43)? mem[58] :
                         (N45)? mem[122] :
                         (N47)? mem[186] :
                         (N49)? mem[250] :
                         (N51)? mem[314] :
                         (N53)? mem[378] :
                         (N55)? mem[442] :
                         (N57)? mem[506] :
                         (N59)? mem[570] :
                         (N61)? mem[634] :
                         (N63)? mem[698] :
                         (N65)? mem[762] :
                         (N67)? mem[826] :
                         (N69)? mem[890] :
                         (N71)? mem[954] :
                         (N73)? mem[1018] :
                         (N44)? mem[1082] :
                         (N46)? mem[1146] :
                         (N48)? mem[1210] :
                         (N50)? mem[1274] :
                         (N52)? mem[1338] :
                         (N54)? mem[1402] :
                         (N56)? mem[1466] :
                         (N58)? mem[1530] :
                         (N60)? mem[1594] :
                         (N62)? mem[1658] :
                         (N64)? mem[1722] :
                         (N66)? mem[1786] :
                         (N68)? mem[1850] :
                         (N70)? mem[1914] :
                         (N72)? mem[1978] :
                         (N74)? mem[2042] : 1'b0;
  assign r0_data_o[57] = (N43)? mem[57] :
                         (N45)? mem[121] :
                         (N47)? mem[185] :
                         (N49)? mem[249] :
                         (N51)? mem[313] :
                         (N53)? mem[377] :
                         (N55)? mem[441] :
                         (N57)? mem[505] :
                         (N59)? mem[569] :
                         (N61)? mem[633] :
                         (N63)? mem[697] :
                         (N65)? mem[761] :
                         (N67)? mem[825] :
                         (N69)? mem[889] :
                         (N71)? mem[953] :
                         (N73)? mem[1017] :
                         (N44)? mem[1081] :
                         (N46)? mem[1145] :
                         (N48)? mem[1209] :
                         (N50)? mem[1273] :
                         (N52)? mem[1337] :
                         (N54)? mem[1401] :
                         (N56)? mem[1465] :
                         (N58)? mem[1529] :
                         (N60)? mem[1593] :
                         (N62)? mem[1657] :
                         (N64)? mem[1721] :
                         (N66)? mem[1785] :
                         (N68)? mem[1849] :
                         (N70)? mem[1913] :
                         (N72)? mem[1977] :
                         (N74)? mem[2041] : 1'b0;
  assign r0_data_o[56] = (N43)? mem[56] :
                         (N45)? mem[120] :
                         (N47)? mem[184] :
                         (N49)? mem[248] :
                         (N51)? mem[312] :
                         (N53)? mem[376] :
                         (N55)? mem[440] :
                         (N57)? mem[504] :
                         (N59)? mem[568] :
                         (N61)? mem[632] :
                         (N63)? mem[696] :
                         (N65)? mem[760] :
                         (N67)? mem[824] :
                         (N69)? mem[888] :
                         (N71)? mem[952] :
                         (N73)? mem[1016] :
                         (N44)? mem[1080] :
                         (N46)? mem[1144] :
                         (N48)? mem[1208] :
                         (N50)? mem[1272] :
                         (N52)? mem[1336] :
                         (N54)? mem[1400] :
                         (N56)? mem[1464] :
                         (N58)? mem[1528] :
                         (N60)? mem[1592] :
                         (N62)? mem[1656] :
                         (N64)? mem[1720] :
                         (N66)? mem[1784] :
                         (N68)? mem[1848] :
                         (N70)? mem[1912] :
                         (N72)? mem[1976] :
                         (N74)? mem[2040] : 1'b0;
  assign r0_data_o[55] = (N43)? mem[55] :
                         (N45)? mem[119] :
                         (N47)? mem[183] :
                         (N49)? mem[247] :
                         (N51)? mem[311] :
                         (N53)? mem[375] :
                         (N55)? mem[439] :
                         (N57)? mem[503] :
                         (N59)? mem[567] :
                         (N61)? mem[631] :
                         (N63)? mem[695] :
                         (N65)? mem[759] :
                         (N67)? mem[823] :
                         (N69)? mem[887] :
                         (N71)? mem[951] :
                         (N73)? mem[1015] :
                         (N44)? mem[1079] :
                         (N46)? mem[1143] :
                         (N48)? mem[1207] :
                         (N50)? mem[1271] :
                         (N52)? mem[1335] :
                         (N54)? mem[1399] :
                         (N56)? mem[1463] :
                         (N58)? mem[1527] :
                         (N60)? mem[1591] :
                         (N62)? mem[1655] :
                         (N64)? mem[1719] :
                         (N66)? mem[1783] :
                         (N68)? mem[1847] :
                         (N70)? mem[1911] :
                         (N72)? mem[1975] :
                         (N74)? mem[2039] : 1'b0;
  assign r0_data_o[54] = (N43)? mem[54] :
                         (N45)? mem[118] :
                         (N47)? mem[182] :
                         (N49)? mem[246] :
                         (N51)? mem[310] :
                         (N53)? mem[374] :
                         (N55)? mem[438] :
                         (N57)? mem[502] :
                         (N59)? mem[566] :
                         (N61)? mem[630] :
                         (N63)? mem[694] :
                         (N65)? mem[758] :
                         (N67)? mem[822] :
                         (N69)? mem[886] :
                         (N71)? mem[950] :
                         (N73)? mem[1014] :
                         (N44)? mem[1078] :
                         (N46)? mem[1142] :
                         (N48)? mem[1206] :
                         (N50)? mem[1270] :
                         (N52)? mem[1334] :
                         (N54)? mem[1398] :
                         (N56)? mem[1462] :
                         (N58)? mem[1526] :
                         (N60)? mem[1590] :
                         (N62)? mem[1654] :
                         (N64)? mem[1718] :
                         (N66)? mem[1782] :
                         (N68)? mem[1846] :
                         (N70)? mem[1910] :
                         (N72)? mem[1974] :
                         (N74)? mem[2038] : 1'b0;
  assign r0_data_o[53] = (N43)? mem[53] :
                         (N45)? mem[117] :
                         (N47)? mem[181] :
                         (N49)? mem[245] :
                         (N51)? mem[309] :
                         (N53)? mem[373] :
                         (N55)? mem[437] :
                         (N57)? mem[501] :
                         (N59)? mem[565] :
                         (N61)? mem[629] :
                         (N63)? mem[693] :
                         (N65)? mem[757] :
                         (N67)? mem[821] :
                         (N69)? mem[885] :
                         (N71)? mem[949] :
                         (N73)? mem[1013] :
                         (N44)? mem[1077] :
                         (N46)? mem[1141] :
                         (N48)? mem[1205] :
                         (N50)? mem[1269] :
                         (N52)? mem[1333] :
                         (N54)? mem[1397] :
                         (N56)? mem[1461] :
                         (N58)? mem[1525] :
                         (N60)? mem[1589] :
                         (N62)? mem[1653] :
                         (N64)? mem[1717] :
                         (N66)? mem[1781] :
                         (N68)? mem[1845] :
                         (N70)? mem[1909] :
                         (N72)? mem[1973] :
                         (N74)? mem[2037] : 1'b0;
  assign r0_data_o[52] = (N43)? mem[52] :
                         (N45)? mem[116] :
                         (N47)? mem[180] :
                         (N49)? mem[244] :
                         (N51)? mem[308] :
                         (N53)? mem[372] :
                         (N55)? mem[436] :
                         (N57)? mem[500] :
                         (N59)? mem[564] :
                         (N61)? mem[628] :
                         (N63)? mem[692] :
                         (N65)? mem[756] :
                         (N67)? mem[820] :
                         (N69)? mem[884] :
                         (N71)? mem[948] :
                         (N73)? mem[1012] :
                         (N44)? mem[1076] :
                         (N46)? mem[1140] :
                         (N48)? mem[1204] :
                         (N50)? mem[1268] :
                         (N52)? mem[1332] :
                         (N54)? mem[1396] :
                         (N56)? mem[1460] :
                         (N58)? mem[1524] :
                         (N60)? mem[1588] :
                         (N62)? mem[1652] :
                         (N64)? mem[1716] :
                         (N66)? mem[1780] :
                         (N68)? mem[1844] :
                         (N70)? mem[1908] :
                         (N72)? mem[1972] :
                         (N74)? mem[2036] : 1'b0;
  assign r0_data_o[51] = (N43)? mem[51] :
                         (N45)? mem[115] :
                         (N47)? mem[179] :
                         (N49)? mem[243] :
                         (N51)? mem[307] :
                         (N53)? mem[371] :
                         (N55)? mem[435] :
                         (N57)? mem[499] :
                         (N59)? mem[563] :
                         (N61)? mem[627] :
                         (N63)? mem[691] :
                         (N65)? mem[755] :
                         (N67)? mem[819] :
                         (N69)? mem[883] :
                         (N71)? mem[947] :
                         (N73)? mem[1011] :
                         (N44)? mem[1075] :
                         (N46)? mem[1139] :
                         (N48)? mem[1203] :
                         (N50)? mem[1267] :
                         (N52)? mem[1331] :
                         (N54)? mem[1395] :
                         (N56)? mem[1459] :
                         (N58)? mem[1523] :
                         (N60)? mem[1587] :
                         (N62)? mem[1651] :
                         (N64)? mem[1715] :
                         (N66)? mem[1779] :
                         (N68)? mem[1843] :
                         (N70)? mem[1907] :
                         (N72)? mem[1971] :
                         (N74)? mem[2035] : 1'b0;
  assign r0_data_o[50] = (N43)? mem[50] :
                         (N45)? mem[114] :
                         (N47)? mem[178] :
                         (N49)? mem[242] :
                         (N51)? mem[306] :
                         (N53)? mem[370] :
                         (N55)? mem[434] :
                         (N57)? mem[498] :
                         (N59)? mem[562] :
                         (N61)? mem[626] :
                         (N63)? mem[690] :
                         (N65)? mem[754] :
                         (N67)? mem[818] :
                         (N69)? mem[882] :
                         (N71)? mem[946] :
                         (N73)? mem[1010] :
                         (N44)? mem[1074] :
                         (N46)? mem[1138] :
                         (N48)? mem[1202] :
                         (N50)? mem[1266] :
                         (N52)? mem[1330] :
                         (N54)? mem[1394] :
                         (N56)? mem[1458] :
                         (N58)? mem[1522] :
                         (N60)? mem[1586] :
                         (N62)? mem[1650] :
                         (N64)? mem[1714] :
                         (N66)? mem[1778] :
                         (N68)? mem[1842] :
                         (N70)? mem[1906] :
                         (N72)? mem[1970] :
                         (N74)? mem[2034] : 1'b0;
  assign r0_data_o[49] = (N43)? mem[49] :
                         (N45)? mem[113] :
                         (N47)? mem[177] :
                         (N49)? mem[241] :
                         (N51)? mem[305] :
                         (N53)? mem[369] :
                         (N55)? mem[433] :
                         (N57)? mem[497] :
                         (N59)? mem[561] :
                         (N61)? mem[625] :
                         (N63)? mem[689] :
                         (N65)? mem[753] :
                         (N67)? mem[817] :
                         (N69)? mem[881] :
                         (N71)? mem[945] :
                         (N73)? mem[1009] :
                         (N44)? mem[1073] :
                         (N46)? mem[1137] :
                         (N48)? mem[1201] :
                         (N50)? mem[1265] :
                         (N52)? mem[1329] :
                         (N54)? mem[1393] :
                         (N56)? mem[1457] :
                         (N58)? mem[1521] :
                         (N60)? mem[1585] :
                         (N62)? mem[1649] :
                         (N64)? mem[1713] :
                         (N66)? mem[1777] :
                         (N68)? mem[1841] :
                         (N70)? mem[1905] :
                         (N72)? mem[1969] :
                         (N74)? mem[2033] : 1'b0;
  assign r0_data_o[48] = (N43)? mem[48] :
                         (N45)? mem[112] :
                         (N47)? mem[176] :
                         (N49)? mem[240] :
                         (N51)? mem[304] :
                         (N53)? mem[368] :
                         (N55)? mem[432] :
                         (N57)? mem[496] :
                         (N59)? mem[560] :
                         (N61)? mem[624] :
                         (N63)? mem[688] :
                         (N65)? mem[752] :
                         (N67)? mem[816] :
                         (N69)? mem[880] :
                         (N71)? mem[944] :
                         (N73)? mem[1008] :
                         (N44)? mem[1072] :
                         (N46)? mem[1136] :
                         (N48)? mem[1200] :
                         (N50)? mem[1264] :
                         (N52)? mem[1328] :
                         (N54)? mem[1392] :
                         (N56)? mem[1456] :
                         (N58)? mem[1520] :
                         (N60)? mem[1584] :
                         (N62)? mem[1648] :
                         (N64)? mem[1712] :
                         (N66)? mem[1776] :
                         (N68)? mem[1840] :
                         (N70)? mem[1904] :
                         (N72)? mem[1968] :
                         (N74)? mem[2032] : 1'b0;
  assign r0_data_o[47] = (N43)? mem[47] :
                         (N45)? mem[111] :
                         (N47)? mem[175] :
                         (N49)? mem[239] :
                         (N51)? mem[303] :
                         (N53)? mem[367] :
                         (N55)? mem[431] :
                         (N57)? mem[495] :
                         (N59)? mem[559] :
                         (N61)? mem[623] :
                         (N63)? mem[687] :
                         (N65)? mem[751] :
                         (N67)? mem[815] :
                         (N69)? mem[879] :
                         (N71)? mem[943] :
                         (N73)? mem[1007] :
                         (N44)? mem[1071] :
                         (N46)? mem[1135] :
                         (N48)? mem[1199] :
                         (N50)? mem[1263] :
                         (N52)? mem[1327] :
                         (N54)? mem[1391] :
                         (N56)? mem[1455] :
                         (N58)? mem[1519] :
                         (N60)? mem[1583] :
                         (N62)? mem[1647] :
                         (N64)? mem[1711] :
                         (N66)? mem[1775] :
                         (N68)? mem[1839] :
                         (N70)? mem[1903] :
                         (N72)? mem[1967] :
                         (N74)? mem[2031] : 1'b0;
  assign r0_data_o[46] = (N43)? mem[46] :
                         (N45)? mem[110] :
                         (N47)? mem[174] :
                         (N49)? mem[238] :
                         (N51)? mem[302] :
                         (N53)? mem[366] :
                         (N55)? mem[430] :
                         (N57)? mem[494] :
                         (N59)? mem[558] :
                         (N61)? mem[622] :
                         (N63)? mem[686] :
                         (N65)? mem[750] :
                         (N67)? mem[814] :
                         (N69)? mem[878] :
                         (N71)? mem[942] :
                         (N73)? mem[1006] :
                         (N44)? mem[1070] :
                         (N46)? mem[1134] :
                         (N48)? mem[1198] :
                         (N50)? mem[1262] :
                         (N52)? mem[1326] :
                         (N54)? mem[1390] :
                         (N56)? mem[1454] :
                         (N58)? mem[1518] :
                         (N60)? mem[1582] :
                         (N62)? mem[1646] :
                         (N64)? mem[1710] :
                         (N66)? mem[1774] :
                         (N68)? mem[1838] :
                         (N70)? mem[1902] :
                         (N72)? mem[1966] :
                         (N74)? mem[2030] : 1'b0;
  assign r0_data_o[45] = (N43)? mem[45] :
                         (N45)? mem[109] :
                         (N47)? mem[173] :
                         (N49)? mem[237] :
                         (N51)? mem[301] :
                         (N53)? mem[365] :
                         (N55)? mem[429] :
                         (N57)? mem[493] :
                         (N59)? mem[557] :
                         (N61)? mem[621] :
                         (N63)? mem[685] :
                         (N65)? mem[749] :
                         (N67)? mem[813] :
                         (N69)? mem[877] :
                         (N71)? mem[941] :
                         (N73)? mem[1005] :
                         (N44)? mem[1069] :
                         (N46)? mem[1133] :
                         (N48)? mem[1197] :
                         (N50)? mem[1261] :
                         (N52)? mem[1325] :
                         (N54)? mem[1389] :
                         (N56)? mem[1453] :
                         (N58)? mem[1517] :
                         (N60)? mem[1581] :
                         (N62)? mem[1645] :
                         (N64)? mem[1709] :
                         (N66)? mem[1773] :
                         (N68)? mem[1837] :
                         (N70)? mem[1901] :
                         (N72)? mem[1965] :
                         (N74)? mem[2029] : 1'b0;
  assign r0_data_o[44] = (N43)? mem[44] :
                         (N45)? mem[108] :
                         (N47)? mem[172] :
                         (N49)? mem[236] :
                         (N51)? mem[300] :
                         (N53)? mem[364] :
                         (N55)? mem[428] :
                         (N57)? mem[492] :
                         (N59)? mem[556] :
                         (N61)? mem[620] :
                         (N63)? mem[684] :
                         (N65)? mem[748] :
                         (N67)? mem[812] :
                         (N69)? mem[876] :
                         (N71)? mem[940] :
                         (N73)? mem[1004] :
                         (N44)? mem[1068] :
                         (N46)? mem[1132] :
                         (N48)? mem[1196] :
                         (N50)? mem[1260] :
                         (N52)? mem[1324] :
                         (N54)? mem[1388] :
                         (N56)? mem[1452] :
                         (N58)? mem[1516] :
                         (N60)? mem[1580] :
                         (N62)? mem[1644] :
                         (N64)? mem[1708] :
                         (N66)? mem[1772] :
                         (N68)? mem[1836] :
                         (N70)? mem[1900] :
                         (N72)? mem[1964] :
                         (N74)? mem[2028] : 1'b0;
  assign r0_data_o[43] = (N43)? mem[43] :
                         (N45)? mem[107] :
                         (N47)? mem[171] :
                         (N49)? mem[235] :
                         (N51)? mem[299] :
                         (N53)? mem[363] :
                         (N55)? mem[427] :
                         (N57)? mem[491] :
                         (N59)? mem[555] :
                         (N61)? mem[619] :
                         (N63)? mem[683] :
                         (N65)? mem[747] :
                         (N67)? mem[811] :
                         (N69)? mem[875] :
                         (N71)? mem[939] :
                         (N73)? mem[1003] :
                         (N44)? mem[1067] :
                         (N46)? mem[1131] :
                         (N48)? mem[1195] :
                         (N50)? mem[1259] :
                         (N52)? mem[1323] :
                         (N54)? mem[1387] :
                         (N56)? mem[1451] :
                         (N58)? mem[1515] :
                         (N60)? mem[1579] :
                         (N62)? mem[1643] :
                         (N64)? mem[1707] :
                         (N66)? mem[1771] :
                         (N68)? mem[1835] :
                         (N70)? mem[1899] :
                         (N72)? mem[1963] :
                         (N74)? mem[2027] : 1'b0;
  assign r0_data_o[42] = (N43)? mem[42] :
                         (N45)? mem[106] :
                         (N47)? mem[170] :
                         (N49)? mem[234] :
                         (N51)? mem[298] :
                         (N53)? mem[362] :
                         (N55)? mem[426] :
                         (N57)? mem[490] :
                         (N59)? mem[554] :
                         (N61)? mem[618] :
                         (N63)? mem[682] :
                         (N65)? mem[746] :
                         (N67)? mem[810] :
                         (N69)? mem[874] :
                         (N71)? mem[938] :
                         (N73)? mem[1002] :
                         (N44)? mem[1066] :
                         (N46)? mem[1130] :
                         (N48)? mem[1194] :
                         (N50)? mem[1258] :
                         (N52)? mem[1322] :
                         (N54)? mem[1386] :
                         (N56)? mem[1450] :
                         (N58)? mem[1514] :
                         (N60)? mem[1578] :
                         (N62)? mem[1642] :
                         (N64)? mem[1706] :
                         (N66)? mem[1770] :
                         (N68)? mem[1834] :
                         (N70)? mem[1898] :
                         (N72)? mem[1962] :
                         (N74)? mem[2026] : 1'b0;
  assign r0_data_o[41] = (N43)? mem[41] :
                         (N45)? mem[105] :
                         (N47)? mem[169] :
                         (N49)? mem[233] :
                         (N51)? mem[297] :
                         (N53)? mem[361] :
                         (N55)? mem[425] :
                         (N57)? mem[489] :
                         (N59)? mem[553] :
                         (N61)? mem[617] :
                         (N63)? mem[681] :
                         (N65)? mem[745] :
                         (N67)? mem[809] :
                         (N69)? mem[873] :
                         (N71)? mem[937] :
                         (N73)? mem[1001] :
                         (N44)? mem[1065] :
                         (N46)? mem[1129] :
                         (N48)? mem[1193] :
                         (N50)? mem[1257] :
                         (N52)? mem[1321] :
                         (N54)? mem[1385] :
                         (N56)? mem[1449] :
                         (N58)? mem[1513] :
                         (N60)? mem[1577] :
                         (N62)? mem[1641] :
                         (N64)? mem[1705] :
                         (N66)? mem[1769] :
                         (N68)? mem[1833] :
                         (N70)? mem[1897] :
                         (N72)? mem[1961] :
                         (N74)? mem[2025] : 1'b0;
  assign r0_data_o[40] = (N43)? mem[40] :
                         (N45)? mem[104] :
                         (N47)? mem[168] :
                         (N49)? mem[232] :
                         (N51)? mem[296] :
                         (N53)? mem[360] :
                         (N55)? mem[424] :
                         (N57)? mem[488] :
                         (N59)? mem[552] :
                         (N61)? mem[616] :
                         (N63)? mem[680] :
                         (N65)? mem[744] :
                         (N67)? mem[808] :
                         (N69)? mem[872] :
                         (N71)? mem[936] :
                         (N73)? mem[1000] :
                         (N44)? mem[1064] :
                         (N46)? mem[1128] :
                         (N48)? mem[1192] :
                         (N50)? mem[1256] :
                         (N52)? mem[1320] :
                         (N54)? mem[1384] :
                         (N56)? mem[1448] :
                         (N58)? mem[1512] :
                         (N60)? mem[1576] :
                         (N62)? mem[1640] :
                         (N64)? mem[1704] :
                         (N66)? mem[1768] :
                         (N68)? mem[1832] :
                         (N70)? mem[1896] :
                         (N72)? mem[1960] :
                         (N74)? mem[2024] : 1'b0;
  assign r0_data_o[39] = (N43)? mem[39] :
                         (N45)? mem[103] :
                         (N47)? mem[167] :
                         (N49)? mem[231] :
                         (N51)? mem[295] :
                         (N53)? mem[359] :
                         (N55)? mem[423] :
                         (N57)? mem[487] :
                         (N59)? mem[551] :
                         (N61)? mem[615] :
                         (N63)? mem[679] :
                         (N65)? mem[743] :
                         (N67)? mem[807] :
                         (N69)? mem[871] :
                         (N71)? mem[935] :
                         (N73)? mem[999] :
                         (N44)? mem[1063] :
                         (N46)? mem[1127] :
                         (N48)? mem[1191] :
                         (N50)? mem[1255] :
                         (N52)? mem[1319] :
                         (N54)? mem[1383] :
                         (N56)? mem[1447] :
                         (N58)? mem[1511] :
                         (N60)? mem[1575] :
                         (N62)? mem[1639] :
                         (N64)? mem[1703] :
                         (N66)? mem[1767] :
                         (N68)? mem[1831] :
                         (N70)? mem[1895] :
                         (N72)? mem[1959] :
                         (N74)? mem[2023] : 1'b0;
  assign r0_data_o[38] = (N43)? mem[38] :
                         (N45)? mem[102] :
                         (N47)? mem[166] :
                         (N49)? mem[230] :
                         (N51)? mem[294] :
                         (N53)? mem[358] :
                         (N55)? mem[422] :
                         (N57)? mem[486] :
                         (N59)? mem[550] :
                         (N61)? mem[614] :
                         (N63)? mem[678] :
                         (N65)? mem[742] :
                         (N67)? mem[806] :
                         (N69)? mem[870] :
                         (N71)? mem[934] :
                         (N73)? mem[998] :
                         (N44)? mem[1062] :
                         (N46)? mem[1126] :
                         (N48)? mem[1190] :
                         (N50)? mem[1254] :
                         (N52)? mem[1318] :
                         (N54)? mem[1382] :
                         (N56)? mem[1446] :
                         (N58)? mem[1510] :
                         (N60)? mem[1574] :
                         (N62)? mem[1638] :
                         (N64)? mem[1702] :
                         (N66)? mem[1766] :
                         (N68)? mem[1830] :
                         (N70)? mem[1894] :
                         (N72)? mem[1958] :
                         (N74)? mem[2022] : 1'b0;
  assign r0_data_o[37] = (N43)? mem[37] :
                         (N45)? mem[101] :
                         (N47)? mem[165] :
                         (N49)? mem[229] :
                         (N51)? mem[293] :
                         (N53)? mem[357] :
                         (N55)? mem[421] :
                         (N57)? mem[485] :
                         (N59)? mem[549] :
                         (N61)? mem[613] :
                         (N63)? mem[677] :
                         (N65)? mem[741] :
                         (N67)? mem[805] :
                         (N69)? mem[869] :
                         (N71)? mem[933] :
                         (N73)? mem[997] :
                         (N44)? mem[1061] :
                         (N46)? mem[1125] :
                         (N48)? mem[1189] :
                         (N50)? mem[1253] :
                         (N52)? mem[1317] :
                         (N54)? mem[1381] :
                         (N56)? mem[1445] :
                         (N58)? mem[1509] :
                         (N60)? mem[1573] :
                         (N62)? mem[1637] :
                         (N64)? mem[1701] :
                         (N66)? mem[1765] :
                         (N68)? mem[1829] :
                         (N70)? mem[1893] :
                         (N72)? mem[1957] :
                         (N74)? mem[2021] : 1'b0;
  assign r0_data_o[36] = (N43)? mem[36] :
                         (N45)? mem[100] :
                         (N47)? mem[164] :
                         (N49)? mem[228] :
                         (N51)? mem[292] :
                         (N53)? mem[356] :
                         (N55)? mem[420] :
                         (N57)? mem[484] :
                         (N59)? mem[548] :
                         (N61)? mem[612] :
                         (N63)? mem[676] :
                         (N65)? mem[740] :
                         (N67)? mem[804] :
                         (N69)? mem[868] :
                         (N71)? mem[932] :
                         (N73)? mem[996] :
                         (N44)? mem[1060] :
                         (N46)? mem[1124] :
                         (N48)? mem[1188] :
                         (N50)? mem[1252] :
                         (N52)? mem[1316] :
                         (N54)? mem[1380] :
                         (N56)? mem[1444] :
                         (N58)? mem[1508] :
                         (N60)? mem[1572] :
                         (N62)? mem[1636] :
                         (N64)? mem[1700] :
                         (N66)? mem[1764] :
                         (N68)? mem[1828] :
                         (N70)? mem[1892] :
                         (N72)? mem[1956] :
                         (N74)? mem[2020] : 1'b0;
  assign r0_data_o[35] = (N43)? mem[35] :
                         (N45)? mem[99] :
                         (N47)? mem[163] :
                         (N49)? mem[227] :
                         (N51)? mem[291] :
                         (N53)? mem[355] :
                         (N55)? mem[419] :
                         (N57)? mem[483] :
                         (N59)? mem[547] :
                         (N61)? mem[611] :
                         (N63)? mem[675] :
                         (N65)? mem[739] :
                         (N67)? mem[803] :
                         (N69)? mem[867] :
                         (N71)? mem[931] :
                         (N73)? mem[995] :
                         (N44)? mem[1059] :
                         (N46)? mem[1123] :
                         (N48)? mem[1187] :
                         (N50)? mem[1251] :
                         (N52)? mem[1315] :
                         (N54)? mem[1379] :
                         (N56)? mem[1443] :
                         (N58)? mem[1507] :
                         (N60)? mem[1571] :
                         (N62)? mem[1635] :
                         (N64)? mem[1699] :
                         (N66)? mem[1763] :
                         (N68)? mem[1827] :
                         (N70)? mem[1891] :
                         (N72)? mem[1955] :
                         (N74)? mem[2019] : 1'b0;
  assign r0_data_o[34] = (N43)? mem[34] :
                         (N45)? mem[98] :
                         (N47)? mem[162] :
                         (N49)? mem[226] :
                         (N51)? mem[290] :
                         (N53)? mem[354] :
                         (N55)? mem[418] :
                         (N57)? mem[482] :
                         (N59)? mem[546] :
                         (N61)? mem[610] :
                         (N63)? mem[674] :
                         (N65)? mem[738] :
                         (N67)? mem[802] :
                         (N69)? mem[866] :
                         (N71)? mem[930] :
                         (N73)? mem[994] :
                         (N44)? mem[1058] :
                         (N46)? mem[1122] :
                         (N48)? mem[1186] :
                         (N50)? mem[1250] :
                         (N52)? mem[1314] :
                         (N54)? mem[1378] :
                         (N56)? mem[1442] :
                         (N58)? mem[1506] :
                         (N60)? mem[1570] :
                         (N62)? mem[1634] :
                         (N64)? mem[1698] :
                         (N66)? mem[1762] :
                         (N68)? mem[1826] :
                         (N70)? mem[1890] :
                         (N72)? mem[1954] :
                         (N74)? mem[2018] : 1'b0;
  assign r0_data_o[33] = (N43)? mem[33] :
                         (N45)? mem[97] :
                         (N47)? mem[161] :
                         (N49)? mem[225] :
                         (N51)? mem[289] :
                         (N53)? mem[353] :
                         (N55)? mem[417] :
                         (N57)? mem[481] :
                         (N59)? mem[545] :
                         (N61)? mem[609] :
                         (N63)? mem[673] :
                         (N65)? mem[737] :
                         (N67)? mem[801] :
                         (N69)? mem[865] :
                         (N71)? mem[929] :
                         (N73)? mem[993] :
                         (N44)? mem[1057] :
                         (N46)? mem[1121] :
                         (N48)? mem[1185] :
                         (N50)? mem[1249] :
                         (N52)? mem[1313] :
                         (N54)? mem[1377] :
                         (N56)? mem[1441] :
                         (N58)? mem[1505] :
                         (N60)? mem[1569] :
                         (N62)? mem[1633] :
                         (N64)? mem[1697] :
                         (N66)? mem[1761] :
                         (N68)? mem[1825] :
                         (N70)? mem[1889] :
                         (N72)? mem[1953] :
                         (N74)? mem[2017] : 1'b0;
  assign r0_data_o[32] = (N43)? mem[32] :
                         (N45)? mem[96] :
                         (N47)? mem[160] :
                         (N49)? mem[224] :
                         (N51)? mem[288] :
                         (N53)? mem[352] :
                         (N55)? mem[416] :
                         (N57)? mem[480] :
                         (N59)? mem[544] :
                         (N61)? mem[608] :
                         (N63)? mem[672] :
                         (N65)? mem[736] :
                         (N67)? mem[800] :
                         (N69)? mem[864] :
                         (N71)? mem[928] :
                         (N73)? mem[992] :
                         (N44)? mem[1056] :
                         (N46)? mem[1120] :
                         (N48)? mem[1184] :
                         (N50)? mem[1248] :
                         (N52)? mem[1312] :
                         (N54)? mem[1376] :
                         (N56)? mem[1440] :
                         (N58)? mem[1504] :
                         (N60)? mem[1568] :
                         (N62)? mem[1632] :
                         (N64)? mem[1696] :
                         (N66)? mem[1760] :
                         (N68)? mem[1824] :
                         (N70)? mem[1888] :
                         (N72)? mem[1952] :
                         (N74)? mem[2016] : 1'b0;
  assign r0_data_o[31] = (N43)? mem[31] :
                         (N45)? mem[95] :
                         (N47)? mem[159] :
                         (N49)? mem[223] :
                         (N51)? mem[287] :
                         (N53)? mem[351] :
                         (N55)? mem[415] :
                         (N57)? mem[479] :
                         (N59)? mem[543] :
                         (N61)? mem[607] :
                         (N63)? mem[671] :
                         (N65)? mem[735] :
                         (N67)? mem[799] :
                         (N69)? mem[863] :
                         (N71)? mem[927] :
                         (N73)? mem[991] :
                         (N44)? mem[1055] :
                         (N46)? mem[1119] :
                         (N48)? mem[1183] :
                         (N50)? mem[1247] :
                         (N52)? mem[1311] :
                         (N54)? mem[1375] :
                         (N56)? mem[1439] :
                         (N58)? mem[1503] :
                         (N60)? mem[1567] :
                         (N62)? mem[1631] :
                         (N64)? mem[1695] :
                         (N66)? mem[1759] :
                         (N68)? mem[1823] :
                         (N70)? mem[1887] :
                         (N72)? mem[1951] :
                         (N74)? mem[2015] : 1'b0;
  assign r0_data_o[30] = (N43)? mem[30] :
                         (N45)? mem[94] :
                         (N47)? mem[158] :
                         (N49)? mem[222] :
                         (N51)? mem[286] :
                         (N53)? mem[350] :
                         (N55)? mem[414] :
                         (N57)? mem[478] :
                         (N59)? mem[542] :
                         (N61)? mem[606] :
                         (N63)? mem[670] :
                         (N65)? mem[734] :
                         (N67)? mem[798] :
                         (N69)? mem[862] :
                         (N71)? mem[926] :
                         (N73)? mem[990] :
                         (N44)? mem[1054] :
                         (N46)? mem[1118] :
                         (N48)? mem[1182] :
                         (N50)? mem[1246] :
                         (N52)? mem[1310] :
                         (N54)? mem[1374] :
                         (N56)? mem[1438] :
                         (N58)? mem[1502] :
                         (N60)? mem[1566] :
                         (N62)? mem[1630] :
                         (N64)? mem[1694] :
                         (N66)? mem[1758] :
                         (N68)? mem[1822] :
                         (N70)? mem[1886] :
                         (N72)? mem[1950] :
                         (N74)? mem[2014] : 1'b0;
  assign r0_data_o[29] = (N43)? mem[29] :
                         (N45)? mem[93] :
                         (N47)? mem[157] :
                         (N49)? mem[221] :
                         (N51)? mem[285] :
                         (N53)? mem[349] :
                         (N55)? mem[413] :
                         (N57)? mem[477] :
                         (N59)? mem[541] :
                         (N61)? mem[605] :
                         (N63)? mem[669] :
                         (N65)? mem[733] :
                         (N67)? mem[797] :
                         (N69)? mem[861] :
                         (N71)? mem[925] :
                         (N73)? mem[989] :
                         (N44)? mem[1053] :
                         (N46)? mem[1117] :
                         (N48)? mem[1181] :
                         (N50)? mem[1245] :
                         (N52)? mem[1309] :
                         (N54)? mem[1373] :
                         (N56)? mem[1437] :
                         (N58)? mem[1501] :
                         (N60)? mem[1565] :
                         (N62)? mem[1629] :
                         (N64)? mem[1693] :
                         (N66)? mem[1757] :
                         (N68)? mem[1821] :
                         (N70)? mem[1885] :
                         (N72)? mem[1949] :
                         (N74)? mem[2013] : 1'b0;
  assign r0_data_o[28] = (N43)? mem[28] :
                         (N45)? mem[92] :
                         (N47)? mem[156] :
                         (N49)? mem[220] :
                         (N51)? mem[284] :
                         (N53)? mem[348] :
                         (N55)? mem[412] :
                         (N57)? mem[476] :
                         (N59)? mem[540] :
                         (N61)? mem[604] :
                         (N63)? mem[668] :
                         (N65)? mem[732] :
                         (N67)? mem[796] :
                         (N69)? mem[860] :
                         (N71)? mem[924] :
                         (N73)? mem[988] :
                         (N44)? mem[1052] :
                         (N46)? mem[1116] :
                         (N48)? mem[1180] :
                         (N50)? mem[1244] :
                         (N52)? mem[1308] :
                         (N54)? mem[1372] :
                         (N56)? mem[1436] :
                         (N58)? mem[1500] :
                         (N60)? mem[1564] :
                         (N62)? mem[1628] :
                         (N64)? mem[1692] :
                         (N66)? mem[1756] :
                         (N68)? mem[1820] :
                         (N70)? mem[1884] :
                         (N72)? mem[1948] :
                         (N74)? mem[2012] : 1'b0;
  assign r0_data_o[27] = (N43)? mem[27] :
                         (N45)? mem[91] :
                         (N47)? mem[155] :
                         (N49)? mem[219] :
                         (N51)? mem[283] :
                         (N53)? mem[347] :
                         (N55)? mem[411] :
                         (N57)? mem[475] :
                         (N59)? mem[539] :
                         (N61)? mem[603] :
                         (N63)? mem[667] :
                         (N65)? mem[731] :
                         (N67)? mem[795] :
                         (N69)? mem[859] :
                         (N71)? mem[923] :
                         (N73)? mem[987] :
                         (N44)? mem[1051] :
                         (N46)? mem[1115] :
                         (N48)? mem[1179] :
                         (N50)? mem[1243] :
                         (N52)? mem[1307] :
                         (N54)? mem[1371] :
                         (N56)? mem[1435] :
                         (N58)? mem[1499] :
                         (N60)? mem[1563] :
                         (N62)? mem[1627] :
                         (N64)? mem[1691] :
                         (N66)? mem[1755] :
                         (N68)? mem[1819] :
                         (N70)? mem[1883] :
                         (N72)? mem[1947] :
                         (N74)? mem[2011] : 1'b0;
  assign r0_data_o[26] = (N43)? mem[26] :
                         (N45)? mem[90] :
                         (N47)? mem[154] :
                         (N49)? mem[218] :
                         (N51)? mem[282] :
                         (N53)? mem[346] :
                         (N55)? mem[410] :
                         (N57)? mem[474] :
                         (N59)? mem[538] :
                         (N61)? mem[602] :
                         (N63)? mem[666] :
                         (N65)? mem[730] :
                         (N67)? mem[794] :
                         (N69)? mem[858] :
                         (N71)? mem[922] :
                         (N73)? mem[986] :
                         (N44)? mem[1050] :
                         (N46)? mem[1114] :
                         (N48)? mem[1178] :
                         (N50)? mem[1242] :
                         (N52)? mem[1306] :
                         (N54)? mem[1370] :
                         (N56)? mem[1434] :
                         (N58)? mem[1498] :
                         (N60)? mem[1562] :
                         (N62)? mem[1626] :
                         (N64)? mem[1690] :
                         (N66)? mem[1754] :
                         (N68)? mem[1818] :
                         (N70)? mem[1882] :
                         (N72)? mem[1946] :
                         (N74)? mem[2010] : 1'b0;
  assign r0_data_o[25] = (N43)? mem[25] :
                         (N45)? mem[89] :
                         (N47)? mem[153] :
                         (N49)? mem[217] :
                         (N51)? mem[281] :
                         (N53)? mem[345] :
                         (N55)? mem[409] :
                         (N57)? mem[473] :
                         (N59)? mem[537] :
                         (N61)? mem[601] :
                         (N63)? mem[665] :
                         (N65)? mem[729] :
                         (N67)? mem[793] :
                         (N69)? mem[857] :
                         (N71)? mem[921] :
                         (N73)? mem[985] :
                         (N44)? mem[1049] :
                         (N46)? mem[1113] :
                         (N48)? mem[1177] :
                         (N50)? mem[1241] :
                         (N52)? mem[1305] :
                         (N54)? mem[1369] :
                         (N56)? mem[1433] :
                         (N58)? mem[1497] :
                         (N60)? mem[1561] :
                         (N62)? mem[1625] :
                         (N64)? mem[1689] :
                         (N66)? mem[1753] :
                         (N68)? mem[1817] :
                         (N70)? mem[1881] :
                         (N72)? mem[1945] :
                         (N74)? mem[2009] : 1'b0;
  assign r0_data_o[24] = (N43)? mem[24] :
                         (N45)? mem[88] :
                         (N47)? mem[152] :
                         (N49)? mem[216] :
                         (N51)? mem[280] :
                         (N53)? mem[344] :
                         (N55)? mem[408] :
                         (N57)? mem[472] :
                         (N59)? mem[536] :
                         (N61)? mem[600] :
                         (N63)? mem[664] :
                         (N65)? mem[728] :
                         (N67)? mem[792] :
                         (N69)? mem[856] :
                         (N71)? mem[920] :
                         (N73)? mem[984] :
                         (N44)? mem[1048] :
                         (N46)? mem[1112] :
                         (N48)? mem[1176] :
                         (N50)? mem[1240] :
                         (N52)? mem[1304] :
                         (N54)? mem[1368] :
                         (N56)? mem[1432] :
                         (N58)? mem[1496] :
                         (N60)? mem[1560] :
                         (N62)? mem[1624] :
                         (N64)? mem[1688] :
                         (N66)? mem[1752] :
                         (N68)? mem[1816] :
                         (N70)? mem[1880] :
                         (N72)? mem[1944] :
                         (N74)? mem[2008] : 1'b0;
  assign r0_data_o[23] = (N43)? mem[23] :
                         (N45)? mem[87] :
                         (N47)? mem[151] :
                         (N49)? mem[215] :
                         (N51)? mem[279] :
                         (N53)? mem[343] :
                         (N55)? mem[407] :
                         (N57)? mem[471] :
                         (N59)? mem[535] :
                         (N61)? mem[599] :
                         (N63)? mem[663] :
                         (N65)? mem[727] :
                         (N67)? mem[791] :
                         (N69)? mem[855] :
                         (N71)? mem[919] :
                         (N73)? mem[983] :
                         (N44)? mem[1047] :
                         (N46)? mem[1111] :
                         (N48)? mem[1175] :
                         (N50)? mem[1239] :
                         (N52)? mem[1303] :
                         (N54)? mem[1367] :
                         (N56)? mem[1431] :
                         (N58)? mem[1495] :
                         (N60)? mem[1559] :
                         (N62)? mem[1623] :
                         (N64)? mem[1687] :
                         (N66)? mem[1751] :
                         (N68)? mem[1815] :
                         (N70)? mem[1879] :
                         (N72)? mem[1943] :
                         (N74)? mem[2007] : 1'b0;
  assign r0_data_o[22] = (N43)? mem[22] :
                         (N45)? mem[86] :
                         (N47)? mem[150] :
                         (N49)? mem[214] :
                         (N51)? mem[278] :
                         (N53)? mem[342] :
                         (N55)? mem[406] :
                         (N57)? mem[470] :
                         (N59)? mem[534] :
                         (N61)? mem[598] :
                         (N63)? mem[662] :
                         (N65)? mem[726] :
                         (N67)? mem[790] :
                         (N69)? mem[854] :
                         (N71)? mem[918] :
                         (N73)? mem[982] :
                         (N44)? mem[1046] :
                         (N46)? mem[1110] :
                         (N48)? mem[1174] :
                         (N50)? mem[1238] :
                         (N52)? mem[1302] :
                         (N54)? mem[1366] :
                         (N56)? mem[1430] :
                         (N58)? mem[1494] :
                         (N60)? mem[1558] :
                         (N62)? mem[1622] :
                         (N64)? mem[1686] :
                         (N66)? mem[1750] :
                         (N68)? mem[1814] :
                         (N70)? mem[1878] :
                         (N72)? mem[1942] :
                         (N74)? mem[2006] : 1'b0;
  assign r0_data_o[21] = (N43)? mem[21] :
                         (N45)? mem[85] :
                         (N47)? mem[149] :
                         (N49)? mem[213] :
                         (N51)? mem[277] :
                         (N53)? mem[341] :
                         (N55)? mem[405] :
                         (N57)? mem[469] :
                         (N59)? mem[533] :
                         (N61)? mem[597] :
                         (N63)? mem[661] :
                         (N65)? mem[725] :
                         (N67)? mem[789] :
                         (N69)? mem[853] :
                         (N71)? mem[917] :
                         (N73)? mem[981] :
                         (N44)? mem[1045] :
                         (N46)? mem[1109] :
                         (N48)? mem[1173] :
                         (N50)? mem[1237] :
                         (N52)? mem[1301] :
                         (N54)? mem[1365] :
                         (N56)? mem[1429] :
                         (N58)? mem[1493] :
                         (N60)? mem[1557] :
                         (N62)? mem[1621] :
                         (N64)? mem[1685] :
                         (N66)? mem[1749] :
                         (N68)? mem[1813] :
                         (N70)? mem[1877] :
                         (N72)? mem[1941] :
                         (N74)? mem[2005] : 1'b0;
  assign r0_data_o[20] = (N43)? mem[20] :
                         (N45)? mem[84] :
                         (N47)? mem[148] :
                         (N49)? mem[212] :
                         (N51)? mem[276] :
                         (N53)? mem[340] :
                         (N55)? mem[404] :
                         (N57)? mem[468] :
                         (N59)? mem[532] :
                         (N61)? mem[596] :
                         (N63)? mem[660] :
                         (N65)? mem[724] :
                         (N67)? mem[788] :
                         (N69)? mem[852] :
                         (N71)? mem[916] :
                         (N73)? mem[980] :
                         (N44)? mem[1044] :
                         (N46)? mem[1108] :
                         (N48)? mem[1172] :
                         (N50)? mem[1236] :
                         (N52)? mem[1300] :
                         (N54)? mem[1364] :
                         (N56)? mem[1428] :
                         (N58)? mem[1492] :
                         (N60)? mem[1556] :
                         (N62)? mem[1620] :
                         (N64)? mem[1684] :
                         (N66)? mem[1748] :
                         (N68)? mem[1812] :
                         (N70)? mem[1876] :
                         (N72)? mem[1940] :
                         (N74)? mem[2004] : 1'b0;
  assign r0_data_o[19] = (N43)? mem[19] :
                         (N45)? mem[83] :
                         (N47)? mem[147] :
                         (N49)? mem[211] :
                         (N51)? mem[275] :
                         (N53)? mem[339] :
                         (N55)? mem[403] :
                         (N57)? mem[467] :
                         (N59)? mem[531] :
                         (N61)? mem[595] :
                         (N63)? mem[659] :
                         (N65)? mem[723] :
                         (N67)? mem[787] :
                         (N69)? mem[851] :
                         (N71)? mem[915] :
                         (N73)? mem[979] :
                         (N44)? mem[1043] :
                         (N46)? mem[1107] :
                         (N48)? mem[1171] :
                         (N50)? mem[1235] :
                         (N52)? mem[1299] :
                         (N54)? mem[1363] :
                         (N56)? mem[1427] :
                         (N58)? mem[1491] :
                         (N60)? mem[1555] :
                         (N62)? mem[1619] :
                         (N64)? mem[1683] :
                         (N66)? mem[1747] :
                         (N68)? mem[1811] :
                         (N70)? mem[1875] :
                         (N72)? mem[1939] :
                         (N74)? mem[2003] : 1'b0;
  assign r0_data_o[18] = (N43)? mem[18] :
                         (N45)? mem[82] :
                         (N47)? mem[146] :
                         (N49)? mem[210] :
                         (N51)? mem[274] :
                         (N53)? mem[338] :
                         (N55)? mem[402] :
                         (N57)? mem[466] :
                         (N59)? mem[530] :
                         (N61)? mem[594] :
                         (N63)? mem[658] :
                         (N65)? mem[722] :
                         (N67)? mem[786] :
                         (N69)? mem[850] :
                         (N71)? mem[914] :
                         (N73)? mem[978] :
                         (N44)? mem[1042] :
                         (N46)? mem[1106] :
                         (N48)? mem[1170] :
                         (N50)? mem[1234] :
                         (N52)? mem[1298] :
                         (N54)? mem[1362] :
                         (N56)? mem[1426] :
                         (N58)? mem[1490] :
                         (N60)? mem[1554] :
                         (N62)? mem[1618] :
                         (N64)? mem[1682] :
                         (N66)? mem[1746] :
                         (N68)? mem[1810] :
                         (N70)? mem[1874] :
                         (N72)? mem[1938] :
                         (N74)? mem[2002] : 1'b0;
  assign r0_data_o[17] = (N43)? mem[17] :
                         (N45)? mem[81] :
                         (N47)? mem[145] :
                         (N49)? mem[209] :
                         (N51)? mem[273] :
                         (N53)? mem[337] :
                         (N55)? mem[401] :
                         (N57)? mem[465] :
                         (N59)? mem[529] :
                         (N61)? mem[593] :
                         (N63)? mem[657] :
                         (N65)? mem[721] :
                         (N67)? mem[785] :
                         (N69)? mem[849] :
                         (N71)? mem[913] :
                         (N73)? mem[977] :
                         (N44)? mem[1041] :
                         (N46)? mem[1105] :
                         (N48)? mem[1169] :
                         (N50)? mem[1233] :
                         (N52)? mem[1297] :
                         (N54)? mem[1361] :
                         (N56)? mem[1425] :
                         (N58)? mem[1489] :
                         (N60)? mem[1553] :
                         (N62)? mem[1617] :
                         (N64)? mem[1681] :
                         (N66)? mem[1745] :
                         (N68)? mem[1809] :
                         (N70)? mem[1873] :
                         (N72)? mem[1937] :
                         (N74)? mem[2001] : 1'b0;
  assign r0_data_o[16] = (N43)? mem[16] :
                         (N45)? mem[80] :
                         (N47)? mem[144] :
                         (N49)? mem[208] :
                         (N51)? mem[272] :
                         (N53)? mem[336] :
                         (N55)? mem[400] :
                         (N57)? mem[464] :
                         (N59)? mem[528] :
                         (N61)? mem[592] :
                         (N63)? mem[656] :
                         (N65)? mem[720] :
                         (N67)? mem[784] :
                         (N69)? mem[848] :
                         (N71)? mem[912] :
                         (N73)? mem[976] :
                         (N44)? mem[1040] :
                         (N46)? mem[1104] :
                         (N48)? mem[1168] :
                         (N50)? mem[1232] :
                         (N52)? mem[1296] :
                         (N54)? mem[1360] :
                         (N56)? mem[1424] :
                         (N58)? mem[1488] :
                         (N60)? mem[1552] :
                         (N62)? mem[1616] :
                         (N64)? mem[1680] :
                         (N66)? mem[1744] :
                         (N68)? mem[1808] :
                         (N70)? mem[1872] :
                         (N72)? mem[1936] :
                         (N74)? mem[2000] : 1'b0;
  assign r0_data_o[15] = (N43)? mem[15] :
                         (N45)? mem[79] :
                         (N47)? mem[143] :
                         (N49)? mem[207] :
                         (N51)? mem[271] :
                         (N53)? mem[335] :
                         (N55)? mem[399] :
                         (N57)? mem[463] :
                         (N59)? mem[527] :
                         (N61)? mem[591] :
                         (N63)? mem[655] :
                         (N65)? mem[719] :
                         (N67)? mem[783] :
                         (N69)? mem[847] :
                         (N71)? mem[911] :
                         (N73)? mem[975] :
                         (N44)? mem[1039] :
                         (N46)? mem[1103] :
                         (N48)? mem[1167] :
                         (N50)? mem[1231] :
                         (N52)? mem[1295] :
                         (N54)? mem[1359] :
                         (N56)? mem[1423] :
                         (N58)? mem[1487] :
                         (N60)? mem[1551] :
                         (N62)? mem[1615] :
                         (N64)? mem[1679] :
                         (N66)? mem[1743] :
                         (N68)? mem[1807] :
                         (N70)? mem[1871] :
                         (N72)? mem[1935] :
                         (N74)? mem[1999] : 1'b0;
  assign r0_data_o[14] = (N43)? mem[14] :
                         (N45)? mem[78] :
                         (N47)? mem[142] :
                         (N49)? mem[206] :
                         (N51)? mem[270] :
                         (N53)? mem[334] :
                         (N55)? mem[398] :
                         (N57)? mem[462] :
                         (N59)? mem[526] :
                         (N61)? mem[590] :
                         (N63)? mem[654] :
                         (N65)? mem[718] :
                         (N67)? mem[782] :
                         (N69)? mem[846] :
                         (N71)? mem[910] :
                         (N73)? mem[974] :
                         (N44)? mem[1038] :
                         (N46)? mem[1102] :
                         (N48)? mem[1166] :
                         (N50)? mem[1230] :
                         (N52)? mem[1294] :
                         (N54)? mem[1358] :
                         (N56)? mem[1422] :
                         (N58)? mem[1486] :
                         (N60)? mem[1550] :
                         (N62)? mem[1614] :
                         (N64)? mem[1678] :
                         (N66)? mem[1742] :
                         (N68)? mem[1806] :
                         (N70)? mem[1870] :
                         (N72)? mem[1934] :
                         (N74)? mem[1998] : 1'b0;
  assign r0_data_o[13] = (N43)? mem[13] :
                         (N45)? mem[77] :
                         (N47)? mem[141] :
                         (N49)? mem[205] :
                         (N51)? mem[269] :
                         (N53)? mem[333] :
                         (N55)? mem[397] :
                         (N57)? mem[461] :
                         (N59)? mem[525] :
                         (N61)? mem[589] :
                         (N63)? mem[653] :
                         (N65)? mem[717] :
                         (N67)? mem[781] :
                         (N69)? mem[845] :
                         (N71)? mem[909] :
                         (N73)? mem[973] :
                         (N44)? mem[1037] :
                         (N46)? mem[1101] :
                         (N48)? mem[1165] :
                         (N50)? mem[1229] :
                         (N52)? mem[1293] :
                         (N54)? mem[1357] :
                         (N56)? mem[1421] :
                         (N58)? mem[1485] :
                         (N60)? mem[1549] :
                         (N62)? mem[1613] :
                         (N64)? mem[1677] :
                         (N66)? mem[1741] :
                         (N68)? mem[1805] :
                         (N70)? mem[1869] :
                         (N72)? mem[1933] :
                         (N74)? mem[1997] : 1'b0;
  assign r0_data_o[12] = (N43)? mem[12] :
                         (N45)? mem[76] :
                         (N47)? mem[140] :
                         (N49)? mem[204] :
                         (N51)? mem[268] :
                         (N53)? mem[332] :
                         (N55)? mem[396] :
                         (N57)? mem[460] :
                         (N59)? mem[524] :
                         (N61)? mem[588] :
                         (N63)? mem[652] :
                         (N65)? mem[716] :
                         (N67)? mem[780] :
                         (N69)? mem[844] :
                         (N71)? mem[908] :
                         (N73)? mem[972] :
                         (N44)? mem[1036] :
                         (N46)? mem[1100] :
                         (N48)? mem[1164] :
                         (N50)? mem[1228] :
                         (N52)? mem[1292] :
                         (N54)? mem[1356] :
                         (N56)? mem[1420] :
                         (N58)? mem[1484] :
                         (N60)? mem[1548] :
                         (N62)? mem[1612] :
                         (N64)? mem[1676] :
                         (N66)? mem[1740] :
                         (N68)? mem[1804] :
                         (N70)? mem[1868] :
                         (N72)? mem[1932] :
                         (N74)? mem[1996] : 1'b0;
  assign r0_data_o[11] = (N43)? mem[11] :
                         (N45)? mem[75] :
                         (N47)? mem[139] :
                         (N49)? mem[203] :
                         (N51)? mem[267] :
                         (N53)? mem[331] :
                         (N55)? mem[395] :
                         (N57)? mem[459] :
                         (N59)? mem[523] :
                         (N61)? mem[587] :
                         (N63)? mem[651] :
                         (N65)? mem[715] :
                         (N67)? mem[779] :
                         (N69)? mem[843] :
                         (N71)? mem[907] :
                         (N73)? mem[971] :
                         (N44)? mem[1035] :
                         (N46)? mem[1099] :
                         (N48)? mem[1163] :
                         (N50)? mem[1227] :
                         (N52)? mem[1291] :
                         (N54)? mem[1355] :
                         (N56)? mem[1419] :
                         (N58)? mem[1483] :
                         (N60)? mem[1547] :
                         (N62)? mem[1611] :
                         (N64)? mem[1675] :
                         (N66)? mem[1739] :
                         (N68)? mem[1803] :
                         (N70)? mem[1867] :
                         (N72)? mem[1931] :
                         (N74)? mem[1995] : 1'b0;
  assign r0_data_o[10] = (N43)? mem[10] :
                         (N45)? mem[74] :
                         (N47)? mem[138] :
                         (N49)? mem[202] :
                         (N51)? mem[266] :
                         (N53)? mem[330] :
                         (N55)? mem[394] :
                         (N57)? mem[458] :
                         (N59)? mem[522] :
                         (N61)? mem[586] :
                         (N63)? mem[650] :
                         (N65)? mem[714] :
                         (N67)? mem[778] :
                         (N69)? mem[842] :
                         (N71)? mem[906] :
                         (N73)? mem[970] :
                         (N44)? mem[1034] :
                         (N46)? mem[1098] :
                         (N48)? mem[1162] :
                         (N50)? mem[1226] :
                         (N52)? mem[1290] :
                         (N54)? mem[1354] :
                         (N56)? mem[1418] :
                         (N58)? mem[1482] :
                         (N60)? mem[1546] :
                         (N62)? mem[1610] :
                         (N64)? mem[1674] :
                         (N66)? mem[1738] :
                         (N68)? mem[1802] :
                         (N70)? mem[1866] :
                         (N72)? mem[1930] :
                         (N74)? mem[1994] : 1'b0;
  assign r0_data_o[9] = (N43)? mem[9] :
                        (N45)? mem[73] :
                        (N47)? mem[137] :
                        (N49)? mem[201] :
                        (N51)? mem[265] :
                        (N53)? mem[329] :
                        (N55)? mem[393] :
                        (N57)? mem[457] :
                        (N59)? mem[521] :
                        (N61)? mem[585] :
                        (N63)? mem[649] :
                        (N65)? mem[713] :
                        (N67)? mem[777] :
                        (N69)? mem[841] :
                        (N71)? mem[905] :
                        (N73)? mem[969] :
                        (N44)? mem[1033] :
                        (N46)? mem[1097] :
                        (N48)? mem[1161] :
                        (N50)? mem[1225] :
                        (N52)? mem[1289] :
                        (N54)? mem[1353] :
                        (N56)? mem[1417] :
                        (N58)? mem[1481] :
                        (N60)? mem[1545] :
                        (N62)? mem[1609] :
                        (N64)? mem[1673] :
                        (N66)? mem[1737] :
                        (N68)? mem[1801] :
                        (N70)? mem[1865] :
                        (N72)? mem[1929] :
                        (N74)? mem[1993] : 1'b0;
  assign r0_data_o[8] = (N43)? mem[8] :
                        (N45)? mem[72] :
                        (N47)? mem[136] :
                        (N49)? mem[200] :
                        (N51)? mem[264] :
                        (N53)? mem[328] :
                        (N55)? mem[392] :
                        (N57)? mem[456] :
                        (N59)? mem[520] :
                        (N61)? mem[584] :
                        (N63)? mem[648] :
                        (N65)? mem[712] :
                        (N67)? mem[776] :
                        (N69)? mem[840] :
                        (N71)? mem[904] :
                        (N73)? mem[968] :
                        (N44)? mem[1032] :
                        (N46)? mem[1096] :
                        (N48)? mem[1160] :
                        (N50)? mem[1224] :
                        (N52)? mem[1288] :
                        (N54)? mem[1352] :
                        (N56)? mem[1416] :
                        (N58)? mem[1480] :
                        (N60)? mem[1544] :
                        (N62)? mem[1608] :
                        (N64)? mem[1672] :
                        (N66)? mem[1736] :
                        (N68)? mem[1800] :
                        (N70)? mem[1864] :
                        (N72)? mem[1928] :
                        (N74)? mem[1992] : 1'b0;
  assign r0_data_o[7] = (N43)? mem[7] :
                        (N45)? mem[71] :
                        (N47)? mem[135] :
                        (N49)? mem[199] :
                        (N51)? mem[263] :
                        (N53)? mem[327] :
                        (N55)? mem[391] :
                        (N57)? mem[455] :
                        (N59)? mem[519] :
                        (N61)? mem[583] :
                        (N63)? mem[647] :
                        (N65)? mem[711] :
                        (N67)? mem[775] :
                        (N69)? mem[839] :
                        (N71)? mem[903] :
                        (N73)? mem[967] :
                        (N44)? mem[1031] :
                        (N46)? mem[1095] :
                        (N48)? mem[1159] :
                        (N50)? mem[1223] :
                        (N52)? mem[1287] :
                        (N54)? mem[1351] :
                        (N56)? mem[1415] :
                        (N58)? mem[1479] :
                        (N60)? mem[1543] :
                        (N62)? mem[1607] :
                        (N64)? mem[1671] :
                        (N66)? mem[1735] :
                        (N68)? mem[1799] :
                        (N70)? mem[1863] :
                        (N72)? mem[1927] :
                        (N74)? mem[1991] : 1'b0;
  assign r0_data_o[6] = (N43)? mem[6] :
                        (N45)? mem[70] :
                        (N47)? mem[134] :
                        (N49)? mem[198] :
                        (N51)? mem[262] :
                        (N53)? mem[326] :
                        (N55)? mem[390] :
                        (N57)? mem[454] :
                        (N59)? mem[518] :
                        (N61)? mem[582] :
                        (N63)? mem[646] :
                        (N65)? mem[710] :
                        (N67)? mem[774] :
                        (N69)? mem[838] :
                        (N71)? mem[902] :
                        (N73)? mem[966] :
                        (N44)? mem[1030] :
                        (N46)? mem[1094] :
                        (N48)? mem[1158] :
                        (N50)? mem[1222] :
                        (N52)? mem[1286] :
                        (N54)? mem[1350] :
                        (N56)? mem[1414] :
                        (N58)? mem[1478] :
                        (N60)? mem[1542] :
                        (N62)? mem[1606] :
                        (N64)? mem[1670] :
                        (N66)? mem[1734] :
                        (N68)? mem[1798] :
                        (N70)? mem[1862] :
                        (N72)? mem[1926] :
                        (N74)? mem[1990] : 1'b0;
  assign r0_data_o[5] = (N43)? mem[5] :
                        (N45)? mem[69] :
                        (N47)? mem[133] :
                        (N49)? mem[197] :
                        (N51)? mem[261] :
                        (N53)? mem[325] :
                        (N55)? mem[389] :
                        (N57)? mem[453] :
                        (N59)? mem[517] :
                        (N61)? mem[581] :
                        (N63)? mem[645] :
                        (N65)? mem[709] :
                        (N67)? mem[773] :
                        (N69)? mem[837] :
                        (N71)? mem[901] :
                        (N73)? mem[965] :
                        (N44)? mem[1029] :
                        (N46)? mem[1093] :
                        (N48)? mem[1157] :
                        (N50)? mem[1221] :
                        (N52)? mem[1285] :
                        (N54)? mem[1349] :
                        (N56)? mem[1413] :
                        (N58)? mem[1477] :
                        (N60)? mem[1541] :
                        (N62)? mem[1605] :
                        (N64)? mem[1669] :
                        (N66)? mem[1733] :
                        (N68)? mem[1797] :
                        (N70)? mem[1861] :
                        (N72)? mem[1925] :
                        (N74)? mem[1989] : 1'b0;
  assign r0_data_o[4] = (N43)? mem[4] :
                        (N45)? mem[68] :
                        (N47)? mem[132] :
                        (N49)? mem[196] :
                        (N51)? mem[260] :
                        (N53)? mem[324] :
                        (N55)? mem[388] :
                        (N57)? mem[452] :
                        (N59)? mem[516] :
                        (N61)? mem[580] :
                        (N63)? mem[644] :
                        (N65)? mem[708] :
                        (N67)? mem[772] :
                        (N69)? mem[836] :
                        (N71)? mem[900] :
                        (N73)? mem[964] :
                        (N44)? mem[1028] :
                        (N46)? mem[1092] :
                        (N48)? mem[1156] :
                        (N50)? mem[1220] :
                        (N52)? mem[1284] :
                        (N54)? mem[1348] :
                        (N56)? mem[1412] :
                        (N58)? mem[1476] :
                        (N60)? mem[1540] :
                        (N62)? mem[1604] :
                        (N64)? mem[1668] :
                        (N66)? mem[1732] :
                        (N68)? mem[1796] :
                        (N70)? mem[1860] :
                        (N72)? mem[1924] :
                        (N74)? mem[1988] : 1'b0;
  assign r0_data_o[3] = (N43)? mem[3] :
                        (N45)? mem[67] :
                        (N47)? mem[131] :
                        (N49)? mem[195] :
                        (N51)? mem[259] :
                        (N53)? mem[323] :
                        (N55)? mem[387] :
                        (N57)? mem[451] :
                        (N59)? mem[515] :
                        (N61)? mem[579] :
                        (N63)? mem[643] :
                        (N65)? mem[707] :
                        (N67)? mem[771] :
                        (N69)? mem[835] :
                        (N71)? mem[899] :
                        (N73)? mem[963] :
                        (N44)? mem[1027] :
                        (N46)? mem[1091] :
                        (N48)? mem[1155] :
                        (N50)? mem[1219] :
                        (N52)? mem[1283] :
                        (N54)? mem[1347] :
                        (N56)? mem[1411] :
                        (N58)? mem[1475] :
                        (N60)? mem[1539] :
                        (N62)? mem[1603] :
                        (N64)? mem[1667] :
                        (N66)? mem[1731] :
                        (N68)? mem[1795] :
                        (N70)? mem[1859] :
                        (N72)? mem[1923] :
                        (N74)? mem[1987] : 1'b0;
  assign r0_data_o[2] = (N43)? mem[2] :
                        (N45)? mem[66] :
                        (N47)? mem[130] :
                        (N49)? mem[194] :
                        (N51)? mem[258] :
                        (N53)? mem[322] :
                        (N55)? mem[386] :
                        (N57)? mem[450] :
                        (N59)? mem[514] :
                        (N61)? mem[578] :
                        (N63)? mem[642] :
                        (N65)? mem[706] :
                        (N67)? mem[770] :
                        (N69)? mem[834] :
                        (N71)? mem[898] :
                        (N73)? mem[962] :
                        (N44)? mem[1026] :
                        (N46)? mem[1090] :
                        (N48)? mem[1154] :
                        (N50)? mem[1218] :
                        (N52)? mem[1282] :
                        (N54)? mem[1346] :
                        (N56)? mem[1410] :
                        (N58)? mem[1474] :
                        (N60)? mem[1538] :
                        (N62)? mem[1602] :
                        (N64)? mem[1666] :
                        (N66)? mem[1730] :
                        (N68)? mem[1794] :
                        (N70)? mem[1858] :
                        (N72)? mem[1922] :
                        (N74)? mem[1986] : 1'b0;
  assign r0_data_o[1] = (N43)? mem[1] :
                        (N45)? mem[65] :
                        (N47)? mem[129] :
                        (N49)? mem[193] :
                        (N51)? mem[257] :
                        (N53)? mem[321] :
                        (N55)? mem[385] :
                        (N57)? mem[449] :
                        (N59)? mem[513] :
                        (N61)? mem[577] :
                        (N63)? mem[641] :
                        (N65)? mem[705] :
                        (N67)? mem[769] :
                        (N69)? mem[833] :
                        (N71)? mem[897] :
                        (N73)? mem[961] :
                        (N44)? mem[1025] :
                        (N46)? mem[1089] :
                        (N48)? mem[1153] :
                        (N50)? mem[1217] :
                        (N52)? mem[1281] :
                        (N54)? mem[1345] :
                        (N56)? mem[1409] :
                        (N58)? mem[1473] :
                        (N60)? mem[1537] :
                        (N62)? mem[1601] :
                        (N64)? mem[1665] :
                        (N66)? mem[1729] :
                        (N68)? mem[1793] :
                        (N70)? mem[1857] :
                        (N72)? mem[1921] :
                        (N74)? mem[1985] : 1'b0;
  assign r0_data_o[0] = (N43)? mem[0] :
                        (N45)? mem[64] :
                        (N47)? mem[128] :
                        (N49)? mem[192] :
                        (N51)? mem[256] :
                        (N53)? mem[320] :
                        (N55)? mem[384] :
                        (N57)? mem[448] :
                        (N59)? mem[512] :
                        (N61)? mem[576] :
                        (N63)? mem[640] :
                        (N65)? mem[704] :
                        (N67)? mem[768] :
                        (N69)? mem[832] :
                        (N71)? mem[896] :
                        (N73)? mem[960] :
                        (N44)? mem[1024] :
                        (N46)? mem[1088] :
                        (N48)? mem[1152] :
                        (N50)? mem[1216] :
                        (N52)? mem[1280] :
                        (N54)? mem[1344] :
                        (N56)? mem[1408] :
                        (N58)? mem[1472] :
                        (N60)? mem[1536] :
                        (N62)? mem[1600] :
                        (N64)? mem[1664] :
                        (N66)? mem[1728] :
                        (N68)? mem[1792] :
                        (N70)? mem[1856] :
                        (N72)? mem[1920] :
                        (N74)? mem[1984] : 1'b0;
  assign r1_data_o[63] = (N108)? mem[63] :
                         (N110)? mem[127] :
                         (N112)? mem[191] :
                         (N114)? mem[255] :
                         (N116)? mem[319] :
                         (N118)? mem[383] :
                         (N120)? mem[447] :
                         (N122)? mem[511] :
                         (N124)? mem[575] :
                         (N126)? mem[639] :
                         (N128)? mem[703] :
                         (N130)? mem[767] :
                         (N132)? mem[831] :
                         (N134)? mem[895] :
                         (N136)? mem[959] :
                         (N138)? mem[1023] :
                         (N109)? mem[1087] :
                         (N111)? mem[1151] :
                         (N113)? mem[1215] :
                         (N115)? mem[1279] :
                         (N117)? mem[1343] :
                         (N119)? mem[1407] :
                         (N121)? mem[1471] :
                         (N123)? mem[1535] :
                         (N125)? mem[1599] :
                         (N127)? mem[1663] :
                         (N129)? mem[1727] :
                         (N131)? mem[1791] :
                         (N133)? mem[1855] :
                         (N135)? mem[1919] :
                         (N137)? mem[1983] :
                         (N139)? mem[2047] : 1'b0;
  assign r1_data_o[62] = (N108)? mem[62] :
                         (N110)? mem[126] :
                         (N112)? mem[190] :
                         (N114)? mem[254] :
                         (N116)? mem[318] :
                         (N118)? mem[382] :
                         (N120)? mem[446] :
                         (N122)? mem[510] :
                         (N124)? mem[574] :
                         (N126)? mem[638] :
                         (N128)? mem[702] :
                         (N130)? mem[766] :
                         (N132)? mem[830] :
                         (N134)? mem[894] :
                         (N136)? mem[958] :
                         (N138)? mem[1022] :
                         (N109)? mem[1086] :
                         (N111)? mem[1150] :
                         (N113)? mem[1214] :
                         (N115)? mem[1278] :
                         (N117)? mem[1342] :
                         (N119)? mem[1406] :
                         (N121)? mem[1470] :
                         (N123)? mem[1534] :
                         (N125)? mem[1598] :
                         (N127)? mem[1662] :
                         (N129)? mem[1726] :
                         (N131)? mem[1790] :
                         (N133)? mem[1854] :
                         (N135)? mem[1918] :
                         (N137)? mem[1982] :
                         (N139)? mem[2046] : 1'b0;
  assign r1_data_o[61] = (N108)? mem[61] :
                         (N110)? mem[125] :
                         (N112)? mem[189] :
                         (N114)? mem[253] :
                         (N116)? mem[317] :
                         (N118)? mem[381] :
                         (N120)? mem[445] :
                         (N122)? mem[509] :
                         (N124)? mem[573] :
                         (N126)? mem[637] :
                         (N128)? mem[701] :
                         (N130)? mem[765] :
                         (N132)? mem[829] :
                         (N134)? mem[893] :
                         (N136)? mem[957] :
                         (N138)? mem[1021] :
                         (N109)? mem[1085] :
                         (N111)? mem[1149] :
                         (N113)? mem[1213] :
                         (N115)? mem[1277] :
                         (N117)? mem[1341] :
                         (N119)? mem[1405] :
                         (N121)? mem[1469] :
                         (N123)? mem[1533] :
                         (N125)? mem[1597] :
                         (N127)? mem[1661] :
                         (N129)? mem[1725] :
                         (N131)? mem[1789] :
                         (N133)? mem[1853] :
                         (N135)? mem[1917] :
                         (N137)? mem[1981] :
                         (N139)? mem[2045] : 1'b0;
  assign r1_data_o[60] = (N108)? mem[60] :
                         (N110)? mem[124] :
                         (N112)? mem[188] :
                         (N114)? mem[252] :
                         (N116)? mem[316] :
                         (N118)? mem[380] :
                         (N120)? mem[444] :
                         (N122)? mem[508] :
                         (N124)? mem[572] :
                         (N126)? mem[636] :
                         (N128)? mem[700] :
                         (N130)? mem[764] :
                         (N132)? mem[828] :
                         (N134)? mem[892] :
                         (N136)? mem[956] :
                         (N138)? mem[1020] :
                         (N109)? mem[1084] :
                         (N111)? mem[1148] :
                         (N113)? mem[1212] :
                         (N115)? mem[1276] :
                         (N117)? mem[1340] :
                         (N119)? mem[1404] :
                         (N121)? mem[1468] :
                         (N123)? mem[1532] :
                         (N125)? mem[1596] :
                         (N127)? mem[1660] :
                         (N129)? mem[1724] :
                         (N131)? mem[1788] :
                         (N133)? mem[1852] :
                         (N135)? mem[1916] :
                         (N137)? mem[1980] :
                         (N139)? mem[2044] : 1'b0;
  assign r1_data_o[59] = (N108)? mem[59] :
                         (N110)? mem[123] :
                         (N112)? mem[187] :
                         (N114)? mem[251] :
                         (N116)? mem[315] :
                         (N118)? mem[379] :
                         (N120)? mem[443] :
                         (N122)? mem[507] :
                         (N124)? mem[571] :
                         (N126)? mem[635] :
                         (N128)? mem[699] :
                         (N130)? mem[763] :
                         (N132)? mem[827] :
                         (N134)? mem[891] :
                         (N136)? mem[955] :
                         (N138)? mem[1019] :
                         (N109)? mem[1083] :
                         (N111)? mem[1147] :
                         (N113)? mem[1211] :
                         (N115)? mem[1275] :
                         (N117)? mem[1339] :
                         (N119)? mem[1403] :
                         (N121)? mem[1467] :
                         (N123)? mem[1531] :
                         (N125)? mem[1595] :
                         (N127)? mem[1659] :
                         (N129)? mem[1723] :
                         (N131)? mem[1787] :
                         (N133)? mem[1851] :
                         (N135)? mem[1915] :
                         (N137)? mem[1979] :
                         (N139)? mem[2043] : 1'b0;
  assign r1_data_o[58] = (N108)? mem[58] :
                         (N110)? mem[122] :
                         (N112)? mem[186] :
                         (N114)? mem[250] :
                         (N116)? mem[314] :
                         (N118)? mem[378] :
                         (N120)? mem[442] :
                         (N122)? mem[506] :
                         (N124)? mem[570] :
                         (N126)? mem[634] :
                         (N128)? mem[698] :
                         (N130)? mem[762] :
                         (N132)? mem[826] :
                         (N134)? mem[890] :
                         (N136)? mem[954] :
                         (N138)? mem[1018] :
                         (N109)? mem[1082] :
                         (N111)? mem[1146] :
                         (N113)? mem[1210] :
                         (N115)? mem[1274] :
                         (N117)? mem[1338] :
                         (N119)? mem[1402] :
                         (N121)? mem[1466] :
                         (N123)? mem[1530] :
                         (N125)? mem[1594] :
                         (N127)? mem[1658] :
                         (N129)? mem[1722] :
                         (N131)? mem[1786] :
                         (N133)? mem[1850] :
                         (N135)? mem[1914] :
                         (N137)? mem[1978] :
                         (N139)? mem[2042] : 1'b0;
  assign r1_data_o[57] = (N108)? mem[57] :
                         (N110)? mem[121] :
                         (N112)? mem[185] :
                         (N114)? mem[249] :
                         (N116)? mem[313] :
                         (N118)? mem[377] :
                         (N120)? mem[441] :
                         (N122)? mem[505] :
                         (N124)? mem[569] :
                         (N126)? mem[633] :
                         (N128)? mem[697] :
                         (N130)? mem[761] :
                         (N132)? mem[825] :
                         (N134)? mem[889] :
                         (N136)? mem[953] :
                         (N138)? mem[1017] :
                         (N109)? mem[1081] :
                         (N111)? mem[1145] :
                         (N113)? mem[1209] :
                         (N115)? mem[1273] :
                         (N117)? mem[1337] :
                         (N119)? mem[1401] :
                         (N121)? mem[1465] :
                         (N123)? mem[1529] :
                         (N125)? mem[1593] :
                         (N127)? mem[1657] :
                         (N129)? mem[1721] :
                         (N131)? mem[1785] :
                         (N133)? mem[1849] :
                         (N135)? mem[1913] :
                         (N137)? mem[1977] :
                         (N139)? mem[2041] : 1'b0;
  assign r1_data_o[56] = (N108)? mem[56] :
                         (N110)? mem[120] :
                         (N112)? mem[184] :
                         (N114)? mem[248] :
                         (N116)? mem[312] :
                         (N118)? mem[376] :
                         (N120)? mem[440] :
                         (N122)? mem[504] :
                         (N124)? mem[568] :
                         (N126)? mem[632] :
                         (N128)? mem[696] :
                         (N130)? mem[760] :
                         (N132)? mem[824] :
                         (N134)? mem[888] :
                         (N136)? mem[952] :
                         (N138)? mem[1016] :
                         (N109)? mem[1080] :
                         (N111)? mem[1144] :
                         (N113)? mem[1208] :
                         (N115)? mem[1272] :
                         (N117)? mem[1336] :
                         (N119)? mem[1400] :
                         (N121)? mem[1464] :
                         (N123)? mem[1528] :
                         (N125)? mem[1592] :
                         (N127)? mem[1656] :
                         (N129)? mem[1720] :
                         (N131)? mem[1784] :
                         (N133)? mem[1848] :
                         (N135)? mem[1912] :
                         (N137)? mem[1976] :
                         (N139)? mem[2040] : 1'b0;
  assign r1_data_o[55] = (N108)? mem[55] :
                         (N110)? mem[119] :
                         (N112)? mem[183] :
                         (N114)? mem[247] :
                         (N116)? mem[311] :
                         (N118)? mem[375] :
                         (N120)? mem[439] :
                         (N122)? mem[503] :
                         (N124)? mem[567] :
                         (N126)? mem[631] :
                         (N128)? mem[695] :
                         (N130)? mem[759] :
                         (N132)? mem[823] :
                         (N134)? mem[887] :
                         (N136)? mem[951] :
                         (N138)? mem[1015] :
                         (N109)? mem[1079] :
                         (N111)? mem[1143] :
                         (N113)? mem[1207] :
                         (N115)? mem[1271] :
                         (N117)? mem[1335] :
                         (N119)? mem[1399] :
                         (N121)? mem[1463] :
                         (N123)? mem[1527] :
                         (N125)? mem[1591] :
                         (N127)? mem[1655] :
                         (N129)? mem[1719] :
                         (N131)? mem[1783] :
                         (N133)? mem[1847] :
                         (N135)? mem[1911] :
                         (N137)? mem[1975] :
                         (N139)? mem[2039] : 1'b0;
  assign r1_data_o[54] = (N108)? mem[54] :
                         (N110)? mem[118] :
                         (N112)? mem[182] :
                         (N114)? mem[246] :
                         (N116)? mem[310] :
                         (N118)? mem[374] :
                         (N120)? mem[438] :
                         (N122)? mem[502] :
                         (N124)? mem[566] :
                         (N126)? mem[630] :
                         (N128)? mem[694] :
                         (N130)? mem[758] :
                         (N132)? mem[822] :
                         (N134)? mem[886] :
                         (N136)? mem[950] :
                         (N138)? mem[1014] :
                         (N109)? mem[1078] :
                         (N111)? mem[1142] :
                         (N113)? mem[1206] :
                         (N115)? mem[1270] :
                         (N117)? mem[1334] :
                         (N119)? mem[1398] :
                         (N121)? mem[1462] :
                         (N123)? mem[1526] :
                         (N125)? mem[1590] :
                         (N127)? mem[1654] :
                         (N129)? mem[1718] :
                         (N131)? mem[1782] :
                         (N133)? mem[1846] :
                         (N135)? mem[1910] :
                         (N137)? mem[1974] :
                         (N139)? mem[2038] : 1'b0;
  assign r1_data_o[53] = (N108)? mem[53] :
                         (N110)? mem[117] :
                         (N112)? mem[181] :
                         (N114)? mem[245] :
                         (N116)? mem[309] :
                         (N118)? mem[373] :
                         (N120)? mem[437] :
                         (N122)? mem[501] :
                         (N124)? mem[565] :
                         (N126)? mem[629] :
                         (N128)? mem[693] :
                         (N130)? mem[757] :
                         (N132)? mem[821] :
                         (N134)? mem[885] :
                         (N136)? mem[949] :
                         (N138)? mem[1013] :
                         (N109)? mem[1077] :
                         (N111)? mem[1141] :
                         (N113)? mem[1205] :
                         (N115)? mem[1269] :
                         (N117)? mem[1333] :
                         (N119)? mem[1397] :
                         (N121)? mem[1461] :
                         (N123)? mem[1525] :
                         (N125)? mem[1589] :
                         (N127)? mem[1653] :
                         (N129)? mem[1717] :
                         (N131)? mem[1781] :
                         (N133)? mem[1845] :
                         (N135)? mem[1909] :
                         (N137)? mem[1973] :
                         (N139)? mem[2037] : 1'b0;
  assign r1_data_o[52] = (N108)? mem[52] :
                         (N110)? mem[116] :
                         (N112)? mem[180] :
                         (N114)? mem[244] :
                         (N116)? mem[308] :
                         (N118)? mem[372] :
                         (N120)? mem[436] :
                         (N122)? mem[500] :
                         (N124)? mem[564] :
                         (N126)? mem[628] :
                         (N128)? mem[692] :
                         (N130)? mem[756] :
                         (N132)? mem[820] :
                         (N134)? mem[884] :
                         (N136)? mem[948] :
                         (N138)? mem[1012] :
                         (N109)? mem[1076] :
                         (N111)? mem[1140] :
                         (N113)? mem[1204] :
                         (N115)? mem[1268] :
                         (N117)? mem[1332] :
                         (N119)? mem[1396] :
                         (N121)? mem[1460] :
                         (N123)? mem[1524] :
                         (N125)? mem[1588] :
                         (N127)? mem[1652] :
                         (N129)? mem[1716] :
                         (N131)? mem[1780] :
                         (N133)? mem[1844] :
                         (N135)? mem[1908] :
                         (N137)? mem[1972] :
                         (N139)? mem[2036] : 1'b0;
  assign r1_data_o[51] = (N108)? mem[51] :
                         (N110)? mem[115] :
                         (N112)? mem[179] :
                         (N114)? mem[243] :
                         (N116)? mem[307] :
                         (N118)? mem[371] :
                         (N120)? mem[435] :
                         (N122)? mem[499] :
                         (N124)? mem[563] :
                         (N126)? mem[627] :
                         (N128)? mem[691] :
                         (N130)? mem[755] :
                         (N132)? mem[819] :
                         (N134)? mem[883] :
                         (N136)? mem[947] :
                         (N138)? mem[1011] :
                         (N109)? mem[1075] :
                         (N111)? mem[1139] :
                         (N113)? mem[1203] :
                         (N115)? mem[1267] :
                         (N117)? mem[1331] :
                         (N119)? mem[1395] :
                         (N121)? mem[1459] :
                         (N123)? mem[1523] :
                         (N125)? mem[1587] :
                         (N127)? mem[1651] :
                         (N129)? mem[1715] :
                         (N131)? mem[1779] :
                         (N133)? mem[1843] :
                         (N135)? mem[1907] :
                         (N137)? mem[1971] :
                         (N139)? mem[2035] : 1'b0;
  assign r1_data_o[50] = (N108)? mem[50] :
                         (N110)? mem[114] :
                         (N112)? mem[178] :
                         (N114)? mem[242] :
                         (N116)? mem[306] :
                         (N118)? mem[370] :
                         (N120)? mem[434] :
                         (N122)? mem[498] :
                         (N124)? mem[562] :
                         (N126)? mem[626] :
                         (N128)? mem[690] :
                         (N130)? mem[754] :
                         (N132)? mem[818] :
                         (N134)? mem[882] :
                         (N136)? mem[946] :
                         (N138)? mem[1010] :
                         (N109)? mem[1074] :
                         (N111)? mem[1138] :
                         (N113)? mem[1202] :
                         (N115)? mem[1266] :
                         (N117)? mem[1330] :
                         (N119)? mem[1394] :
                         (N121)? mem[1458] :
                         (N123)? mem[1522] :
                         (N125)? mem[1586] :
                         (N127)? mem[1650] :
                         (N129)? mem[1714] :
                         (N131)? mem[1778] :
                         (N133)? mem[1842] :
                         (N135)? mem[1906] :
                         (N137)? mem[1970] :
                         (N139)? mem[2034] : 1'b0;
  assign r1_data_o[49] = (N108)? mem[49] :
                         (N110)? mem[113] :
                         (N112)? mem[177] :
                         (N114)? mem[241] :
                         (N116)? mem[305] :
                         (N118)? mem[369] :
                         (N120)? mem[433] :
                         (N122)? mem[497] :
                         (N124)? mem[561] :
                         (N126)? mem[625] :
                         (N128)? mem[689] :
                         (N130)? mem[753] :
                         (N132)? mem[817] :
                         (N134)? mem[881] :
                         (N136)? mem[945] :
                         (N138)? mem[1009] :
                         (N109)? mem[1073] :
                         (N111)? mem[1137] :
                         (N113)? mem[1201] :
                         (N115)? mem[1265] :
                         (N117)? mem[1329] :
                         (N119)? mem[1393] :
                         (N121)? mem[1457] :
                         (N123)? mem[1521] :
                         (N125)? mem[1585] :
                         (N127)? mem[1649] :
                         (N129)? mem[1713] :
                         (N131)? mem[1777] :
                         (N133)? mem[1841] :
                         (N135)? mem[1905] :
                         (N137)? mem[1969] :
                         (N139)? mem[2033] : 1'b0;
  assign r1_data_o[48] = (N108)? mem[48] :
                         (N110)? mem[112] :
                         (N112)? mem[176] :
                         (N114)? mem[240] :
                         (N116)? mem[304] :
                         (N118)? mem[368] :
                         (N120)? mem[432] :
                         (N122)? mem[496] :
                         (N124)? mem[560] :
                         (N126)? mem[624] :
                         (N128)? mem[688] :
                         (N130)? mem[752] :
                         (N132)? mem[816] :
                         (N134)? mem[880] :
                         (N136)? mem[944] :
                         (N138)? mem[1008] :
                         (N109)? mem[1072] :
                         (N111)? mem[1136] :
                         (N113)? mem[1200] :
                         (N115)? mem[1264] :
                         (N117)? mem[1328] :
                         (N119)? mem[1392] :
                         (N121)? mem[1456] :
                         (N123)? mem[1520] :
                         (N125)? mem[1584] :
                         (N127)? mem[1648] :
                         (N129)? mem[1712] :
                         (N131)? mem[1776] :
                         (N133)? mem[1840] :
                         (N135)? mem[1904] :
                         (N137)? mem[1968] :
                         (N139)? mem[2032] : 1'b0;
  assign r1_data_o[47] = (N108)? mem[47] :
                         (N110)? mem[111] :
                         (N112)? mem[175] :
                         (N114)? mem[239] :
                         (N116)? mem[303] :
                         (N118)? mem[367] :
                         (N120)? mem[431] :
                         (N122)? mem[495] :
                         (N124)? mem[559] :
                         (N126)? mem[623] :
                         (N128)? mem[687] :
                         (N130)? mem[751] :
                         (N132)? mem[815] :
                         (N134)? mem[879] :
                         (N136)? mem[943] :
                         (N138)? mem[1007] :
                         (N109)? mem[1071] :
                         (N111)? mem[1135] :
                         (N113)? mem[1199] :
                         (N115)? mem[1263] :
                         (N117)? mem[1327] :
                         (N119)? mem[1391] :
                         (N121)? mem[1455] :
                         (N123)? mem[1519] :
                         (N125)? mem[1583] :
                         (N127)? mem[1647] :
                         (N129)? mem[1711] :
                         (N131)? mem[1775] :
                         (N133)? mem[1839] :
                         (N135)? mem[1903] :
                         (N137)? mem[1967] :
                         (N139)? mem[2031] : 1'b0;
  assign r1_data_o[46] = (N108)? mem[46] :
                         (N110)? mem[110] :
                         (N112)? mem[174] :
                         (N114)? mem[238] :
                         (N116)? mem[302] :
                         (N118)? mem[366] :
                         (N120)? mem[430] :
                         (N122)? mem[494] :
                         (N124)? mem[558] :
                         (N126)? mem[622] :
                         (N128)? mem[686] :
                         (N130)? mem[750] :
                         (N132)? mem[814] :
                         (N134)? mem[878] :
                         (N136)? mem[942] :
                         (N138)? mem[1006] :
                         (N109)? mem[1070] :
                         (N111)? mem[1134] :
                         (N113)? mem[1198] :
                         (N115)? mem[1262] :
                         (N117)? mem[1326] :
                         (N119)? mem[1390] :
                         (N121)? mem[1454] :
                         (N123)? mem[1518] :
                         (N125)? mem[1582] :
                         (N127)? mem[1646] :
                         (N129)? mem[1710] :
                         (N131)? mem[1774] :
                         (N133)? mem[1838] :
                         (N135)? mem[1902] :
                         (N137)? mem[1966] :
                         (N139)? mem[2030] : 1'b0;
  assign r1_data_o[45] = (N108)? mem[45] :
                         (N110)? mem[109] :
                         (N112)? mem[173] :
                         (N114)? mem[237] :
                         (N116)? mem[301] :
                         (N118)? mem[365] :
                         (N120)? mem[429] :
                         (N122)? mem[493] :
                         (N124)? mem[557] :
                         (N126)? mem[621] :
                         (N128)? mem[685] :
                         (N130)? mem[749] :
                         (N132)? mem[813] :
                         (N134)? mem[877] :
                         (N136)? mem[941] :
                         (N138)? mem[1005] :
                         (N109)? mem[1069] :
                         (N111)? mem[1133] :
                         (N113)? mem[1197] :
                         (N115)? mem[1261] :
                         (N117)? mem[1325] :
                         (N119)? mem[1389] :
                         (N121)? mem[1453] :
                         (N123)? mem[1517] :
                         (N125)? mem[1581] :
                         (N127)? mem[1645] :
                         (N129)? mem[1709] :
                         (N131)? mem[1773] :
                         (N133)? mem[1837] :
                         (N135)? mem[1901] :
                         (N137)? mem[1965] :
                         (N139)? mem[2029] : 1'b0;
  assign r1_data_o[44] = (N108)? mem[44] :
                         (N110)? mem[108] :
                         (N112)? mem[172] :
                         (N114)? mem[236] :
                         (N116)? mem[300] :
                         (N118)? mem[364] :
                         (N120)? mem[428] :
                         (N122)? mem[492] :
                         (N124)? mem[556] :
                         (N126)? mem[620] :
                         (N128)? mem[684] :
                         (N130)? mem[748] :
                         (N132)? mem[812] :
                         (N134)? mem[876] :
                         (N136)? mem[940] :
                         (N138)? mem[1004] :
                         (N109)? mem[1068] :
                         (N111)? mem[1132] :
                         (N113)? mem[1196] :
                         (N115)? mem[1260] :
                         (N117)? mem[1324] :
                         (N119)? mem[1388] :
                         (N121)? mem[1452] :
                         (N123)? mem[1516] :
                         (N125)? mem[1580] :
                         (N127)? mem[1644] :
                         (N129)? mem[1708] :
                         (N131)? mem[1772] :
                         (N133)? mem[1836] :
                         (N135)? mem[1900] :
                         (N137)? mem[1964] :
                         (N139)? mem[2028] : 1'b0;
  assign r1_data_o[43] = (N108)? mem[43] :
                         (N110)? mem[107] :
                         (N112)? mem[171] :
                         (N114)? mem[235] :
                         (N116)? mem[299] :
                         (N118)? mem[363] :
                         (N120)? mem[427] :
                         (N122)? mem[491] :
                         (N124)? mem[555] :
                         (N126)? mem[619] :
                         (N128)? mem[683] :
                         (N130)? mem[747] :
                         (N132)? mem[811] :
                         (N134)? mem[875] :
                         (N136)? mem[939] :
                         (N138)? mem[1003] :
                         (N109)? mem[1067] :
                         (N111)? mem[1131] :
                         (N113)? mem[1195] :
                         (N115)? mem[1259] :
                         (N117)? mem[1323] :
                         (N119)? mem[1387] :
                         (N121)? mem[1451] :
                         (N123)? mem[1515] :
                         (N125)? mem[1579] :
                         (N127)? mem[1643] :
                         (N129)? mem[1707] :
                         (N131)? mem[1771] :
                         (N133)? mem[1835] :
                         (N135)? mem[1899] :
                         (N137)? mem[1963] :
                         (N139)? mem[2027] : 1'b0;
  assign r1_data_o[42] = (N108)? mem[42] :
                         (N110)? mem[106] :
                         (N112)? mem[170] :
                         (N114)? mem[234] :
                         (N116)? mem[298] :
                         (N118)? mem[362] :
                         (N120)? mem[426] :
                         (N122)? mem[490] :
                         (N124)? mem[554] :
                         (N126)? mem[618] :
                         (N128)? mem[682] :
                         (N130)? mem[746] :
                         (N132)? mem[810] :
                         (N134)? mem[874] :
                         (N136)? mem[938] :
                         (N138)? mem[1002] :
                         (N109)? mem[1066] :
                         (N111)? mem[1130] :
                         (N113)? mem[1194] :
                         (N115)? mem[1258] :
                         (N117)? mem[1322] :
                         (N119)? mem[1386] :
                         (N121)? mem[1450] :
                         (N123)? mem[1514] :
                         (N125)? mem[1578] :
                         (N127)? mem[1642] :
                         (N129)? mem[1706] :
                         (N131)? mem[1770] :
                         (N133)? mem[1834] :
                         (N135)? mem[1898] :
                         (N137)? mem[1962] :
                         (N139)? mem[2026] : 1'b0;
  assign r1_data_o[41] = (N108)? mem[41] :
                         (N110)? mem[105] :
                         (N112)? mem[169] :
                         (N114)? mem[233] :
                         (N116)? mem[297] :
                         (N118)? mem[361] :
                         (N120)? mem[425] :
                         (N122)? mem[489] :
                         (N124)? mem[553] :
                         (N126)? mem[617] :
                         (N128)? mem[681] :
                         (N130)? mem[745] :
                         (N132)? mem[809] :
                         (N134)? mem[873] :
                         (N136)? mem[937] :
                         (N138)? mem[1001] :
                         (N109)? mem[1065] :
                         (N111)? mem[1129] :
                         (N113)? mem[1193] :
                         (N115)? mem[1257] :
                         (N117)? mem[1321] :
                         (N119)? mem[1385] :
                         (N121)? mem[1449] :
                         (N123)? mem[1513] :
                         (N125)? mem[1577] :
                         (N127)? mem[1641] :
                         (N129)? mem[1705] :
                         (N131)? mem[1769] :
                         (N133)? mem[1833] :
                         (N135)? mem[1897] :
                         (N137)? mem[1961] :
                         (N139)? mem[2025] : 1'b0;
  assign r1_data_o[40] = (N108)? mem[40] :
                         (N110)? mem[104] :
                         (N112)? mem[168] :
                         (N114)? mem[232] :
                         (N116)? mem[296] :
                         (N118)? mem[360] :
                         (N120)? mem[424] :
                         (N122)? mem[488] :
                         (N124)? mem[552] :
                         (N126)? mem[616] :
                         (N128)? mem[680] :
                         (N130)? mem[744] :
                         (N132)? mem[808] :
                         (N134)? mem[872] :
                         (N136)? mem[936] :
                         (N138)? mem[1000] :
                         (N109)? mem[1064] :
                         (N111)? mem[1128] :
                         (N113)? mem[1192] :
                         (N115)? mem[1256] :
                         (N117)? mem[1320] :
                         (N119)? mem[1384] :
                         (N121)? mem[1448] :
                         (N123)? mem[1512] :
                         (N125)? mem[1576] :
                         (N127)? mem[1640] :
                         (N129)? mem[1704] :
                         (N131)? mem[1768] :
                         (N133)? mem[1832] :
                         (N135)? mem[1896] :
                         (N137)? mem[1960] :
                         (N139)? mem[2024] : 1'b0;
  assign r1_data_o[39] = (N108)? mem[39] :
                         (N110)? mem[103] :
                         (N112)? mem[167] :
                         (N114)? mem[231] :
                         (N116)? mem[295] :
                         (N118)? mem[359] :
                         (N120)? mem[423] :
                         (N122)? mem[487] :
                         (N124)? mem[551] :
                         (N126)? mem[615] :
                         (N128)? mem[679] :
                         (N130)? mem[743] :
                         (N132)? mem[807] :
                         (N134)? mem[871] :
                         (N136)? mem[935] :
                         (N138)? mem[999] :
                         (N109)? mem[1063] :
                         (N111)? mem[1127] :
                         (N113)? mem[1191] :
                         (N115)? mem[1255] :
                         (N117)? mem[1319] :
                         (N119)? mem[1383] :
                         (N121)? mem[1447] :
                         (N123)? mem[1511] :
                         (N125)? mem[1575] :
                         (N127)? mem[1639] :
                         (N129)? mem[1703] :
                         (N131)? mem[1767] :
                         (N133)? mem[1831] :
                         (N135)? mem[1895] :
                         (N137)? mem[1959] :
                         (N139)? mem[2023] : 1'b0;
  assign r1_data_o[38] = (N108)? mem[38] :
                         (N110)? mem[102] :
                         (N112)? mem[166] :
                         (N114)? mem[230] :
                         (N116)? mem[294] :
                         (N118)? mem[358] :
                         (N120)? mem[422] :
                         (N122)? mem[486] :
                         (N124)? mem[550] :
                         (N126)? mem[614] :
                         (N128)? mem[678] :
                         (N130)? mem[742] :
                         (N132)? mem[806] :
                         (N134)? mem[870] :
                         (N136)? mem[934] :
                         (N138)? mem[998] :
                         (N109)? mem[1062] :
                         (N111)? mem[1126] :
                         (N113)? mem[1190] :
                         (N115)? mem[1254] :
                         (N117)? mem[1318] :
                         (N119)? mem[1382] :
                         (N121)? mem[1446] :
                         (N123)? mem[1510] :
                         (N125)? mem[1574] :
                         (N127)? mem[1638] :
                         (N129)? mem[1702] :
                         (N131)? mem[1766] :
                         (N133)? mem[1830] :
                         (N135)? mem[1894] :
                         (N137)? mem[1958] :
                         (N139)? mem[2022] : 1'b0;
  assign r1_data_o[37] = (N108)? mem[37] :
                         (N110)? mem[101] :
                         (N112)? mem[165] :
                         (N114)? mem[229] :
                         (N116)? mem[293] :
                         (N118)? mem[357] :
                         (N120)? mem[421] :
                         (N122)? mem[485] :
                         (N124)? mem[549] :
                         (N126)? mem[613] :
                         (N128)? mem[677] :
                         (N130)? mem[741] :
                         (N132)? mem[805] :
                         (N134)? mem[869] :
                         (N136)? mem[933] :
                         (N138)? mem[997] :
                         (N109)? mem[1061] :
                         (N111)? mem[1125] :
                         (N113)? mem[1189] :
                         (N115)? mem[1253] :
                         (N117)? mem[1317] :
                         (N119)? mem[1381] :
                         (N121)? mem[1445] :
                         (N123)? mem[1509] :
                         (N125)? mem[1573] :
                         (N127)? mem[1637] :
                         (N129)? mem[1701] :
                         (N131)? mem[1765] :
                         (N133)? mem[1829] :
                         (N135)? mem[1893] :
                         (N137)? mem[1957] :
                         (N139)? mem[2021] : 1'b0;
  assign r1_data_o[36] = (N108)? mem[36] :
                         (N110)? mem[100] :
                         (N112)? mem[164] :
                         (N114)? mem[228] :
                         (N116)? mem[292] :
                         (N118)? mem[356] :
                         (N120)? mem[420] :
                         (N122)? mem[484] :
                         (N124)? mem[548] :
                         (N126)? mem[612] :
                         (N128)? mem[676] :
                         (N130)? mem[740] :
                         (N132)? mem[804] :
                         (N134)? mem[868] :
                         (N136)? mem[932] :
                         (N138)? mem[996] :
                         (N109)? mem[1060] :
                         (N111)? mem[1124] :
                         (N113)? mem[1188] :
                         (N115)? mem[1252] :
                         (N117)? mem[1316] :
                         (N119)? mem[1380] :
                         (N121)? mem[1444] :
                         (N123)? mem[1508] :
                         (N125)? mem[1572] :
                         (N127)? mem[1636] :
                         (N129)? mem[1700] :
                         (N131)? mem[1764] :
                         (N133)? mem[1828] :
                         (N135)? mem[1892] :
                         (N137)? mem[1956] :
                         (N139)? mem[2020] : 1'b0;
  assign r1_data_o[35] = (N108)? mem[35] :
                         (N110)? mem[99] :
                         (N112)? mem[163] :
                         (N114)? mem[227] :
                         (N116)? mem[291] :
                         (N118)? mem[355] :
                         (N120)? mem[419] :
                         (N122)? mem[483] :
                         (N124)? mem[547] :
                         (N126)? mem[611] :
                         (N128)? mem[675] :
                         (N130)? mem[739] :
                         (N132)? mem[803] :
                         (N134)? mem[867] :
                         (N136)? mem[931] :
                         (N138)? mem[995] :
                         (N109)? mem[1059] :
                         (N111)? mem[1123] :
                         (N113)? mem[1187] :
                         (N115)? mem[1251] :
                         (N117)? mem[1315] :
                         (N119)? mem[1379] :
                         (N121)? mem[1443] :
                         (N123)? mem[1507] :
                         (N125)? mem[1571] :
                         (N127)? mem[1635] :
                         (N129)? mem[1699] :
                         (N131)? mem[1763] :
                         (N133)? mem[1827] :
                         (N135)? mem[1891] :
                         (N137)? mem[1955] :
                         (N139)? mem[2019] : 1'b0;
  assign r1_data_o[34] = (N108)? mem[34] :
                         (N110)? mem[98] :
                         (N112)? mem[162] :
                         (N114)? mem[226] :
                         (N116)? mem[290] :
                         (N118)? mem[354] :
                         (N120)? mem[418] :
                         (N122)? mem[482] :
                         (N124)? mem[546] :
                         (N126)? mem[610] :
                         (N128)? mem[674] :
                         (N130)? mem[738] :
                         (N132)? mem[802] :
                         (N134)? mem[866] :
                         (N136)? mem[930] :
                         (N138)? mem[994] :
                         (N109)? mem[1058] :
                         (N111)? mem[1122] :
                         (N113)? mem[1186] :
                         (N115)? mem[1250] :
                         (N117)? mem[1314] :
                         (N119)? mem[1378] :
                         (N121)? mem[1442] :
                         (N123)? mem[1506] :
                         (N125)? mem[1570] :
                         (N127)? mem[1634] :
                         (N129)? mem[1698] :
                         (N131)? mem[1762] :
                         (N133)? mem[1826] :
                         (N135)? mem[1890] :
                         (N137)? mem[1954] :
                         (N139)? mem[2018] : 1'b0;
  assign r1_data_o[33] = (N108)? mem[33] :
                         (N110)? mem[97] :
                         (N112)? mem[161] :
                         (N114)? mem[225] :
                         (N116)? mem[289] :
                         (N118)? mem[353] :
                         (N120)? mem[417] :
                         (N122)? mem[481] :
                         (N124)? mem[545] :
                         (N126)? mem[609] :
                         (N128)? mem[673] :
                         (N130)? mem[737] :
                         (N132)? mem[801] :
                         (N134)? mem[865] :
                         (N136)? mem[929] :
                         (N138)? mem[993] :
                         (N109)? mem[1057] :
                         (N111)? mem[1121] :
                         (N113)? mem[1185] :
                         (N115)? mem[1249] :
                         (N117)? mem[1313] :
                         (N119)? mem[1377] :
                         (N121)? mem[1441] :
                         (N123)? mem[1505] :
                         (N125)? mem[1569] :
                         (N127)? mem[1633] :
                         (N129)? mem[1697] :
                         (N131)? mem[1761] :
                         (N133)? mem[1825] :
                         (N135)? mem[1889] :
                         (N137)? mem[1953] :
                         (N139)? mem[2017] : 1'b0;
  assign r1_data_o[32] = (N108)? mem[32] :
                         (N110)? mem[96] :
                         (N112)? mem[160] :
                         (N114)? mem[224] :
                         (N116)? mem[288] :
                         (N118)? mem[352] :
                         (N120)? mem[416] :
                         (N122)? mem[480] :
                         (N124)? mem[544] :
                         (N126)? mem[608] :
                         (N128)? mem[672] :
                         (N130)? mem[736] :
                         (N132)? mem[800] :
                         (N134)? mem[864] :
                         (N136)? mem[928] :
                         (N138)? mem[992] :
                         (N109)? mem[1056] :
                         (N111)? mem[1120] :
                         (N113)? mem[1184] :
                         (N115)? mem[1248] :
                         (N117)? mem[1312] :
                         (N119)? mem[1376] :
                         (N121)? mem[1440] :
                         (N123)? mem[1504] :
                         (N125)? mem[1568] :
                         (N127)? mem[1632] :
                         (N129)? mem[1696] :
                         (N131)? mem[1760] :
                         (N133)? mem[1824] :
                         (N135)? mem[1888] :
                         (N137)? mem[1952] :
                         (N139)? mem[2016] : 1'b0;
  assign r1_data_o[31] = (N108)? mem[31] :
                         (N110)? mem[95] :
                         (N112)? mem[159] :
                         (N114)? mem[223] :
                         (N116)? mem[287] :
                         (N118)? mem[351] :
                         (N120)? mem[415] :
                         (N122)? mem[479] :
                         (N124)? mem[543] :
                         (N126)? mem[607] :
                         (N128)? mem[671] :
                         (N130)? mem[735] :
                         (N132)? mem[799] :
                         (N134)? mem[863] :
                         (N136)? mem[927] :
                         (N138)? mem[991] :
                         (N109)? mem[1055] :
                         (N111)? mem[1119] :
                         (N113)? mem[1183] :
                         (N115)? mem[1247] :
                         (N117)? mem[1311] :
                         (N119)? mem[1375] :
                         (N121)? mem[1439] :
                         (N123)? mem[1503] :
                         (N125)? mem[1567] :
                         (N127)? mem[1631] :
                         (N129)? mem[1695] :
                         (N131)? mem[1759] :
                         (N133)? mem[1823] :
                         (N135)? mem[1887] :
                         (N137)? mem[1951] :
                         (N139)? mem[2015] : 1'b0;
  assign r1_data_o[30] = (N108)? mem[30] :
                         (N110)? mem[94] :
                         (N112)? mem[158] :
                         (N114)? mem[222] :
                         (N116)? mem[286] :
                         (N118)? mem[350] :
                         (N120)? mem[414] :
                         (N122)? mem[478] :
                         (N124)? mem[542] :
                         (N126)? mem[606] :
                         (N128)? mem[670] :
                         (N130)? mem[734] :
                         (N132)? mem[798] :
                         (N134)? mem[862] :
                         (N136)? mem[926] :
                         (N138)? mem[990] :
                         (N109)? mem[1054] :
                         (N111)? mem[1118] :
                         (N113)? mem[1182] :
                         (N115)? mem[1246] :
                         (N117)? mem[1310] :
                         (N119)? mem[1374] :
                         (N121)? mem[1438] :
                         (N123)? mem[1502] :
                         (N125)? mem[1566] :
                         (N127)? mem[1630] :
                         (N129)? mem[1694] :
                         (N131)? mem[1758] :
                         (N133)? mem[1822] :
                         (N135)? mem[1886] :
                         (N137)? mem[1950] :
                         (N139)? mem[2014] : 1'b0;
  assign r1_data_o[29] = (N108)? mem[29] :
                         (N110)? mem[93] :
                         (N112)? mem[157] :
                         (N114)? mem[221] :
                         (N116)? mem[285] :
                         (N118)? mem[349] :
                         (N120)? mem[413] :
                         (N122)? mem[477] :
                         (N124)? mem[541] :
                         (N126)? mem[605] :
                         (N128)? mem[669] :
                         (N130)? mem[733] :
                         (N132)? mem[797] :
                         (N134)? mem[861] :
                         (N136)? mem[925] :
                         (N138)? mem[989] :
                         (N109)? mem[1053] :
                         (N111)? mem[1117] :
                         (N113)? mem[1181] :
                         (N115)? mem[1245] :
                         (N117)? mem[1309] :
                         (N119)? mem[1373] :
                         (N121)? mem[1437] :
                         (N123)? mem[1501] :
                         (N125)? mem[1565] :
                         (N127)? mem[1629] :
                         (N129)? mem[1693] :
                         (N131)? mem[1757] :
                         (N133)? mem[1821] :
                         (N135)? mem[1885] :
                         (N137)? mem[1949] :
                         (N139)? mem[2013] : 1'b0;
  assign r1_data_o[28] = (N108)? mem[28] :
                         (N110)? mem[92] :
                         (N112)? mem[156] :
                         (N114)? mem[220] :
                         (N116)? mem[284] :
                         (N118)? mem[348] :
                         (N120)? mem[412] :
                         (N122)? mem[476] :
                         (N124)? mem[540] :
                         (N126)? mem[604] :
                         (N128)? mem[668] :
                         (N130)? mem[732] :
                         (N132)? mem[796] :
                         (N134)? mem[860] :
                         (N136)? mem[924] :
                         (N138)? mem[988] :
                         (N109)? mem[1052] :
                         (N111)? mem[1116] :
                         (N113)? mem[1180] :
                         (N115)? mem[1244] :
                         (N117)? mem[1308] :
                         (N119)? mem[1372] :
                         (N121)? mem[1436] :
                         (N123)? mem[1500] :
                         (N125)? mem[1564] :
                         (N127)? mem[1628] :
                         (N129)? mem[1692] :
                         (N131)? mem[1756] :
                         (N133)? mem[1820] :
                         (N135)? mem[1884] :
                         (N137)? mem[1948] :
                         (N139)? mem[2012] : 1'b0;
  assign r1_data_o[27] = (N108)? mem[27] :
                         (N110)? mem[91] :
                         (N112)? mem[155] :
                         (N114)? mem[219] :
                         (N116)? mem[283] :
                         (N118)? mem[347] :
                         (N120)? mem[411] :
                         (N122)? mem[475] :
                         (N124)? mem[539] :
                         (N126)? mem[603] :
                         (N128)? mem[667] :
                         (N130)? mem[731] :
                         (N132)? mem[795] :
                         (N134)? mem[859] :
                         (N136)? mem[923] :
                         (N138)? mem[987] :
                         (N109)? mem[1051] :
                         (N111)? mem[1115] :
                         (N113)? mem[1179] :
                         (N115)? mem[1243] :
                         (N117)? mem[1307] :
                         (N119)? mem[1371] :
                         (N121)? mem[1435] :
                         (N123)? mem[1499] :
                         (N125)? mem[1563] :
                         (N127)? mem[1627] :
                         (N129)? mem[1691] :
                         (N131)? mem[1755] :
                         (N133)? mem[1819] :
                         (N135)? mem[1883] :
                         (N137)? mem[1947] :
                         (N139)? mem[2011] : 1'b0;
  assign r1_data_o[26] = (N108)? mem[26] :
                         (N110)? mem[90] :
                         (N112)? mem[154] :
                         (N114)? mem[218] :
                         (N116)? mem[282] :
                         (N118)? mem[346] :
                         (N120)? mem[410] :
                         (N122)? mem[474] :
                         (N124)? mem[538] :
                         (N126)? mem[602] :
                         (N128)? mem[666] :
                         (N130)? mem[730] :
                         (N132)? mem[794] :
                         (N134)? mem[858] :
                         (N136)? mem[922] :
                         (N138)? mem[986] :
                         (N109)? mem[1050] :
                         (N111)? mem[1114] :
                         (N113)? mem[1178] :
                         (N115)? mem[1242] :
                         (N117)? mem[1306] :
                         (N119)? mem[1370] :
                         (N121)? mem[1434] :
                         (N123)? mem[1498] :
                         (N125)? mem[1562] :
                         (N127)? mem[1626] :
                         (N129)? mem[1690] :
                         (N131)? mem[1754] :
                         (N133)? mem[1818] :
                         (N135)? mem[1882] :
                         (N137)? mem[1946] :
                         (N139)? mem[2010] : 1'b0;
  assign r1_data_o[25] = (N108)? mem[25] :
                         (N110)? mem[89] :
                         (N112)? mem[153] :
                         (N114)? mem[217] :
                         (N116)? mem[281] :
                         (N118)? mem[345] :
                         (N120)? mem[409] :
                         (N122)? mem[473] :
                         (N124)? mem[537] :
                         (N126)? mem[601] :
                         (N128)? mem[665] :
                         (N130)? mem[729] :
                         (N132)? mem[793] :
                         (N134)? mem[857] :
                         (N136)? mem[921] :
                         (N138)? mem[985] :
                         (N109)? mem[1049] :
                         (N111)? mem[1113] :
                         (N113)? mem[1177] :
                         (N115)? mem[1241] :
                         (N117)? mem[1305] :
                         (N119)? mem[1369] :
                         (N121)? mem[1433] :
                         (N123)? mem[1497] :
                         (N125)? mem[1561] :
                         (N127)? mem[1625] :
                         (N129)? mem[1689] :
                         (N131)? mem[1753] :
                         (N133)? mem[1817] :
                         (N135)? mem[1881] :
                         (N137)? mem[1945] :
                         (N139)? mem[2009] : 1'b0;
  assign r1_data_o[24] = (N108)? mem[24] :
                         (N110)? mem[88] :
                         (N112)? mem[152] :
                         (N114)? mem[216] :
                         (N116)? mem[280] :
                         (N118)? mem[344] :
                         (N120)? mem[408] :
                         (N122)? mem[472] :
                         (N124)? mem[536] :
                         (N126)? mem[600] :
                         (N128)? mem[664] :
                         (N130)? mem[728] :
                         (N132)? mem[792] :
                         (N134)? mem[856] :
                         (N136)? mem[920] :
                         (N138)? mem[984] :
                         (N109)? mem[1048] :
                         (N111)? mem[1112] :
                         (N113)? mem[1176] :
                         (N115)? mem[1240] :
                         (N117)? mem[1304] :
                         (N119)? mem[1368] :
                         (N121)? mem[1432] :
                         (N123)? mem[1496] :
                         (N125)? mem[1560] :
                         (N127)? mem[1624] :
                         (N129)? mem[1688] :
                         (N131)? mem[1752] :
                         (N133)? mem[1816] :
                         (N135)? mem[1880] :
                         (N137)? mem[1944] :
                         (N139)? mem[2008] : 1'b0;
  assign r1_data_o[23] = (N108)? mem[23] :
                         (N110)? mem[87] :
                         (N112)? mem[151] :
                         (N114)? mem[215] :
                         (N116)? mem[279] :
                         (N118)? mem[343] :
                         (N120)? mem[407] :
                         (N122)? mem[471] :
                         (N124)? mem[535] :
                         (N126)? mem[599] :
                         (N128)? mem[663] :
                         (N130)? mem[727] :
                         (N132)? mem[791] :
                         (N134)? mem[855] :
                         (N136)? mem[919] :
                         (N138)? mem[983] :
                         (N109)? mem[1047] :
                         (N111)? mem[1111] :
                         (N113)? mem[1175] :
                         (N115)? mem[1239] :
                         (N117)? mem[1303] :
                         (N119)? mem[1367] :
                         (N121)? mem[1431] :
                         (N123)? mem[1495] :
                         (N125)? mem[1559] :
                         (N127)? mem[1623] :
                         (N129)? mem[1687] :
                         (N131)? mem[1751] :
                         (N133)? mem[1815] :
                         (N135)? mem[1879] :
                         (N137)? mem[1943] :
                         (N139)? mem[2007] : 1'b0;
  assign r1_data_o[22] = (N108)? mem[22] :
                         (N110)? mem[86] :
                         (N112)? mem[150] :
                         (N114)? mem[214] :
                         (N116)? mem[278] :
                         (N118)? mem[342] :
                         (N120)? mem[406] :
                         (N122)? mem[470] :
                         (N124)? mem[534] :
                         (N126)? mem[598] :
                         (N128)? mem[662] :
                         (N130)? mem[726] :
                         (N132)? mem[790] :
                         (N134)? mem[854] :
                         (N136)? mem[918] :
                         (N138)? mem[982] :
                         (N109)? mem[1046] :
                         (N111)? mem[1110] :
                         (N113)? mem[1174] :
                         (N115)? mem[1238] :
                         (N117)? mem[1302] :
                         (N119)? mem[1366] :
                         (N121)? mem[1430] :
                         (N123)? mem[1494] :
                         (N125)? mem[1558] :
                         (N127)? mem[1622] :
                         (N129)? mem[1686] :
                         (N131)? mem[1750] :
                         (N133)? mem[1814] :
                         (N135)? mem[1878] :
                         (N137)? mem[1942] :
                         (N139)? mem[2006] : 1'b0;
  assign r1_data_o[21] = (N108)? mem[21] :
                         (N110)? mem[85] :
                         (N112)? mem[149] :
                         (N114)? mem[213] :
                         (N116)? mem[277] :
                         (N118)? mem[341] :
                         (N120)? mem[405] :
                         (N122)? mem[469] :
                         (N124)? mem[533] :
                         (N126)? mem[597] :
                         (N128)? mem[661] :
                         (N130)? mem[725] :
                         (N132)? mem[789] :
                         (N134)? mem[853] :
                         (N136)? mem[917] :
                         (N138)? mem[981] :
                         (N109)? mem[1045] :
                         (N111)? mem[1109] :
                         (N113)? mem[1173] :
                         (N115)? mem[1237] :
                         (N117)? mem[1301] :
                         (N119)? mem[1365] :
                         (N121)? mem[1429] :
                         (N123)? mem[1493] :
                         (N125)? mem[1557] :
                         (N127)? mem[1621] :
                         (N129)? mem[1685] :
                         (N131)? mem[1749] :
                         (N133)? mem[1813] :
                         (N135)? mem[1877] :
                         (N137)? mem[1941] :
                         (N139)? mem[2005] : 1'b0;
  assign r1_data_o[20] = (N108)? mem[20] :
                         (N110)? mem[84] :
                         (N112)? mem[148] :
                         (N114)? mem[212] :
                         (N116)? mem[276] :
                         (N118)? mem[340] :
                         (N120)? mem[404] :
                         (N122)? mem[468] :
                         (N124)? mem[532] :
                         (N126)? mem[596] :
                         (N128)? mem[660] :
                         (N130)? mem[724] :
                         (N132)? mem[788] :
                         (N134)? mem[852] :
                         (N136)? mem[916] :
                         (N138)? mem[980] :
                         (N109)? mem[1044] :
                         (N111)? mem[1108] :
                         (N113)? mem[1172] :
                         (N115)? mem[1236] :
                         (N117)? mem[1300] :
                         (N119)? mem[1364] :
                         (N121)? mem[1428] :
                         (N123)? mem[1492] :
                         (N125)? mem[1556] :
                         (N127)? mem[1620] :
                         (N129)? mem[1684] :
                         (N131)? mem[1748] :
                         (N133)? mem[1812] :
                         (N135)? mem[1876] :
                         (N137)? mem[1940] :
                         (N139)? mem[2004] : 1'b0;
  assign r1_data_o[19] = (N108)? mem[19] :
                         (N110)? mem[83] :
                         (N112)? mem[147] :
                         (N114)? mem[211] :
                         (N116)? mem[275] :
                         (N118)? mem[339] :
                         (N120)? mem[403] :
                         (N122)? mem[467] :
                         (N124)? mem[531] :
                         (N126)? mem[595] :
                         (N128)? mem[659] :
                         (N130)? mem[723] :
                         (N132)? mem[787] :
                         (N134)? mem[851] :
                         (N136)? mem[915] :
                         (N138)? mem[979] :
                         (N109)? mem[1043] :
                         (N111)? mem[1107] :
                         (N113)? mem[1171] :
                         (N115)? mem[1235] :
                         (N117)? mem[1299] :
                         (N119)? mem[1363] :
                         (N121)? mem[1427] :
                         (N123)? mem[1491] :
                         (N125)? mem[1555] :
                         (N127)? mem[1619] :
                         (N129)? mem[1683] :
                         (N131)? mem[1747] :
                         (N133)? mem[1811] :
                         (N135)? mem[1875] :
                         (N137)? mem[1939] :
                         (N139)? mem[2003] : 1'b0;
  assign r1_data_o[18] = (N108)? mem[18] :
                         (N110)? mem[82] :
                         (N112)? mem[146] :
                         (N114)? mem[210] :
                         (N116)? mem[274] :
                         (N118)? mem[338] :
                         (N120)? mem[402] :
                         (N122)? mem[466] :
                         (N124)? mem[530] :
                         (N126)? mem[594] :
                         (N128)? mem[658] :
                         (N130)? mem[722] :
                         (N132)? mem[786] :
                         (N134)? mem[850] :
                         (N136)? mem[914] :
                         (N138)? mem[978] :
                         (N109)? mem[1042] :
                         (N111)? mem[1106] :
                         (N113)? mem[1170] :
                         (N115)? mem[1234] :
                         (N117)? mem[1298] :
                         (N119)? mem[1362] :
                         (N121)? mem[1426] :
                         (N123)? mem[1490] :
                         (N125)? mem[1554] :
                         (N127)? mem[1618] :
                         (N129)? mem[1682] :
                         (N131)? mem[1746] :
                         (N133)? mem[1810] :
                         (N135)? mem[1874] :
                         (N137)? mem[1938] :
                         (N139)? mem[2002] : 1'b0;
  assign r1_data_o[17] = (N108)? mem[17] :
                         (N110)? mem[81] :
                         (N112)? mem[145] :
                         (N114)? mem[209] :
                         (N116)? mem[273] :
                         (N118)? mem[337] :
                         (N120)? mem[401] :
                         (N122)? mem[465] :
                         (N124)? mem[529] :
                         (N126)? mem[593] :
                         (N128)? mem[657] :
                         (N130)? mem[721] :
                         (N132)? mem[785] :
                         (N134)? mem[849] :
                         (N136)? mem[913] :
                         (N138)? mem[977] :
                         (N109)? mem[1041] :
                         (N111)? mem[1105] :
                         (N113)? mem[1169] :
                         (N115)? mem[1233] :
                         (N117)? mem[1297] :
                         (N119)? mem[1361] :
                         (N121)? mem[1425] :
                         (N123)? mem[1489] :
                         (N125)? mem[1553] :
                         (N127)? mem[1617] :
                         (N129)? mem[1681] :
                         (N131)? mem[1745] :
                         (N133)? mem[1809] :
                         (N135)? mem[1873] :
                         (N137)? mem[1937] :
                         (N139)? mem[2001] : 1'b0;
  assign r1_data_o[16] = (N108)? mem[16] :
                         (N110)? mem[80] :
                         (N112)? mem[144] :
                         (N114)? mem[208] :
                         (N116)? mem[272] :
                         (N118)? mem[336] :
                         (N120)? mem[400] :
                         (N122)? mem[464] :
                         (N124)? mem[528] :
                         (N126)? mem[592] :
                         (N128)? mem[656] :
                         (N130)? mem[720] :
                         (N132)? mem[784] :
                         (N134)? mem[848] :
                         (N136)? mem[912] :
                         (N138)? mem[976] :
                         (N109)? mem[1040] :
                         (N111)? mem[1104] :
                         (N113)? mem[1168] :
                         (N115)? mem[1232] :
                         (N117)? mem[1296] :
                         (N119)? mem[1360] :
                         (N121)? mem[1424] :
                         (N123)? mem[1488] :
                         (N125)? mem[1552] :
                         (N127)? mem[1616] :
                         (N129)? mem[1680] :
                         (N131)? mem[1744] :
                         (N133)? mem[1808] :
                         (N135)? mem[1872] :
                         (N137)? mem[1936] :
                         (N139)? mem[2000] : 1'b0;
  assign r1_data_o[15] = (N108)? mem[15] :
                         (N110)? mem[79] :
                         (N112)? mem[143] :
                         (N114)? mem[207] :
                         (N116)? mem[271] :
                         (N118)? mem[335] :
                         (N120)? mem[399] :
                         (N122)? mem[463] :
                         (N124)? mem[527] :
                         (N126)? mem[591] :
                         (N128)? mem[655] :
                         (N130)? mem[719] :
                         (N132)? mem[783] :
                         (N134)? mem[847] :
                         (N136)? mem[911] :
                         (N138)? mem[975] :
                         (N109)? mem[1039] :
                         (N111)? mem[1103] :
                         (N113)? mem[1167] :
                         (N115)? mem[1231] :
                         (N117)? mem[1295] :
                         (N119)? mem[1359] :
                         (N121)? mem[1423] :
                         (N123)? mem[1487] :
                         (N125)? mem[1551] :
                         (N127)? mem[1615] :
                         (N129)? mem[1679] :
                         (N131)? mem[1743] :
                         (N133)? mem[1807] :
                         (N135)? mem[1871] :
                         (N137)? mem[1935] :
                         (N139)? mem[1999] : 1'b0;
  assign r1_data_o[14] = (N108)? mem[14] :
                         (N110)? mem[78] :
                         (N112)? mem[142] :
                         (N114)? mem[206] :
                         (N116)? mem[270] :
                         (N118)? mem[334] :
                         (N120)? mem[398] :
                         (N122)? mem[462] :
                         (N124)? mem[526] :
                         (N126)? mem[590] :
                         (N128)? mem[654] :
                         (N130)? mem[718] :
                         (N132)? mem[782] :
                         (N134)? mem[846] :
                         (N136)? mem[910] :
                         (N138)? mem[974] :
                         (N109)? mem[1038] :
                         (N111)? mem[1102] :
                         (N113)? mem[1166] :
                         (N115)? mem[1230] :
                         (N117)? mem[1294] :
                         (N119)? mem[1358] :
                         (N121)? mem[1422] :
                         (N123)? mem[1486] :
                         (N125)? mem[1550] :
                         (N127)? mem[1614] :
                         (N129)? mem[1678] :
                         (N131)? mem[1742] :
                         (N133)? mem[1806] :
                         (N135)? mem[1870] :
                         (N137)? mem[1934] :
                         (N139)? mem[1998] : 1'b0;
  assign r1_data_o[13] = (N108)? mem[13] :
                         (N110)? mem[77] :
                         (N112)? mem[141] :
                         (N114)? mem[205] :
                         (N116)? mem[269] :
                         (N118)? mem[333] :
                         (N120)? mem[397] :
                         (N122)? mem[461] :
                         (N124)? mem[525] :
                         (N126)? mem[589] :
                         (N128)? mem[653] :
                         (N130)? mem[717] :
                         (N132)? mem[781] :
                         (N134)? mem[845] :
                         (N136)? mem[909] :
                         (N138)? mem[973] :
                         (N109)? mem[1037] :
                         (N111)? mem[1101] :
                         (N113)? mem[1165] :
                         (N115)? mem[1229] :
                         (N117)? mem[1293] :
                         (N119)? mem[1357] :
                         (N121)? mem[1421] :
                         (N123)? mem[1485] :
                         (N125)? mem[1549] :
                         (N127)? mem[1613] :
                         (N129)? mem[1677] :
                         (N131)? mem[1741] :
                         (N133)? mem[1805] :
                         (N135)? mem[1869] :
                         (N137)? mem[1933] :
                         (N139)? mem[1997] : 1'b0;
  assign r1_data_o[12] = (N108)? mem[12] :
                         (N110)? mem[76] :
                         (N112)? mem[140] :
                         (N114)? mem[204] :
                         (N116)? mem[268] :
                         (N118)? mem[332] :
                         (N120)? mem[396] :
                         (N122)? mem[460] :
                         (N124)? mem[524] :
                         (N126)? mem[588] :
                         (N128)? mem[652] :
                         (N130)? mem[716] :
                         (N132)? mem[780] :
                         (N134)? mem[844] :
                         (N136)? mem[908] :
                         (N138)? mem[972] :
                         (N109)? mem[1036] :
                         (N111)? mem[1100] :
                         (N113)? mem[1164] :
                         (N115)? mem[1228] :
                         (N117)? mem[1292] :
                         (N119)? mem[1356] :
                         (N121)? mem[1420] :
                         (N123)? mem[1484] :
                         (N125)? mem[1548] :
                         (N127)? mem[1612] :
                         (N129)? mem[1676] :
                         (N131)? mem[1740] :
                         (N133)? mem[1804] :
                         (N135)? mem[1868] :
                         (N137)? mem[1932] :
                         (N139)? mem[1996] : 1'b0;
  assign r1_data_o[11] = (N108)? mem[11] :
                         (N110)? mem[75] :
                         (N112)? mem[139] :
                         (N114)? mem[203] :
                         (N116)? mem[267] :
                         (N118)? mem[331] :
                         (N120)? mem[395] :
                         (N122)? mem[459] :
                         (N124)? mem[523] :
                         (N126)? mem[587] :
                         (N128)? mem[651] :
                         (N130)? mem[715] :
                         (N132)? mem[779] :
                         (N134)? mem[843] :
                         (N136)? mem[907] :
                         (N138)? mem[971] :
                         (N109)? mem[1035] :
                         (N111)? mem[1099] :
                         (N113)? mem[1163] :
                         (N115)? mem[1227] :
                         (N117)? mem[1291] :
                         (N119)? mem[1355] :
                         (N121)? mem[1419] :
                         (N123)? mem[1483] :
                         (N125)? mem[1547] :
                         (N127)? mem[1611] :
                         (N129)? mem[1675] :
                         (N131)? mem[1739] :
                         (N133)? mem[1803] :
                         (N135)? mem[1867] :
                         (N137)? mem[1931] :
                         (N139)? mem[1995] : 1'b0;
  assign r1_data_o[10] = (N108)? mem[10] :
                         (N110)? mem[74] :
                         (N112)? mem[138] :
                         (N114)? mem[202] :
                         (N116)? mem[266] :
                         (N118)? mem[330] :
                         (N120)? mem[394] :
                         (N122)? mem[458] :
                         (N124)? mem[522] :
                         (N126)? mem[586] :
                         (N128)? mem[650] :
                         (N130)? mem[714] :
                         (N132)? mem[778] :
                         (N134)? mem[842] :
                         (N136)? mem[906] :
                         (N138)? mem[970] :
                         (N109)? mem[1034] :
                         (N111)? mem[1098] :
                         (N113)? mem[1162] :
                         (N115)? mem[1226] :
                         (N117)? mem[1290] :
                         (N119)? mem[1354] :
                         (N121)? mem[1418] :
                         (N123)? mem[1482] :
                         (N125)? mem[1546] :
                         (N127)? mem[1610] :
                         (N129)? mem[1674] :
                         (N131)? mem[1738] :
                         (N133)? mem[1802] :
                         (N135)? mem[1866] :
                         (N137)? mem[1930] :
                         (N139)? mem[1994] : 1'b0;
  assign r1_data_o[9] = (N108)? mem[9] :
                        (N110)? mem[73] :
                        (N112)? mem[137] :
                        (N114)? mem[201] :
                        (N116)? mem[265] :
                        (N118)? mem[329] :
                        (N120)? mem[393] :
                        (N122)? mem[457] :
                        (N124)? mem[521] :
                        (N126)? mem[585] :
                        (N128)? mem[649] :
                        (N130)? mem[713] :
                        (N132)? mem[777] :
                        (N134)? mem[841] :
                        (N136)? mem[905] :
                        (N138)? mem[969] :
                        (N109)? mem[1033] :
                        (N111)? mem[1097] :
                        (N113)? mem[1161] :
                        (N115)? mem[1225] :
                        (N117)? mem[1289] :
                        (N119)? mem[1353] :
                        (N121)? mem[1417] :
                        (N123)? mem[1481] :
                        (N125)? mem[1545] :
                        (N127)? mem[1609] :
                        (N129)? mem[1673] :
                        (N131)? mem[1737] :
                        (N133)? mem[1801] :
                        (N135)? mem[1865] :
                        (N137)? mem[1929] :
                        (N139)? mem[1993] : 1'b0;
  assign r1_data_o[8] = (N108)? mem[8] :
                        (N110)? mem[72] :
                        (N112)? mem[136] :
                        (N114)? mem[200] :
                        (N116)? mem[264] :
                        (N118)? mem[328] :
                        (N120)? mem[392] :
                        (N122)? mem[456] :
                        (N124)? mem[520] :
                        (N126)? mem[584] :
                        (N128)? mem[648] :
                        (N130)? mem[712] :
                        (N132)? mem[776] :
                        (N134)? mem[840] :
                        (N136)? mem[904] :
                        (N138)? mem[968] :
                        (N109)? mem[1032] :
                        (N111)? mem[1096] :
                        (N113)? mem[1160] :
                        (N115)? mem[1224] :
                        (N117)? mem[1288] :
                        (N119)? mem[1352] :
                        (N121)? mem[1416] :
                        (N123)? mem[1480] :
                        (N125)? mem[1544] :
                        (N127)? mem[1608] :
                        (N129)? mem[1672] :
                        (N131)? mem[1736] :
                        (N133)? mem[1800] :
                        (N135)? mem[1864] :
                        (N137)? mem[1928] :
                        (N139)? mem[1992] : 1'b0;
  assign r1_data_o[7] = (N108)? mem[7] :
                        (N110)? mem[71] :
                        (N112)? mem[135] :
                        (N114)? mem[199] :
                        (N116)? mem[263] :
                        (N118)? mem[327] :
                        (N120)? mem[391] :
                        (N122)? mem[455] :
                        (N124)? mem[519] :
                        (N126)? mem[583] :
                        (N128)? mem[647] :
                        (N130)? mem[711] :
                        (N132)? mem[775] :
                        (N134)? mem[839] :
                        (N136)? mem[903] :
                        (N138)? mem[967] :
                        (N109)? mem[1031] :
                        (N111)? mem[1095] :
                        (N113)? mem[1159] :
                        (N115)? mem[1223] :
                        (N117)? mem[1287] :
                        (N119)? mem[1351] :
                        (N121)? mem[1415] :
                        (N123)? mem[1479] :
                        (N125)? mem[1543] :
                        (N127)? mem[1607] :
                        (N129)? mem[1671] :
                        (N131)? mem[1735] :
                        (N133)? mem[1799] :
                        (N135)? mem[1863] :
                        (N137)? mem[1927] :
                        (N139)? mem[1991] : 1'b0;
  assign r1_data_o[6] = (N108)? mem[6] :
                        (N110)? mem[70] :
                        (N112)? mem[134] :
                        (N114)? mem[198] :
                        (N116)? mem[262] :
                        (N118)? mem[326] :
                        (N120)? mem[390] :
                        (N122)? mem[454] :
                        (N124)? mem[518] :
                        (N126)? mem[582] :
                        (N128)? mem[646] :
                        (N130)? mem[710] :
                        (N132)? mem[774] :
                        (N134)? mem[838] :
                        (N136)? mem[902] :
                        (N138)? mem[966] :
                        (N109)? mem[1030] :
                        (N111)? mem[1094] :
                        (N113)? mem[1158] :
                        (N115)? mem[1222] :
                        (N117)? mem[1286] :
                        (N119)? mem[1350] :
                        (N121)? mem[1414] :
                        (N123)? mem[1478] :
                        (N125)? mem[1542] :
                        (N127)? mem[1606] :
                        (N129)? mem[1670] :
                        (N131)? mem[1734] :
                        (N133)? mem[1798] :
                        (N135)? mem[1862] :
                        (N137)? mem[1926] :
                        (N139)? mem[1990] : 1'b0;
  assign r1_data_o[5] = (N108)? mem[5] :
                        (N110)? mem[69] :
                        (N112)? mem[133] :
                        (N114)? mem[197] :
                        (N116)? mem[261] :
                        (N118)? mem[325] :
                        (N120)? mem[389] :
                        (N122)? mem[453] :
                        (N124)? mem[517] :
                        (N126)? mem[581] :
                        (N128)? mem[645] :
                        (N130)? mem[709] :
                        (N132)? mem[773] :
                        (N134)? mem[837] :
                        (N136)? mem[901] :
                        (N138)? mem[965] :
                        (N109)? mem[1029] :
                        (N111)? mem[1093] :
                        (N113)? mem[1157] :
                        (N115)? mem[1221] :
                        (N117)? mem[1285] :
                        (N119)? mem[1349] :
                        (N121)? mem[1413] :
                        (N123)? mem[1477] :
                        (N125)? mem[1541] :
                        (N127)? mem[1605] :
                        (N129)? mem[1669] :
                        (N131)? mem[1733] :
                        (N133)? mem[1797] :
                        (N135)? mem[1861] :
                        (N137)? mem[1925] :
                        (N139)? mem[1989] : 1'b0;
  assign r1_data_o[4] = (N108)? mem[4] :
                        (N110)? mem[68] :
                        (N112)? mem[132] :
                        (N114)? mem[196] :
                        (N116)? mem[260] :
                        (N118)? mem[324] :
                        (N120)? mem[388] :
                        (N122)? mem[452] :
                        (N124)? mem[516] :
                        (N126)? mem[580] :
                        (N128)? mem[644] :
                        (N130)? mem[708] :
                        (N132)? mem[772] :
                        (N134)? mem[836] :
                        (N136)? mem[900] :
                        (N138)? mem[964] :
                        (N109)? mem[1028] :
                        (N111)? mem[1092] :
                        (N113)? mem[1156] :
                        (N115)? mem[1220] :
                        (N117)? mem[1284] :
                        (N119)? mem[1348] :
                        (N121)? mem[1412] :
                        (N123)? mem[1476] :
                        (N125)? mem[1540] :
                        (N127)? mem[1604] :
                        (N129)? mem[1668] :
                        (N131)? mem[1732] :
                        (N133)? mem[1796] :
                        (N135)? mem[1860] :
                        (N137)? mem[1924] :
                        (N139)? mem[1988] : 1'b0;
  assign r1_data_o[3] = (N108)? mem[3] :
                        (N110)? mem[67] :
                        (N112)? mem[131] :
                        (N114)? mem[195] :
                        (N116)? mem[259] :
                        (N118)? mem[323] :
                        (N120)? mem[387] :
                        (N122)? mem[451] :
                        (N124)? mem[515] :
                        (N126)? mem[579] :
                        (N128)? mem[643] :
                        (N130)? mem[707] :
                        (N132)? mem[771] :
                        (N134)? mem[835] :
                        (N136)? mem[899] :
                        (N138)? mem[963] :
                        (N109)? mem[1027] :
                        (N111)? mem[1091] :
                        (N113)? mem[1155] :
                        (N115)? mem[1219] :
                        (N117)? mem[1283] :
                        (N119)? mem[1347] :
                        (N121)? mem[1411] :
                        (N123)? mem[1475] :
                        (N125)? mem[1539] :
                        (N127)? mem[1603] :
                        (N129)? mem[1667] :
                        (N131)? mem[1731] :
                        (N133)? mem[1795] :
                        (N135)? mem[1859] :
                        (N137)? mem[1923] :
                        (N139)? mem[1987] : 1'b0;
  assign r1_data_o[2] = (N108)? mem[2] :
                        (N110)? mem[66] :
                        (N112)? mem[130] :
                        (N114)? mem[194] :
                        (N116)? mem[258] :
                        (N118)? mem[322] :
                        (N120)? mem[386] :
                        (N122)? mem[450] :
                        (N124)? mem[514] :
                        (N126)? mem[578] :
                        (N128)? mem[642] :
                        (N130)? mem[706] :
                        (N132)? mem[770] :
                        (N134)? mem[834] :
                        (N136)? mem[898] :
                        (N138)? mem[962] :
                        (N109)? mem[1026] :
                        (N111)? mem[1090] :
                        (N113)? mem[1154] :
                        (N115)? mem[1218] :
                        (N117)? mem[1282] :
                        (N119)? mem[1346] :
                        (N121)? mem[1410] :
                        (N123)? mem[1474] :
                        (N125)? mem[1538] :
                        (N127)? mem[1602] :
                        (N129)? mem[1666] :
                        (N131)? mem[1730] :
                        (N133)? mem[1794] :
                        (N135)? mem[1858] :
                        (N137)? mem[1922] :
                        (N139)? mem[1986] : 1'b0;
  assign r1_data_o[1] = (N108)? mem[1] :
                        (N110)? mem[65] :
                        (N112)? mem[129] :
                        (N114)? mem[193] :
                        (N116)? mem[257] :
                        (N118)? mem[321] :
                        (N120)? mem[385] :
                        (N122)? mem[449] :
                        (N124)? mem[513] :
                        (N126)? mem[577] :
                        (N128)? mem[641] :
                        (N130)? mem[705] :
                        (N132)? mem[769] :
                        (N134)? mem[833] :
                        (N136)? mem[897] :
                        (N138)? mem[961] :
                        (N109)? mem[1025] :
                        (N111)? mem[1089] :
                        (N113)? mem[1153] :
                        (N115)? mem[1217] :
                        (N117)? mem[1281] :
                        (N119)? mem[1345] :
                        (N121)? mem[1409] :
                        (N123)? mem[1473] :
                        (N125)? mem[1537] :
                        (N127)? mem[1601] :
                        (N129)? mem[1665] :
                        (N131)? mem[1729] :
                        (N133)? mem[1793] :
                        (N135)? mem[1857] :
                        (N137)? mem[1921] :
                        (N139)? mem[1985] : 1'b0;
  assign r1_data_o[0] = (N108)? mem[0] :
                        (N110)? mem[64] :
                        (N112)? mem[128] :
                        (N114)? mem[192] :
                        (N116)? mem[256] :
                        (N118)? mem[320] :
                        (N120)? mem[384] :
                        (N122)? mem[448] :
                        (N124)? mem[512] :
                        (N126)? mem[576] :
                        (N128)? mem[640] :
                        (N130)? mem[704] :
                        (N132)? mem[768] :
                        (N134)? mem[832] :
                        (N136)? mem[896] :
                        (N138)? mem[960] :
                        (N109)? mem[1024] :
                        (N111)? mem[1088] :
                        (N113)? mem[1152] :
                        (N115)? mem[1216] :
                        (N117)? mem[1280] :
                        (N119)? mem[1344] :
                        (N121)? mem[1408] :
                        (N123)? mem[1472] :
                        (N125)? mem[1536] :
                        (N127)? mem[1600] :
                        (N129)? mem[1664] :
                        (N131)? mem[1728] :
                        (N133)? mem[1792] :
                        (N135)? mem[1856] :
                        (N137)? mem[1920] :
                        (N139)? mem[1984] : 1'b0;
  assign N205 = w_addr_i[3] & w_addr_i[4];
  assign N206 = N0 & w_addr_i[4];
  assign N0 = ~w_addr_i[3];
  assign N207 = w_addr_i[3] & N1;
  assign N1 = ~w_addr_i[4];
  assign N208 = N2 & N3;
  assign N2 = ~w_addr_i[3];
  assign N3 = ~w_addr_i[4];
  assign N209 = ~w_addr_i[2];
  assign N210 = w_addr_i[0] & w_addr_i[1];
  assign N211 = N4 & w_addr_i[1];
  assign N4 = ~w_addr_i[0];
  assign N212 = w_addr_i[0] & N5;
  assign N5 = ~w_addr_i[1];
  assign N213 = N6 & N7;
  assign N6 = ~w_addr_i[0];
  assign N7 = ~w_addr_i[1];
  assign N214 = w_addr_i[2] & N210;
  assign N215 = w_addr_i[2] & N211;
  assign N216 = w_addr_i[2] & N212;
  assign N217 = w_addr_i[2] & N213;
  assign N218 = N209 & N210;
  assign N219 = N209 & N211;
  assign N220 = N209 & N212;
  assign N221 = N209 & N213;
  assign N172 = N205 & N214;
  assign N171 = N205 & N215;
  assign N170 = N205 & N216;
  assign N169 = N205 & N217;
  assign N168 = N205 & N218;
  assign N167 = N205 & N219;
  assign N166 = N205 & N220;
  assign N165 = N205 & N221;
  assign N164 = N206 & N214;
  assign N163 = N206 & N215;
  assign N162 = N206 & N216;
  assign N161 = N206 & N217;
  assign N160 = N206 & N218;
  assign N159 = N206 & N219;
  assign N158 = N206 & N220;
  assign N157 = N206 & N221;
  assign N156 = N207 & N214;
  assign N155 = N207 & N215;
  assign N154 = N207 & N216;
  assign N153 = N207 & N217;
  assign N152 = N207 & N218;
  assign N151 = N207 & N219;
  assign N150 = N207 & N220;
  assign N149 = N207 & N221;
  assign N148 = N208 & N214;
  assign N147 = N208 & N215;
  assign N146 = N208 & N216;
  assign N145 = N208 & N217;
  assign N144 = N208 & N218;
  assign N143 = N208 & N219;
  assign N142 = N208 & N220;
  assign N141 = N208 & N221;
  assign { N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173 } = (N8)? { N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141 } :
                                                                                                                                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N140;
  assign N10 = ~r0_addr_r[0];
  assign N11 = ~r0_addr_r[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r0_addr_r[1];
  assign N14 = r0_addr_r[0] & N11;
  assign N15 = r0_addr_r[0] & r0_addr_r[1];
  assign N16 = ~r0_addr_r[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r0_addr_r[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r0_addr_r[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r0_addr_r[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r0_addr_r[2];
  assign N25 = ~r0_addr_r[3];
  assign N26 = N17 & N25;
  assign N27 = N17 & r0_addr_r[3];
  assign N28 = N19 & N25;
  assign N29 = N19 & r0_addr_r[3];
  assign N30 = N21 & N25;
  assign N31 = N21 & r0_addr_r[3];
  assign N32 = N23 & N25;
  assign N33 = N23 & r0_addr_r[3];
  assign N34 = N18 & N25;
  assign N35 = N18 & r0_addr_r[3];
  assign N36 = N20 & N25;
  assign N37 = N20 & r0_addr_r[3];
  assign N38 = N22 & N25;
  assign N39 = N22 & r0_addr_r[3];
  assign N40 = N24 & N25;
  assign N41 = N24 & r0_addr_r[3];
  assign N42 = ~r0_addr_r[4];
  assign N43 = N26 & N42;
  assign N44 = N26 & r0_addr_r[4];
  assign N45 = N28 & N42;
  assign N46 = N28 & r0_addr_r[4];
  assign N47 = N30 & N42;
  assign N48 = N30 & r0_addr_r[4];
  assign N49 = N32 & N42;
  assign N50 = N32 & r0_addr_r[4];
  assign N51 = N34 & N42;
  assign N52 = N34 & r0_addr_r[4];
  assign N53 = N36 & N42;
  assign N54 = N36 & r0_addr_r[4];
  assign N55 = N38 & N42;
  assign N56 = N38 & r0_addr_r[4];
  assign N57 = N40 & N42;
  assign N58 = N40 & r0_addr_r[4];
  assign N59 = N27 & N42;
  assign N60 = N27 & r0_addr_r[4];
  assign N61 = N29 & N42;
  assign N62 = N29 & r0_addr_r[4];
  assign N63 = N31 & N42;
  assign N64 = N31 & r0_addr_r[4];
  assign N65 = N33 & N42;
  assign N66 = N33 & r0_addr_r[4];
  assign N67 = N35 & N42;
  assign N68 = N35 & r0_addr_r[4];
  assign N69 = N37 & N42;
  assign N70 = N37 & r0_addr_r[4];
  assign N71 = N39 & N42;
  assign N72 = N39 & r0_addr_r[4];
  assign N73 = N41 & N42;
  assign N74 = N41 & r0_addr_r[4];
  assign N75 = ~r1_addr_r[0];
  assign N76 = ~r1_addr_r[1];
  assign N77 = N75 & N76;
  assign N78 = N75 & r1_addr_r[1];
  assign N79 = r1_addr_r[0] & N76;
  assign N80 = r1_addr_r[0] & r1_addr_r[1];
  assign N81 = ~r1_addr_r[2];
  assign N82 = N77 & N81;
  assign N83 = N77 & r1_addr_r[2];
  assign N84 = N79 & N81;
  assign N85 = N79 & r1_addr_r[2];
  assign N86 = N78 & N81;
  assign N87 = N78 & r1_addr_r[2];
  assign N88 = N80 & N81;
  assign N89 = N80 & r1_addr_r[2];
  assign N90 = ~r1_addr_r[3];
  assign N91 = N82 & N90;
  assign N92 = N82 & r1_addr_r[3];
  assign N93 = N84 & N90;
  assign N94 = N84 & r1_addr_r[3];
  assign N95 = N86 & N90;
  assign N96 = N86 & r1_addr_r[3];
  assign N97 = N88 & N90;
  assign N98 = N88 & r1_addr_r[3];
  assign N99 = N83 & N90;
  assign N100 = N83 & r1_addr_r[3];
  assign N101 = N85 & N90;
  assign N102 = N85 & r1_addr_r[3];
  assign N103 = N87 & N90;
  assign N104 = N87 & r1_addr_r[3];
  assign N105 = N89 & N90;
  assign N106 = N89 & r1_addr_r[3];
  assign N107 = ~r1_addr_r[4];
  assign N108 = N91 & N107;
  assign N109 = N91 & r1_addr_r[4];
  assign N110 = N93 & N107;
  assign N111 = N93 & r1_addr_r[4];
  assign N112 = N95 & N107;
  assign N113 = N95 & r1_addr_r[4];
  assign N114 = N97 & N107;
  assign N115 = N97 & r1_addr_r[4];
  assign N116 = N99 & N107;
  assign N117 = N99 & r1_addr_r[4];
  assign N118 = N101 & N107;
  assign N119 = N101 & r1_addr_r[4];
  assign N120 = N103 & N107;
  assign N121 = N103 & r1_addr_r[4];
  assign N122 = N105 & N107;
  assign N123 = N105 & r1_addr_r[4];
  assign N124 = N92 & N107;
  assign N125 = N92 & r1_addr_r[4];
  assign N126 = N94 & N107;
  assign N127 = N94 & r1_addr_r[4];
  assign N128 = N96 & N107;
  assign N129 = N96 & r1_addr_r[4];
  assign N130 = N98 & N107;
  assign N131 = N98 & r1_addr_r[4];
  assign N132 = N100 & N107;
  assign N133 = N100 & r1_addr_r[4];
  assign N134 = N102 & N107;
  assign N135 = N102 & r1_addr_r[4];
  assign N136 = N104 & N107;
  assign N137 = N104 & r1_addr_r[4];
  assign N138 = N106 & N107;
  assign N139 = N106 & r1_addr_r[4];
  assign N140 = ~w_v_i;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { r0_addr_r[4:0] } <= { r0_addr_i[4:0] };
      { r1_addr_r[4:0] } <= { r1_addr_i[4:0] };
    end
    if(N204) begin
      { mem[2047:1984] } <= { w_data_i[63:0] };
    end
    if(N203) begin
      { mem[1983:1920] } <= { w_data_i[63:0] };
    end
    if(N202) begin
      { mem[1919:1856] } <= { w_data_i[63:0] };
    end
    if(N201) begin
      { mem[1855:1792] } <= { w_data_i[63:0] };
    end
    if(N200) begin
      { mem[1791:1728] } <= { w_data_i[63:0] };
    end
    if(N199) begin
      { mem[1727:1664] } <= { w_data_i[63:0] };
    end
    if(N198) begin
      { mem[1663:1600] } <= { w_data_i[63:0] };
    end
    if(N197) begin
      { mem[1599:1536] } <= { w_data_i[63:0] };
    end
    if(N196) begin
      { mem[1535:1472] } <= { w_data_i[63:0] };
    end
    if(N195) begin
      { mem[1471:1408] } <= { w_data_i[63:0] };
    end
    if(N194) begin
      { mem[1407:1344] } <= { w_data_i[63:0] };
    end
    if(N193) begin
      { mem[1343:1280] } <= { w_data_i[63:0] };
    end
    if(N192) begin
      { mem[1279:1216] } <= { w_data_i[63:0] };
    end
    if(N191) begin
      { mem[1215:1152] } <= { w_data_i[63:0] };
    end
    if(N190) begin
      { mem[1151:1088] } <= { w_data_i[63:0] };
    end
    if(N189) begin
      { mem[1087:1024] } <= { w_data_i[63:0] };
    end
    if(N188) begin
      { mem[1023:960] } <= { w_data_i[63:0] };
    end
    if(N187) begin
      { mem[959:896] } <= { w_data_i[63:0] };
    end
    if(N186) begin
      { mem[895:832] } <= { w_data_i[63:0] };
    end
    if(N185) begin
      { mem[831:768] } <= { w_data_i[63:0] };
    end
    if(N184) begin
      { mem[767:704] } <= { w_data_i[63:0] };
    end
    if(N183) begin
      { mem[703:640] } <= { w_data_i[63:0] };
    end
    if(N182) begin
      { mem[639:576] } <= { w_data_i[63:0] };
    end
    if(N181) begin
      { mem[575:512] } <= { w_data_i[63:0] };
    end
    if(N180) begin
      { mem[511:448] } <= { w_data_i[63:0] };
    end
    if(N179) begin
      { mem[447:384] } <= { w_data_i[63:0] };
    end
    if(N178) begin
      { mem[383:320] } <= { w_data_i[63:0] };
    end
    if(N177) begin
      { mem[319:256] } <= { w_data_i[63:0] };
    end
    if(N176) begin
      { mem[255:192] } <= { w_data_i[63:0] };
    end
    if(N175) begin
      { mem[191:128] } <= { w_data_i[63:0] };
    end
    if(N174) begin
      { mem[127:64] } <= { w_data_i[63:0] };
    end
    if(N173) begin
      { mem[63:0] } <= { w_data_i[63:0] };
    end
  end


endmodule



module bsg_mem_2r1w_sync_width_p64_els_p32_read_write_same_addr_p1_harden_p0
(
  clk_i,
  reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r0_v_i,
  r0_addr_i,
  r0_data_o,
  r1_v_i,
  r1_addr_i,
  r1_data_o
);

  input [4:0] w_addr_i;
  input [63:0] w_data_i;
  input [4:0] r0_addr_i;
  output [63:0] r0_data_o;
  input [4:0] r1_addr_i;
  output [63:0] r1_data_o;
  input clk_i;
  input reset_i;
  input w_v_i;
  input r0_v_i;
  input r1_v_i;
  wire [63:0] r0_data_o,r1_data_o;

  bsg_mem_2r1w_sync_synth_width_p64_els_p32_read_write_same_addr_p1_harden_p0
  z_notmacro_synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r0_v_i(r0_v_i),
    .r0_addr_i(r0_addr_i),
    .r0_data_o(r0_data_o),
    .r1_v_i(r1_v_i),
    .r1_addr_i(r1_addr_i),
    .r1_data_o(r1_data_o)
  );


endmodule



module bp_be_regfile_harden_p0
(
  clk_i,
  reset_i,
  issue_v_i,
  dispatch_v_i,
  rd_w_v_i,
  rd_addr_i,
  rd_data_i,
  rs1_r_v_i,
  rs1_addr_i,
  rs1_data_o,
  rs2_r_v_i,
  rs2_addr_i,
  rs2_data_o
);

  input [4:0] rd_addr_i;
  input [63:0] rd_data_i;
  input [4:0] rs1_addr_i;
  output [63:0] rs1_data_o;
  input [4:0] rs2_addr_i;
  output [63:0] rs2_data_o;
  input clk_i;
  input reset_i;
  input issue_v_i;
  input dispatch_v_i;
  input rd_w_v_i;
  input rs1_r_v_i;
  input rs2_r_v_i;
  wire [63:0] rs1_data_o,rs2_data_o,rs1_reg_data,rs2_reg_data;
  wire N0,N1,N2,N3,N4,N5,N6,N7,rs1_read_v,rs2_read_v,rs1_issue_v,rs2_issue_v,N8,N9,N10,
  N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22;
  wire [4:0] rs1_reread_addr,rs2_reread_addr,rs1_addr_r,rs2_addr_r;

  bsg_mem_2r1w_sync_width_p64_els_p32_read_write_same_addr_p1_harden_p0
  rf
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(rd_w_v_i),
    .w_addr_i(rd_addr_i),
    .w_data_i(rd_data_i),
    .r0_v_i(rs1_read_v),
    .r0_addr_i(rs1_reread_addr),
    .r0_data_o(rs1_reg_data),
    .r1_v_i(rs2_read_v),
    .r1_addr_i(rs2_reread_addr),
    .r1_data_o(rs2_reg_data)
  );


  bsg_dff_en_width_p5
  rs1_addr
  (
    .clk_i(clk_i),
    .data_i(rs1_addr_i),
    .en_i(rs1_issue_v),
    .data_o(rs1_addr_r)
  );


  bsg_dff_en_width_p5
  rs2_addr
  (
    .clk_i(clk_i),
    .data_i(rs2_addr_i),
    .en_i(rs2_issue_v),
    .data_o(rs2_addr_r)
  );

  assign N12 = rs1_addr_r[3] | rs1_addr_r[4];
  assign N13 = rs1_addr_r[2] | N12;
  assign N14 = rs1_addr_r[1] | N13;
  assign N15 = rs1_addr_r[0] | N14;
  assign N16 = ~N15;
  assign N17 = rs2_addr_r[3] | rs2_addr_r[4];
  assign N18 = rs2_addr_r[2] | N17;
  assign N19 = rs2_addr_r[1] | N18;
  assign N20 = rs2_addr_r[0] | N19;
  assign N21 = ~N20;
  assign rs1_reread_addr = (N0)? rs1_addr_i :
                           (N1)? rs1_addr_r : 1'b0;
  assign N0 = N9;
  assign N1 = N8;
  assign rs2_reread_addr = (N2)? rs2_addr_i :
                           (N3)? rs2_addr_r : 1'b0;
  assign N2 = N11;
  assign N3 = N10;
  assign rs1_data_o = (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                      (N5)? rs1_reg_data : 1'b0;
  assign N4 = N16;
  assign N5 = N15;
  assign rs2_data_o = (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                      (N7)? rs2_reg_data : 1'b0;
  assign N6 = N21;
  assign N7 = N20;
  assign rs1_issue_v = issue_v_i & rs1_r_v_i;
  assign rs2_issue_v = issue_v_i & rs2_r_v_i;
  assign rs1_read_v = rs1_issue_v | N22;
  assign N22 = ~dispatch_v_i;
  assign rs2_read_v = rs2_issue_v | N22;
  assign N8 = ~rs1_issue_v;
  assign N9 = rs1_issue_v;
  assign N10 = ~rs2_issue_v;
  assign N11 = rs2_issue_v;

endmodule



module bsg_dff_reset_en_width_p222
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [221:0] data_i;
  output [221:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229;
  reg [221:0] data_o;
  assign { N7, N5, N3 } = (N0)? { 1'b1, 1'b1, 1'b1 } :
                          (N229)? { 1'b1, 1'b1, 1'b1 } :
                          (N2)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = reset_i;
  assign { N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N6, N4 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                (N229)? data_i : 1'b0;
  assign N1 = en_i | reset_i;
  assign N2 = ~N1;
  assign N228 = ~reset_i;
  assign N229 = en_i & N228;

  always @(posedge clk_i) begin
    if(N3) begin
      { data_o[221:123], data_o[0:0] } <= { N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N4 };
    end
    if(N5) begin
      { data_o[122:24], data_o[1:1] } <= { N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N6 };
    end
    if(N7) begin
      { data_o[23:2] } <= { N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8 };
    end
  end


endmodule



module bp_be_instr_decoder
(
  instr_i,
  decode_o,
  illegal_instr_o,
  ret_instr_o,
  csr_instr_o
);

  input [31:0] instr_i;
  output [50:0] decode_o;
  output illegal_instr_o;
  output ret_instr_o;
  output csr_instr_o;
  wire [50:0] decode_o;
  wire illegal_instr_o,ret_instr_o,csr_instr_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,
  N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,
  N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,
  N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,
  N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,
  N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,
  N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,
  N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,
  N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,
  N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,
  N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,
  N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,
  N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,
  N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,
  N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,
  N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
  N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,
  N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,
  N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,
  N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,
  N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,
  N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,
  N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,
  N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,
  N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,
  N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,
  N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,
  N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458;
  assign decode_o[50] = 1'b1;
  assign decode_o[26] = 1'b0;
  assign decode_o[28] = 1'b0;
  assign decode_o[40] = 1'b0;
  assign decode_o[42] = 1'b0;
  assign decode_o[44] = 1'b0;
  assign decode_o[47] = 1'b0;
  assign decode_o[48] = 1'b0;
  assign decode_o[49] = 1'b0;
  assign csr_instr_o = decode_o[39];
  assign ret_instr_o = decode_o[27];
  assign N65 = instr_i[1] & instr_i[0];
  assign N67 = instr_i[6] | N427;
  assign N68 = N428 | instr_i[3];
  assign N69 = N67 | N68;
  assign N70 = N69 | instr_i[2];
  assign N71 = N428 | N429;
  assign N72 = N67 | N71;
  assign N73 = N72 | instr_i[2];
  assign N75 = instr_i[6] | instr_i[5];
  assign N76 = N75 | N68;
  assign N77 = N76 | instr_i[2];
  assign N78 = N75 | N71;
  assign N79 = N78 | instr_i[2];
  assign N81 = N69 | N97;
  assign N83 = N76 | N97;
  assign N85 = N96 | N427;
  assign N86 = instr_i[4] | N429;
  assign N87 = N85 | N86;
  assign N88 = N87 | N97;
  assign N90 = instr_i[4] | instr_i[3];
  assign N91 = N85 | N90;
  assign N92 = N91 | N97;
  assign N94 = N91 | instr_i[2];
  assign N98 = N96 & N427;
  assign N99 = N428 & N429;
  assign N100 = N98 & N99;
  assign N101 = N100 & N97;
  assign N102 = N67 | N90;
  assign N103 = N102 | instr_i[2];
  assign N105 = N75 | N86;
  assign N106 = N105 | N97;
  assign N108 = N85 | N68;
  assign N109 = N108 | instr_i[2];
  assign N111 = instr_i[6] & instr_i[4];
  assign N112 = N111 & instr_i[2];
  assign N113 = N111 & instr_i[3];
  assign N114 = instr_i[4] & instr_i[3];
  assign N115 = N114 & instr_i[2];
  assign N116 = N96 & instr_i[5];
  assign N117 = N428 & instr_i[2];
  assign N118 = N116 & N117;
  assign N119 = N96 & N428;
  assign N120 = N429 & instr_i[2];
  assign N121 = N119 & N120;
  assign N122 = N427 & N428;
  assign N123 = N122 & N120;
  assign N124 = N428 & instr_i[3];
  assign N125 = N124 & N97;
  assign N126 = instr_i[6] & N427;
  assign N132 = N128 & N129;
  assign N133 = N130 & N303;
  assign N134 = N131 & N304;
  assign N135 = instr_i[4] & N97;
  assign N136 = N132 & N133;
  assign N137 = N134 & N116;
  assign N138 = N135 & N65;
  assign N139 = N136 & N137;
  assign N140 = N139 & N138;
  assign N142 = N163 & N294;
  assign N143 = N142 & N429;
  assign N144 = N142 & instr_i[3];
  assign N146 = N175 & N294;
  assign N147 = N146 & N429;
  assign N148 = N146 & instr_i[3];
  assign N150 = N163 & N295;
  assign N151 = N150 & N429;
  assign N152 = N150 & instr_i[3];
  assign N154 = N168 & N295;
  assign N155 = N154 & N429;
  assign N156 = N154 & instr_i[3];
  assign N158 = N181 & N295;
  assign N159 = N158 & N429;
  assign N160 = N158 & instr_i[3];
  assign N163 = N162 & N260;
  assign N164 = N163 & N296;
  assign N165 = N164 & N429;
  assign N166 = N163 & N297;
  assign N167 = N166 & N429;
  assign N168 = N162 & instr_i[14];
  assign N169 = N168 & N294;
  assign N170 = N169 & N429;
  assign N171 = N168 & N296;
  assign N172 = N171 & N429;
  assign N173 = N168 & N297;
  assign N174 = N173 & N429;
  assign N175 = instr_i[30] & N260;
  assign N176 = N175 & instr_i[12];
  assign N177 = instr_i[14] & N293;
  assign N178 = N177 & instr_i[3];
  assign N179 = instr_i[13] & instr_i[3];
  assign N180 = instr_i[30] & instr_i[13];
  assign N181 = instr_i[30] & instr_i[14];
  assign N182 = N181 & N293;
  assign N194 = N98 & N135;
  assign N195 = N194 & N65;
  assign N197 = N251 & N225;
  assign N198 = N293 & instr_i[3];
  assign N199 = N251 & N198;
  assign N201 = N214 & N251;
  assign N202 = N207 & N201;
  assign N203 = N202 & N227;
  assign N204 = N202 & N219;
  assign N206 = N128 & N162;
  assign N207 = N206 & N213;
  assign N208 = N207 & N216;
  assign N209 = N208 & N227;
  assign N210 = N208 & N219;
  assign N212 = N128 & instr_i[30];
  assign N213 = N129 & N130;
  assign N214 = N303 & N131;
  assign N215 = N212 & N213;
  assign N216 = N214 & N254;
  assign N217 = N215 & N216;
  assign N218 = N217 & N227;
  assign N219 = instr_i[12] & instr_i[3];
  assign N220 = N217 & N219;
  assign N222 = N261 & N225;
  assign N223 = N261 & N227;
  assign N224 = N254 & N225;
  assign N225 = N293 & N429;
  assign N226 = N257 & N225;
  assign N227 = instr_i[12] & N429;
  assign N228 = N257 & N227;
  assign N247 = instr_i[2] | N430;
  assign N248 = N247 | N431;
  assign N249 = N91 | N248;
  assign N251 = N260 & N292;
  assign N252 = N251 & N293;
  assign N253 = N251 & instr_i[12];
  assign N254 = instr_i[14] & N292;
  assign N255 = N254 & N293;
  assign N256 = N254 & instr_i[12];
  assign N257 = instr_i[14] & instr_i[13];
  assign N258 = N257 & N293;
  assign N259 = N257 & instr_i[12];
  assign N261 = N260 & instr_i[13];
  assign N272 = N75 | N90;
  assign N273 = N272 | N248;
  assign N275 = N261 & N293;
  assign N276 = N261 & instr_i[12];
  assign N285 = N260 & N96;
  assign N286 = instr_i[5] & N428;
  assign N287 = N429 & N97;
  assign N288 = N285 & N286;
  assign N289 = N287 & N65;
  assign N290 = N288 & N289;
  assign N294 = N292 & N293;
  assign N295 = N292 & instr_i[12];
  assign N296 = instr_i[13] & N293;
  assign N297 = instr_i[13] & instr_i[12];
  assign N306 = N303 & N304;
  assign N307 = N306 & N305;
  assign N310 = instr_i[26] | N309;
  assign N311 = N322 | N349;
  assign N312 = N310 | N329;
  assign N313 = N311 | N312;
  assign N314 = N313 | instr_i[20];
  assign N316 = N319 | instr_i[20];
  assign N318 = N350 | N342;
  assign N319 = N324 | N318;
  assign N320 = N319 | N338;
  assign N322 = N128 | N162;
  assign N323 = instr_i[29] | instr_i[28];
  assign N324 = N322 | N323;
  assign N325 = N324 | N353;
  assign N326 = N325 | instr_i[20];
  assign N329 = N328 | instr_i[21];
  assign N330 = N350 | N329;
  assign N331 = N352 | N330;
  assign N332 = N331 | N338;
  assign N334 = N341 | N351;
  assign N335 = N352 | N334;
  assign N336 = N335 | N338;
  assign N339 = N344 | N338;
  assign N341 = N131 | instr_i[24];
  assign N342 = instr_i[22] | instr_i[21];
  assign N343 = N341 | N342;
  assign N344 = N352 | N343;
  assign N345 = N344 | instr_i[20];
  assign N348 = instr_i[31] | instr_i[30];
  assign N349 = N129 | N130;
  assign N350 = instr_i[26] | instr_i[24];
  assign N351 = instr_i[22] | N347;
  assign N352 = N348 | N349;
  assign N353 = N350 | N351;
  assign N354 = N352 | N353;
  assign N355 = N354 | instr_i[20];
  assign N427 = ~instr_i[5];
  assign N428 = ~instr_i[4];
  assign N429 = ~instr_i[3];
  assign N430 = ~instr_i[1];
  assign N431 = ~instr_i[0];
  assign N432 = N427 | instr_i[6];
  assign N433 = N428 | N432;
  assign N434 = N429 | N433;
  assign N435 = instr_i[2] | N434;
  assign N436 = N430 | N435;
  assign N437 = N431 | N436;
  assign N438 = ~N437;
  assign N439 = instr_i[5] | instr_i[6];
  assign N440 = N428 | N439;
  assign N441 = N429 | N440;
  assign N442 = instr_i[2] | N441;
  assign N443 = N430 | N442;
  assign N444 = N431 | N443;
  assign N445 = ~N444;
  assign { N187, N186, N185, N184 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0 } :
                                      (N1)? { 1'b1, 1'b0, 1'b0, 1'b0 } :
                                      (N2)? { 1'b0, 1'b0, 1'b0, 1'b1 } :
                                      (N3)? { 1'b0, 1'b1, 1'b0, 1'b1 } :
                                      (N4)? { 1'b1, 1'b1, 1'b0, 1'b1 } :
                                      (N5)? { 1'b0, 1'b0, 1'b1, 1'b0 } :
                                      (N6)? { 1'b0, 1'b0, 1'b1, 1'b1 } :
                                      (N7)? { 1'b0, 1'b1, 1'b0, 1'b0 } :
                                      (N8)? { 1'b0, 1'b1, 1'b1, 1'b0 } :
                                      (N9)? { 1'b0, 1'b1, 1'b1, 1'b1 } :
                                      (N10)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N145;
  assign N1 = N149;
  assign N2 = N153;
  assign N3 = N157;
  assign N4 = N161;
  assign N5 = N165;
  assign N6 = N167;
  assign N7 = N170;
  assign N8 = N172;
  assign N9 = N174;
  assign N10 = N183;
  assign N188 = (N0)? 1'b0 :
                (N1)? 1'b0 :
                (N2)? 1'b0 :
                (N3)? 1'b0 :
                (N4)? 1'b0 :
                (N5)? 1'b0 :
                (N6)? 1'b0 :
                (N7)? 1'b0 :
                (N8)? 1'b0 :
                (N9)? 1'b0 :
                (N10)? 1'b1 : 1'b0;
  assign { N192, N191, N190, N189 } = (N11)? { N187, N186, N185, N184 } :
                                      (N141)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = N140;
  assign N193 = (N11)? N188 :
                (N141)? 1'b1 : 1'b0;
  assign { N240, N239, N238 } = (N12)? { 1'b0, 1'b0, 1'b0 } :
                                (N13)? { 1'b0, 1'b0, 1'b1 } :
                                (N14)? { 1'b1, 1'b0, 1'b1 } :
                                (N15)? { 1'b1, 1'b0, 1'b1 } :
                                (N16)? { 1'b0, 1'b1, 1'b0 } :
                                (N17)? { 1'b0, 1'b1, 1'b1 } :
                                (N18)? { 1'b1, 1'b0, 1'b0 } :
                                (N19)? { 1'b1, 1'b1, 1'b0 } :
                                (N20)? { 1'b1, 1'b1, 1'b1 } :
                                (N237)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = N200;
  assign N13 = N205;
  assign N14 = N211;
  assign N15 = N221;
  assign N16 = N222;
  assign N17 = N223;
  assign N18 = N224;
  assign N19 = N226;
  assign N20 = N228;
  assign N241 = (N12)? 1'b0 :
                (N13)? 1'b0 :
                (N14)? 1'b0 :
                (N15)? 1'b0 :
                (N16)? 1'b0 :
                (N17)? 1'b0 :
                (N18)? 1'b0 :
                (N19)? 1'b0 :
                (N20)? 1'b0 :
                (N237)? 1'b1 : 1'b0;
  assign { N245, N244, N243, N242 } = (N21)? { N221, N240, N239, N238 } :
                                      (N196)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N21 = N195;
  assign N246 = (N21)? N241 :
                (N196)? 1'b1 : 1'b0;
  assign { N265, N264, N263, N262 } = (N22)? { 1'b1, 1'b1, 1'b0, 1'b0 } :
                                      (N23)? { 1'b1, 1'b1, 1'b1, 1'b0 } :
                                      (N24)? { 1'b0, 1'b0, 1'b1, 1'b0 } :
                                      (N25)? { 1'b1, 1'b0, 1'b1, 1'b0 } :
                                      (N26)? { 1'b0, 1'b0, 1'b1, 1'b1 } :
                                      (N27)? { 1'b1, 1'b0, 1'b1, 1'b1 } :
                                      (N28)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N22 = N252;
  assign N23 = N253;
  assign N24 = N255;
  assign N25 = N256;
  assign N26 = N258;
  assign N27 = N259;
  assign N28 = N261;
  assign N266 = (N22)? 1'b0 :
                (N23)? 1'b0 :
                (N24)? 1'b0 :
                (N25)? 1'b0 :
                (N26)? 1'b0 :
                (N27)? 1'b0 :
                (N28)? 1'b1 : 1'b0;
  assign { N270, N269, N268, N267 } = (N29)? { N265, N264, N263, N262 } :
                                      (N30)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N29 = N250;
  assign N30 = N249;
  assign N271 = (N29)? N266 :
                (N30)? 1'b1 : 1'b0;
  assign { N279, N278, N277 } = (N22)? { 1'b0, 1'b0, 1'b0 } :
                                (N23)? { 1'b0, 1'b0, 1'b1 } :
                                (N31)? { 1'b0, 1'b1, 1'b0 } :
                                (N24)? { 1'b1, 1'b0, 1'b0 } :
                                (N25)? { 1'b1, 1'b0, 1'b1 } :
                                (N26)? { 1'b1, 1'b1, 1'b0 } :
                                (N32)? { 1'b0, 1'b1, 1'b1 } :
                                (N27)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N31 = N275;
  assign N32 = N276;
  assign N280 = (N22)? 1'b0 :
                (N23)? 1'b0 :
                (N31)? 1'b0 :
                (N24)? 1'b0 :
                (N25)? 1'b0 :
                (N26)? 1'b0 :
                (N32)? 1'b0 :
                (N27)? 1'b1 : 1'b0;
  assign { N283, N282, N281 } = (N33)? { N279, N278, N277 } :
                                (N34)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N33 = N274;
  assign N34 = N273;
  assign N284 = (N33)? N280 :
                (N34)? 1'b1 : 1'b0;
  assign { N299, N298 } = (N35)? { 1'b0, 1'b0 } :
                          (N36)? { 1'b0, 1'b1 } :
                          (N37)? { 1'b1, 1'b0 } :
                          (N38)? { 1'b1, 1'b1 } : 1'b0;
  assign N35 = N294;
  assign N36 = N295;
  assign N37 = N296;
  assign N38 = N297;
  assign { N301, N300 } = (N39)? { N299, N298 } :
                          (N291)? { 1'b0, 1'b0 } : 1'b0;
  assign N39 = N290;
  assign N302 = ~N290;
  assign N366 = (N40)? 1'b1 :
                (N41)? 1'b1 :
                (N42)? 1'b1 :
                (N43)? 1'b1 :
                (N44)? 1'b1 :
                (N45)? 1'b1 :
                (N46)? 1'b1 :
                (N47)? 1'b1 :
                (N48)? 1'b0 :
                (N365)? 1'b0 : 1'b0;
  assign N40 = N315;
  assign N41 = N317;
  assign N42 = N321;
  assign N43 = N327;
  assign N44 = N333;
  assign N45 = N337;
  assign N46 = N340;
  assign N47 = N346;
  assign N48 = N356;
  assign N367 = (N40)? 1'b0 :
                (N41)? 1'b0 :
                (N42)? 1'b0 :
                (N43)? 1'b0 :
                (N44)? 1'b0 :
                (N45)? 1'b0 :
                (N46)? 1'b0 :
                (N47)? 1'b0 :
                (N48)? 1'b0 :
                (N365)? 1'b1 : 1'b0;
  assign { N377, N376, N375, N374, N373, N372, N371, N370, N369, N368 } = (N49)? { N366, N315, N317, N321, N327, N333, N337, N340, N346, N356 } :
                                                                          (N308)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N49 = N307;
  assign N378 = (N49)? N367 :
                (N308)? 1'b1 : 1'b0;
  assign { N399, N398, N397, N385, N384, N383, N382, N381, N380, N379 } = (N50)? { 1'b1, 1'b0, 1'b1, N438, N192, N191, N190, N189, 1'b0, 1'b0 } :
                                                                          (N51)? { 1'b1, 1'b0, 1'b1, N445, N245, N244, N243, N242, 1'b1, 1'b0 } :
                                                                          (N52)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } :
                                                                          (N53)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } :
                                                                          (N54)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } :
                                                                          (N55)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } :
                                                                          (N56)? { 1'b1, 1'b0, 1'b0, 1'b0, N270, N269, N268, N267, 1'b0, 1'b0 } :
                                                                          (N57)? { 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, N283, N282, N281, 1'b0, 1'b0 } :
                                                                          (N58)? { 1'b0, 1'b1, 1'b0, 1'b0, N290, 1'b0, N301, N300, 1'b0, 1'b0 } :
                                                                          (N59)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                          (N60)? { 1'b0, 1'b1, N377, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                          (N61)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N50 = N74;
  assign N51 = N80;
  assign N52 = N82;
  assign N53 = N84;
  assign N54 = N89;
  assign N55 = N93;
  assign N56 = N95;
  assign N57 = N101;
  assign N58 = N104;
  assign N59 = N107;
  assign N60 = N110;
  assign N61 = N127;
  assign { N396, N395, N394, N393, N392, N391, N390, N389, N388, N387 } = (N60)? { N377, N376, N375, N374, N373, N372, N371, N370, N369, N368 } :
                                                                          (N386)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N400 = (N50)? N193 :
                (N51)? N246 :
                (N52)? 1'b0 :
                (N53)? 1'b0 :
                (N54)? 1'b0 :
                (N55)? 1'b0 :
                (N56)? N271 :
                (N57)? N284 :
                (N58)? N302 :
                (N59)? 1'b0 :
                (N60)? N378 :
                (N61)? 1'b1 : 1'b0;
  assign { N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401 } = (N62)? { N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N104, N101, N387, N95, N385, N384, N383, N382, N381, N84, N380, N93, N379 } :
                                                                                                                                                                    (N66)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N62 = N65;
  assign illegal_instr_o = (N62)? N400 :
                           (N66)? 1'b1 : 1'b0;
  assign { decode_o[45:45], decode_o[43:43], decode_o[41:41], decode_o[39:29], decode_o[27:27], decode_o[25:0] } = (N63)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                   (N64)? { N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N401, N410, N409, N408, N407, N406, N405, instr_i[19:15], instr_i[24:20], instr_i[11:7], N404, N403, N402, N401 } : 1'b0;
  assign N63 = decode_o[46];
  assign N64 = N426;
  assign N66 = ~N65;
  assign N74 = N446 | N447;
  assign N446 = ~N70;
  assign N447 = ~N73;
  assign N80 = N448 | N449;
  assign N448 = ~N77;
  assign N449 = ~N79;
  assign N82 = ~N81;
  assign N84 = ~N83;
  assign N89 = ~N88;
  assign N93 = ~N92;
  assign N95 = ~N94;
  assign N96 = ~instr_i[6];
  assign N97 = ~instr_i[2];
  assign N104 = ~N103;
  assign N107 = ~N106;
  assign N110 = ~N109;
  assign N127 = N112 | N455;
  assign N455 = N113 | N454;
  assign N454 = N115 | N453;
  assign N453 = N118 | N452;
  assign N452 = N121 | N451;
  assign N451 = N123 | N450;
  assign N450 = N125 | N126;
  assign N128 = ~instr_i[31];
  assign N129 = ~instr_i[29];
  assign N130 = ~instr_i[28];
  assign N131 = ~instr_i[26];
  assign N141 = ~N140;
  assign N145 = N143 | N144;
  assign N149 = N147 | N148;
  assign N153 = N151 | N152;
  assign N157 = N155 | N156;
  assign N161 = N159 | N160;
  assign N162 = ~instr_i[30];
  assign N183 = N176 | N458;
  assign N458 = N178 | N457;
  assign N457 = N179 | N456;
  assign N456 = N180 | N182;
  assign N196 = ~N195;
  assign N200 = N197 | N199;
  assign N205 = N203 | N204;
  assign N211 = N209 | N210;
  assign N221 = N218 | N220;
  assign N229 = N205 | N200;
  assign N230 = N211 | N229;
  assign N231 = N221 | N230;
  assign N232 = N222 | N231;
  assign N233 = N223 | N232;
  assign N234 = N224 | N233;
  assign N235 = N226 | N234;
  assign N236 = N228 | N235;
  assign N237 = ~N236;
  assign N250 = ~N249;
  assign N260 = ~instr_i[14];
  assign N274 = ~N273;
  assign N291 = ~N290;
  assign N292 = ~instr_i[13];
  assign N293 = ~instr_i[12];
  assign N303 = ~instr_i[27];
  assign N304 = ~instr_i[25];
  assign N305 = ~instr_i[23];
  assign N308 = ~N307;
  assign N309 = ~instr_i[24];
  assign N315 = ~N314;
  assign N317 = ~N316;
  assign N321 = ~N320;
  assign N327 = ~N326;
  assign N328 = ~instr_i[22];
  assign N333 = ~N332;
  assign N337 = ~N336;
  assign N338 = ~instr_i[20];
  assign N340 = ~N339;
  assign N346 = ~N345;
  assign N347 = ~instr_i[21];
  assign N356 = ~N355;
  assign N357 = N317 | N315;
  assign N358 = N321 | N357;
  assign N359 = N327 | N358;
  assign N360 = N333 | N359;
  assign N361 = N337 | N360;
  assign N362 = N340 | N361;
  assign N363 = N346 | N362;
  assign N364 = N356 | N363;
  assign N365 = ~N364;
  assign N386 = N109;
  assign N426 = ~illegal_instr_o;
  assign decode_o[46] = illegal_instr_o;

endmodule



module bsg_scan_width_p5_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [4:0] i;
  output [4:0] o;
  wire [4:0] o;
  wire t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__4_ = i[0] | 1'b0;
  assign t_1__3_ = i[1] | i[0];
  assign t_1__2_ = i[2] | i[1];
  assign t_1__1_ = i[3] | i[2];
  assign t_1__0_ = i[4] | i[3];
  assign t_2__4_ = t_1__4_ | 1'b0;
  assign t_2__3_ = t_1__3_ | 1'b0;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign o[0] = t_2__4_ | 1'b0;
  assign o[1] = t_2__3_ | 1'b0;
  assign o[2] = t_2__2_ | 1'b0;
  assign o[3] = t_2__1_ | 1'b0;
  assign o[4] = t_2__0_ | t_2__4_;

endmodule



module bsg_priority_encode_one_hot_out_width_p5_lo_to_hi_p1
(
  i,
  o
);

  input [4:0] i;
  output [4:0] o;
  wire [4:0] o;
  wire N0,N1,N2,N3;
  wire [4:1] scan_lo;

  bsg_scan_width_p5_or_p1_lo_to_hi_p1
  scan
  (
    .i(i),
    .o({ scan_lo, o[0:0] })
  );

  assign o[4] = scan_lo[4] & N0;
  assign N0 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N1;
  assign N1 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N2;
  assign N2 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N3;
  assign N3 = ~o[0];

endmodule



module bsg_mux_one_hot_width_p64_els_p5
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [319:0] data_i;
  input [4:0] sel_one_hot_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191;
  wire [319:0] data_masked;
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[1];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[1];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[1];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[2];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[2];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[2];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[2];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[2];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[2];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[2];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[2];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[2];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[2];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[2];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[2];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[2];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[2];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[2];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[2];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[2];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[2];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[2];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[2];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[2];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[2];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[2];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[2];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[2];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[2];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[2];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[2];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[2];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[2];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[2];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[2];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[2];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[2];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[2];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[2];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[2];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[2];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[2];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[2];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[2];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[2];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[2];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[2];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[2];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[2];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[2];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[2];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[2];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[2];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[2];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[2];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[2];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[2];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[2];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[2];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[2];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[2];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[2];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[2];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[2];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[2];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[2];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[2];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[3];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[3];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[3];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[3];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[3];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[3];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[3];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[3];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[3];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[3];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[3];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[3];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[3];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[3];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[3];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[3];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[3];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[3];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[3];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[3];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[3];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[3];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[3];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[3];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[3];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[3];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[3];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[3];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[3];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[3];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[3];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[3];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[3];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[3];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[3];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[3];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[3];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[3];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[3];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[3];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[3];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[3];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[3];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[3];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[3];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[3];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[3];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[3];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[3];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[3];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[3];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[3];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[3];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[3];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[3];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[3];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[3];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[3];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[3];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[3];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[3];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[3];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[3];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[3];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[4];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[4];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[4];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[4];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[4];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[4];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[4];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[4];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[4];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[4];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[4];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[4];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[4];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[4];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[4];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[4];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[4];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[4];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[4];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[4];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[4];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[4];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[4];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[4];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[4];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[4];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[4];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[4];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[4];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[4];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[4];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[4];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[4];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[4];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[4];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[4];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[4];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[4];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[4];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[4];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[4];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[4];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[4];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[4];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[4];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[4];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[4];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[4];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[4];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[4];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[4];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[4];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[4];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[4];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[4];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[4];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[4];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[4];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[4];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[4];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[4];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[4];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[4];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[4];
  assign data_o[0] = N2 | data_masked[0];
  assign N2 = N1 | data_masked[64];
  assign N1 = N0 | data_masked[128];
  assign N0 = data_masked[256] | data_masked[192];
  assign data_o[1] = N5 | data_masked[1];
  assign N5 = N4 | data_masked[65];
  assign N4 = N3 | data_masked[129];
  assign N3 = data_masked[257] | data_masked[193];
  assign data_o[2] = N8 | data_masked[2];
  assign N8 = N7 | data_masked[66];
  assign N7 = N6 | data_masked[130];
  assign N6 = data_masked[258] | data_masked[194];
  assign data_o[3] = N11 | data_masked[3];
  assign N11 = N10 | data_masked[67];
  assign N10 = N9 | data_masked[131];
  assign N9 = data_masked[259] | data_masked[195];
  assign data_o[4] = N14 | data_masked[4];
  assign N14 = N13 | data_masked[68];
  assign N13 = N12 | data_masked[132];
  assign N12 = data_masked[260] | data_masked[196];
  assign data_o[5] = N17 | data_masked[5];
  assign N17 = N16 | data_masked[69];
  assign N16 = N15 | data_masked[133];
  assign N15 = data_masked[261] | data_masked[197];
  assign data_o[6] = N20 | data_masked[6];
  assign N20 = N19 | data_masked[70];
  assign N19 = N18 | data_masked[134];
  assign N18 = data_masked[262] | data_masked[198];
  assign data_o[7] = N23 | data_masked[7];
  assign N23 = N22 | data_masked[71];
  assign N22 = N21 | data_masked[135];
  assign N21 = data_masked[263] | data_masked[199];
  assign data_o[8] = N26 | data_masked[8];
  assign N26 = N25 | data_masked[72];
  assign N25 = N24 | data_masked[136];
  assign N24 = data_masked[264] | data_masked[200];
  assign data_o[9] = N29 | data_masked[9];
  assign N29 = N28 | data_masked[73];
  assign N28 = N27 | data_masked[137];
  assign N27 = data_masked[265] | data_masked[201];
  assign data_o[10] = N32 | data_masked[10];
  assign N32 = N31 | data_masked[74];
  assign N31 = N30 | data_masked[138];
  assign N30 = data_masked[266] | data_masked[202];
  assign data_o[11] = N35 | data_masked[11];
  assign N35 = N34 | data_masked[75];
  assign N34 = N33 | data_masked[139];
  assign N33 = data_masked[267] | data_masked[203];
  assign data_o[12] = N38 | data_masked[12];
  assign N38 = N37 | data_masked[76];
  assign N37 = N36 | data_masked[140];
  assign N36 = data_masked[268] | data_masked[204];
  assign data_o[13] = N41 | data_masked[13];
  assign N41 = N40 | data_masked[77];
  assign N40 = N39 | data_masked[141];
  assign N39 = data_masked[269] | data_masked[205];
  assign data_o[14] = N44 | data_masked[14];
  assign N44 = N43 | data_masked[78];
  assign N43 = N42 | data_masked[142];
  assign N42 = data_masked[270] | data_masked[206];
  assign data_o[15] = N47 | data_masked[15];
  assign N47 = N46 | data_masked[79];
  assign N46 = N45 | data_masked[143];
  assign N45 = data_masked[271] | data_masked[207];
  assign data_o[16] = N50 | data_masked[16];
  assign N50 = N49 | data_masked[80];
  assign N49 = N48 | data_masked[144];
  assign N48 = data_masked[272] | data_masked[208];
  assign data_o[17] = N53 | data_masked[17];
  assign N53 = N52 | data_masked[81];
  assign N52 = N51 | data_masked[145];
  assign N51 = data_masked[273] | data_masked[209];
  assign data_o[18] = N56 | data_masked[18];
  assign N56 = N55 | data_masked[82];
  assign N55 = N54 | data_masked[146];
  assign N54 = data_masked[274] | data_masked[210];
  assign data_o[19] = N59 | data_masked[19];
  assign N59 = N58 | data_masked[83];
  assign N58 = N57 | data_masked[147];
  assign N57 = data_masked[275] | data_masked[211];
  assign data_o[20] = N62 | data_masked[20];
  assign N62 = N61 | data_masked[84];
  assign N61 = N60 | data_masked[148];
  assign N60 = data_masked[276] | data_masked[212];
  assign data_o[21] = N65 | data_masked[21];
  assign N65 = N64 | data_masked[85];
  assign N64 = N63 | data_masked[149];
  assign N63 = data_masked[277] | data_masked[213];
  assign data_o[22] = N68 | data_masked[22];
  assign N68 = N67 | data_masked[86];
  assign N67 = N66 | data_masked[150];
  assign N66 = data_masked[278] | data_masked[214];
  assign data_o[23] = N71 | data_masked[23];
  assign N71 = N70 | data_masked[87];
  assign N70 = N69 | data_masked[151];
  assign N69 = data_masked[279] | data_masked[215];
  assign data_o[24] = N74 | data_masked[24];
  assign N74 = N73 | data_masked[88];
  assign N73 = N72 | data_masked[152];
  assign N72 = data_masked[280] | data_masked[216];
  assign data_o[25] = N77 | data_masked[25];
  assign N77 = N76 | data_masked[89];
  assign N76 = N75 | data_masked[153];
  assign N75 = data_masked[281] | data_masked[217];
  assign data_o[26] = N80 | data_masked[26];
  assign N80 = N79 | data_masked[90];
  assign N79 = N78 | data_masked[154];
  assign N78 = data_masked[282] | data_masked[218];
  assign data_o[27] = N83 | data_masked[27];
  assign N83 = N82 | data_masked[91];
  assign N82 = N81 | data_masked[155];
  assign N81 = data_masked[283] | data_masked[219];
  assign data_o[28] = N86 | data_masked[28];
  assign N86 = N85 | data_masked[92];
  assign N85 = N84 | data_masked[156];
  assign N84 = data_masked[284] | data_masked[220];
  assign data_o[29] = N89 | data_masked[29];
  assign N89 = N88 | data_masked[93];
  assign N88 = N87 | data_masked[157];
  assign N87 = data_masked[285] | data_masked[221];
  assign data_o[30] = N92 | data_masked[30];
  assign N92 = N91 | data_masked[94];
  assign N91 = N90 | data_masked[158];
  assign N90 = data_masked[286] | data_masked[222];
  assign data_o[31] = N95 | data_masked[31];
  assign N95 = N94 | data_masked[95];
  assign N94 = N93 | data_masked[159];
  assign N93 = data_masked[287] | data_masked[223];
  assign data_o[32] = N98 | data_masked[32];
  assign N98 = N97 | data_masked[96];
  assign N97 = N96 | data_masked[160];
  assign N96 = data_masked[288] | data_masked[224];
  assign data_o[33] = N101 | data_masked[33];
  assign N101 = N100 | data_masked[97];
  assign N100 = N99 | data_masked[161];
  assign N99 = data_masked[289] | data_masked[225];
  assign data_o[34] = N104 | data_masked[34];
  assign N104 = N103 | data_masked[98];
  assign N103 = N102 | data_masked[162];
  assign N102 = data_masked[290] | data_masked[226];
  assign data_o[35] = N107 | data_masked[35];
  assign N107 = N106 | data_masked[99];
  assign N106 = N105 | data_masked[163];
  assign N105 = data_masked[291] | data_masked[227];
  assign data_o[36] = N110 | data_masked[36];
  assign N110 = N109 | data_masked[100];
  assign N109 = N108 | data_masked[164];
  assign N108 = data_masked[292] | data_masked[228];
  assign data_o[37] = N113 | data_masked[37];
  assign N113 = N112 | data_masked[101];
  assign N112 = N111 | data_masked[165];
  assign N111 = data_masked[293] | data_masked[229];
  assign data_o[38] = N116 | data_masked[38];
  assign N116 = N115 | data_masked[102];
  assign N115 = N114 | data_masked[166];
  assign N114 = data_masked[294] | data_masked[230];
  assign data_o[39] = N119 | data_masked[39];
  assign N119 = N118 | data_masked[103];
  assign N118 = N117 | data_masked[167];
  assign N117 = data_masked[295] | data_masked[231];
  assign data_o[40] = N122 | data_masked[40];
  assign N122 = N121 | data_masked[104];
  assign N121 = N120 | data_masked[168];
  assign N120 = data_masked[296] | data_masked[232];
  assign data_o[41] = N125 | data_masked[41];
  assign N125 = N124 | data_masked[105];
  assign N124 = N123 | data_masked[169];
  assign N123 = data_masked[297] | data_masked[233];
  assign data_o[42] = N128 | data_masked[42];
  assign N128 = N127 | data_masked[106];
  assign N127 = N126 | data_masked[170];
  assign N126 = data_masked[298] | data_masked[234];
  assign data_o[43] = N131 | data_masked[43];
  assign N131 = N130 | data_masked[107];
  assign N130 = N129 | data_masked[171];
  assign N129 = data_masked[299] | data_masked[235];
  assign data_o[44] = N134 | data_masked[44];
  assign N134 = N133 | data_masked[108];
  assign N133 = N132 | data_masked[172];
  assign N132 = data_masked[300] | data_masked[236];
  assign data_o[45] = N137 | data_masked[45];
  assign N137 = N136 | data_masked[109];
  assign N136 = N135 | data_masked[173];
  assign N135 = data_masked[301] | data_masked[237];
  assign data_o[46] = N140 | data_masked[46];
  assign N140 = N139 | data_masked[110];
  assign N139 = N138 | data_masked[174];
  assign N138 = data_masked[302] | data_masked[238];
  assign data_o[47] = N143 | data_masked[47];
  assign N143 = N142 | data_masked[111];
  assign N142 = N141 | data_masked[175];
  assign N141 = data_masked[303] | data_masked[239];
  assign data_o[48] = N146 | data_masked[48];
  assign N146 = N145 | data_masked[112];
  assign N145 = N144 | data_masked[176];
  assign N144 = data_masked[304] | data_masked[240];
  assign data_o[49] = N149 | data_masked[49];
  assign N149 = N148 | data_masked[113];
  assign N148 = N147 | data_masked[177];
  assign N147 = data_masked[305] | data_masked[241];
  assign data_o[50] = N152 | data_masked[50];
  assign N152 = N151 | data_masked[114];
  assign N151 = N150 | data_masked[178];
  assign N150 = data_masked[306] | data_masked[242];
  assign data_o[51] = N155 | data_masked[51];
  assign N155 = N154 | data_masked[115];
  assign N154 = N153 | data_masked[179];
  assign N153 = data_masked[307] | data_masked[243];
  assign data_o[52] = N158 | data_masked[52];
  assign N158 = N157 | data_masked[116];
  assign N157 = N156 | data_masked[180];
  assign N156 = data_masked[308] | data_masked[244];
  assign data_o[53] = N161 | data_masked[53];
  assign N161 = N160 | data_masked[117];
  assign N160 = N159 | data_masked[181];
  assign N159 = data_masked[309] | data_masked[245];
  assign data_o[54] = N164 | data_masked[54];
  assign N164 = N163 | data_masked[118];
  assign N163 = N162 | data_masked[182];
  assign N162 = data_masked[310] | data_masked[246];
  assign data_o[55] = N167 | data_masked[55];
  assign N167 = N166 | data_masked[119];
  assign N166 = N165 | data_masked[183];
  assign N165 = data_masked[311] | data_masked[247];
  assign data_o[56] = N170 | data_masked[56];
  assign N170 = N169 | data_masked[120];
  assign N169 = N168 | data_masked[184];
  assign N168 = data_masked[312] | data_masked[248];
  assign data_o[57] = N173 | data_masked[57];
  assign N173 = N172 | data_masked[121];
  assign N172 = N171 | data_masked[185];
  assign N171 = data_masked[313] | data_masked[249];
  assign data_o[58] = N176 | data_masked[58];
  assign N176 = N175 | data_masked[122];
  assign N175 = N174 | data_masked[186];
  assign N174 = data_masked[314] | data_masked[250];
  assign data_o[59] = N179 | data_masked[59];
  assign N179 = N178 | data_masked[123];
  assign N178 = N177 | data_masked[187];
  assign N177 = data_masked[315] | data_masked[251];
  assign data_o[60] = N182 | data_masked[60];
  assign N182 = N181 | data_masked[124];
  assign N181 = N180 | data_masked[188];
  assign N180 = data_masked[316] | data_masked[252];
  assign data_o[61] = N185 | data_masked[61];
  assign N185 = N184 | data_masked[125];
  assign N184 = N183 | data_masked[189];
  assign N183 = data_masked[317] | data_masked[253];
  assign data_o[62] = N188 | data_masked[62];
  assign N188 = N187 | data_masked[126];
  assign N187 = N186 | data_masked[190];
  assign N186 = data_masked[318] | data_masked[254];
  assign data_o[63] = N191 | data_masked[63];
  assign N191 = N190 | data_masked[127];
  assign N190 = N189 | data_masked[191];
  assign N189 = data_masked[319] | data_masked[255];

endmodule



module bsg_crossbar_o_by_i_i_els_p5_o_els_p1_width_p64
(
  i,
  sel_oi_one_hot_i,
  o
);

  input [319:0] i;
  input [4:0] sel_oi_one_hot_i;
  output [63:0] o;
  wire [63:0] o;

  bsg_mux_one_hot_width_p64_els_p5
  genblk1_0__mux_one_hot
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i),
    .data_o(o)
  );


endmodule



module bp_be_bypass_fwd_els_p4
(
  id_rs1_v_i,
  id_rs1_addr_i,
  id_rs1_i,
  id_rs2_v_i,
  id_rs2_addr_i,
  id_rs2_i,
  fwd_rd_v_i,
  fwd_rd_addr_i,
  fwd_rd_i,
  bypass_rs1_o,
  bypass_rs2_o
);

  input [4:0] id_rs1_addr_i;
  input [63:0] id_rs1_i;
  input [4:0] id_rs2_addr_i;
  input [63:0] id_rs2_i;
  input [3:0] fwd_rd_v_i;
  input [19:0] fwd_rd_addr_i;
  input [255:0] fwd_rd_i;
  output [63:0] bypass_rs1_o;
  output [63:0] bypass_rs2_o;
  input id_rs1_v_i;
  input id_rs2_v_i;
  wire [63:0] bypass_rs1_o,bypass_rs2_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55;
  wire [3:0] rs1_match_vector,rs2_match_vector;
  wire [4:0] rs1_match_vector_onehot,rs2_match_vector_onehot;

  bsg_priority_encode_one_hot_out_width_p5_lo_to_hi_p1
  bypass_match_one_hot_rs1
  (
    .i({ 1'b1, rs1_match_vector }),
    .o(rs1_match_vector_onehot)
  );


  bsg_priority_encode_one_hot_out_width_p5_lo_to_hi_p1
  bypass_match_one_hot_rs2
  (
    .i({ 1'b1, rs2_match_vector }),
    .o(rs2_match_vector_onehot)
  );


  bsg_crossbar_o_by_i_i_els_p5_o_els_p1_width_p64
  bypass_rs1_crossbar
  (
    .i({ id_rs1_i, fwd_rd_i }),
    .sel_oi_one_hot_i(rs1_match_vector_onehot),
    .o(bypass_rs1_o)
  );


  bsg_crossbar_o_by_i_i_els_p5_o_els_p1_width_p64
  bypass_rs2_crossbar
  (
    .i({ id_rs2_i, fwd_rd_i }),
    .sel_oi_one_hot_i(rs2_match_vector_onehot),
    .o(bypass_rs2_o)
  );

  assign N0 = id_rs1_addr_i == fwd_rd_addr_i[4:0];
  assign N1 = id_rs2_addr_i == fwd_rd_addr_i[4:0];
  assign N2 = id_rs1_addr_i == fwd_rd_addr_i[9:5];
  assign N3 = id_rs2_addr_i == fwd_rd_addr_i[9:5];
  assign N4 = id_rs1_addr_i == fwd_rd_addr_i[14:10];
  assign N5 = id_rs2_addr_i == fwd_rd_addr_i[14:10];
  assign N6 = id_rs1_addr_i == fwd_rd_addr_i[19:15];
  assign N7 = id_rs2_addr_i == fwd_rd_addr_i[19:15];
  assign N8 = id_rs1_addr_i[3] | id_rs1_addr_i[4];
  assign N9 = id_rs1_addr_i[2] | N8;
  assign N10 = id_rs1_addr_i[1] | N9;
  assign N11 = id_rs1_addr_i[0] | N10;
  assign N12 = id_rs1_addr_i[3] | id_rs1_addr_i[4];
  assign N13 = id_rs1_addr_i[2] | N12;
  assign N14 = id_rs1_addr_i[1] | N13;
  assign N15 = id_rs1_addr_i[0] | N14;
  assign N16 = id_rs1_addr_i[3] | id_rs1_addr_i[4];
  assign N17 = id_rs1_addr_i[2] | N16;
  assign N18 = id_rs1_addr_i[1] | N17;
  assign N19 = id_rs1_addr_i[0] | N18;
  assign N20 = id_rs1_addr_i[3] | id_rs1_addr_i[4];
  assign N21 = id_rs1_addr_i[2] | N20;
  assign N22 = id_rs1_addr_i[1] | N21;
  assign N23 = id_rs1_addr_i[0] | N22;
  assign N24 = id_rs2_addr_i[3] | id_rs2_addr_i[4];
  assign N25 = id_rs2_addr_i[2] | N24;
  assign N26 = id_rs2_addr_i[1] | N25;
  assign N27 = id_rs2_addr_i[0] | N26;
  assign N28 = id_rs2_addr_i[3] | id_rs2_addr_i[4];
  assign N29 = id_rs2_addr_i[2] | N28;
  assign N30 = id_rs2_addr_i[1] | N29;
  assign N31 = id_rs2_addr_i[0] | N30;
  assign N32 = id_rs2_addr_i[3] | id_rs2_addr_i[4];
  assign N33 = id_rs2_addr_i[2] | N32;
  assign N34 = id_rs2_addr_i[1] | N33;
  assign N35 = id_rs2_addr_i[0] | N34;
  assign N36 = id_rs2_addr_i[3] | id_rs2_addr_i[4];
  assign N37 = id_rs2_addr_i[2] | N36;
  assign N38 = id_rs2_addr_i[1] | N37;
  assign N39 = id_rs2_addr_i[0] | N38;
  assign rs1_match_vector[0] = N41 & N23;
  assign N41 = N0 & N40;
  assign N40 = id_rs1_v_i & fwd_rd_v_i[0];
  assign rs2_match_vector[0] = N43 & N39;
  assign N43 = N1 & N42;
  assign N42 = id_rs2_v_i & fwd_rd_v_i[0];
  assign rs1_match_vector[1] = N45 & N19;
  assign N45 = N2 & N44;
  assign N44 = id_rs1_v_i & fwd_rd_v_i[1];
  assign rs2_match_vector[1] = N47 & N35;
  assign N47 = N3 & N46;
  assign N46 = id_rs2_v_i & fwd_rd_v_i[1];
  assign rs1_match_vector[2] = N49 & N15;
  assign N49 = N4 & N48;
  assign N48 = id_rs1_v_i & fwd_rd_v_i[2];
  assign rs2_match_vector[2] = N51 & N31;
  assign N51 = N5 & N50;
  assign N50 = id_rs2_v_i & fwd_rd_v_i[2];
  assign rs1_match_vector[3] = N53 & N11;
  assign N53 = N6 & N52;
  assign N52 = id_rs1_v_i & fwd_rd_v_i[3];
  assign rs2_match_vector[3] = N55 & N27;
  assign N55 = N7 & N54;
  assign N54 = id_rs2_v_i & fwd_rd_v_i[3];

endmodule



module bp_be_int_alu
(
  src1_i,
  src2_i,
  op_i,
  opw_v_i,
  result_o
);

  input [63:0] src1_i;
  input [63:0] src2_i;
  input [3:0] op_i;
  output [63:0] result_o;
  input opw_v_i;
  wire [63:0] result_o,result_sgn;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795;
  wire [31:0] resultw_sgn;
  assign N27 = N231 & N35;
  assign N28 = N272 | op_i[0];
  assign N30 = N248 | N35;
  assign N32 = N237 | N35;
  assign N34 = N256 & op_i[0];
  assign N36 = N272 | N35;
  assign N37 = op_i[2] & N35;
  assign { N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103 } = src1_i[31:0] << src2_i[4:0];
  assign { N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135 } = src1_i[31:0] >> src2_i[4:0];
  assign { N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167 } = $signed(src1_i[31:0]) >>> src2_i[4:0];
  assign N231 = N271 & N236;
  assign N232 = N241 & N35;
  assign N233 = N231 & N232;
  assign N234 = N272 | N238;
  assign N237 = op_i[3] | N236;
  assign N238 = op_i[1] | op_i[0];
  assign N239 = N237 | N238;
  assign N242 = N241 | op_i[0];
  assign N243 = N237 | N242;
  assign N245 = N241 | N35;
  assign N246 = N237 | N245;
  assign N248 = op_i[3] | op_i[2];
  assign N249 = N248 | N273;
  assign N251 = N237 | N273;
  assign N253 = N271 | N236;
  assign N254 = N253 | N273;
  assign N256 = op_i[3] & op_i[2];
  assign N257 = op_i[1] & op_i[0];
  assign N258 = N256 & N257;
  assign N259 = N248 | N242;
  assign N261 = N272 | N242;
  assign N263 = N253 | N238;
  assign N265 = N253 | N242;
  assign N267 = N248 | N245;
  assign N269 = N272 | N245;
  assign N272 = N271 | op_i[2];
  assign N273 = op_i[1] | N35;
  assign N274 = N272 | N273;
  assign { N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596 } = src1_i << src2_i[5:0];
  assign { N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660 } = src1_i >> src2_i[5:0];
  assign { N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724 } = $signed(src1_i) >>> src2_i[5:0];
  assign N788 = $signed(src1_i) < $signed(src2_i);
  assign N789 = $signed(src1_i) >= $signed(src2_i);
  assign N790 = src1_i == src2_i;
  assign N791 = src1_i != src2_i;
  assign N792 = src1_i < src2_i;
  assign N793 = src1_i >= src2_i;
  assign { N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276 } = $signed(src1_i) + $signed(src2_i);
  assign { N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39 } = $signed(src1_i[31:0]) + $signed(src2_i[31:0]);
  assign { N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340 } = $signed(src1_i) - $signed(src2_i);
  assign { N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71 } = $signed(src1_i[31:0]) - $signed(src2_i[31:0]);
  assign { N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199 } = (N0)? { N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39 } :
                                                                                                                                                                                                              (N1)? { N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71 } :
                                                                                                                                                                                                              (N2)? { N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103 } :
                                                                                                                                                                                                              (N3)? { N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135 } :
                                                                                                                                                                                                              (N4)? { N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167 } :
                                                                                                                                                                                                              (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N27;
  assign N1 = N29;
  assign N2 = N31;
  assign N3 = N33;
  assign N4 = N34;
  assign N5 = N38;
  assign resultw_sgn = (N6)? { N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199 } :
                       (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N6 = N241;
  assign N7 = op_i[1];
  assign result_sgn = (N8)? { N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276 } :
                      (N9)? { N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340 } :
                      (N10)? { N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467 } :
                      (N11)? { N468, N469, N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530, N531 } :
                      (N12)? { N532, N533, N534, N535, N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595 } :
                      (N13)? { N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596 } :
                      (N14)? { N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660 } :
                      (N15)? { N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724 } :
                      (N16)? src2_i :
                      (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N788 } :
                      (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N789 } :
                      (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N790 } :
                      (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N791 } :
                      (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N792 } :
                      (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N793 } :
                      (N23)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = N233;
  assign N9 = N235;
  assign N10 = N240;
  assign N11 = N244;
  assign N12 = N247;
  assign N13 = N250;
  assign N14 = N252;
  assign N15 = N255;
  assign N16 = N258;
  assign N17 = N260;
  assign N18 = N262;
  assign N19 = N264;
  assign N20 = N266;
  assign N21 = N268;
  assign N22 = N270;
  assign N23 = N275;
  assign result_o = (N24)? { resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn[31:31], resultw_sgn } :
                    (N25)? result_sgn : 1'b0;
  assign N24 = opw_v_i;
  assign N25 = N794;
  assign N26 = N241;
  assign N29 = ~N28;
  assign N31 = ~N30;
  assign N33 = ~N32;
  assign N35 = ~op_i[0];
  assign N38 = N795 | N37;
  assign N795 = ~N36;
  assign N235 = ~N234;
  assign N236 = ~op_i[2];
  assign N240 = ~N239;
  assign N241 = ~op_i[1];
  assign N244 = ~N243;
  assign N247 = ~N246;
  assign N250 = ~N249;
  assign N252 = ~N251;
  assign N255 = ~N254;
  assign N260 = ~N259;
  assign N262 = ~N261;
  assign N264 = ~N263;
  assign N266 = ~N265;
  assign N268 = ~N267;
  assign N270 = ~N269;
  assign N271 = ~op_i[3];
  assign N275 = ~N274;
  assign N404 = src1_i[63] ^ src2_i[63];
  assign N405 = src1_i[62] ^ src2_i[62];
  assign N406 = src1_i[61] ^ src2_i[61];
  assign N407 = src1_i[60] ^ src2_i[60];
  assign N408 = src1_i[59] ^ src2_i[59];
  assign N409 = src1_i[58] ^ src2_i[58];
  assign N410 = src1_i[57] ^ src2_i[57];
  assign N411 = src1_i[56] ^ src2_i[56];
  assign N412 = src1_i[55] ^ src2_i[55];
  assign N413 = src1_i[54] ^ src2_i[54];
  assign N414 = src1_i[53] ^ src2_i[53];
  assign N415 = src1_i[52] ^ src2_i[52];
  assign N416 = src1_i[51] ^ src2_i[51];
  assign N417 = src1_i[50] ^ src2_i[50];
  assign N418 = src1_i[49] ^ src2_i[49];
  assign N419 = src1_i[48] ^ src2_i[48];
  assign N420 = src1_i[47] ^ src2_i[47];
  assign N421 = src1_i[46] ^ src2_i[46];
  assign N422 = src1_i[45] ^ src2_i[45];
  assign N423 = src1_i[44] ^ src2_i[44];
  assign N424 = src1_i[43] ^ src2_i[43];
  assign N425 = src1_i[42] ^ src2_i[42];
  assign N426 = src1_i[41] ^ src2_i[41];
  assign N427 = src1_i[40] ^ src2_i[40];
  assign N428 = src1_i[39] ^ src2_i[39];
  assign N429 = src1_i[38] ^ src2_i[38];
  assign N430 = src1_i[37] ^ src2_i[37];
  assign N431 = src1_i[36] ^ src2_i[36];
  assign N432 = src1_i[35] ^ src2_i[35];
  assign N433 = src1_i[34] ^ src2_i[34];
  assign N434 = src1_i[33] ^ src2_i[33];
  assign N435 = src1_i[32] ^ src2_i[32];
  assign N436 = src1_i[31] ^ src2_i[31];
  assign N437 = src1_i[30] ^ src2_i[30];
  assign N438 = src1_i[29] ^ src2_i[29];
  assign N439 = src1_i[28] ^ src2_i[28];
  assign N440 = src1_i[27] ^ src2_i[27];
  assign N441 = src1_i[26] ^ src2_i[26];
  assign N442 = src1_i[25] ^ src2_i[25];
  assign N443 = src1_i[24] ^ src2_i[24];
  assign N444 = src1_i[23] ^ src2_i[23];
  assign N445 = src1_i[22] ^ src2_i[22];
  assign N446 = src1_i[21] ^ src2_i[21];
  assign N447 = src1_i[20] ^ src2_i[20];
  assign N448 = src1_i[19] ^ src2_i[19];
  assign N449 = src1_i[18] ^ src2_i[18];
  assign N450 = src1_i[17] ^ src2_i[17];
  assign N451 = src1_i[16] ^ src2_i[16];
  assign N452 = src1_i[15] ^ src2_i[15];
  assign N453 = src1_i[14] ^ src2_i[14];
  assign N454 = src1_i[13] ^ src2_i[13];
  assign N455 = src1_i[12] ^ src2_i[12];
  assign N456 = src1_i[11] ^ src2_i[11];
  assign N457 = src1_i[10] ^ src2_i[10];
  assign N458 = src1_i[9] ^ src2_i[9];
  assign N459 = src1_i[8] ^ src2_i[8];
  assign N460 = src1_i[7] ^ src2_i[7];
  assign N461 = src1_i[6] ^ src2_i[6];
  assign N462 = src1_i[5] ^ src2_i[5];
  assign N463 = src1_i[4] ^ src2_i[4];
  assign N464 = src1_i[3] ^ src2_i[3];
  assign N465 = src1_i[2] ^ src2_i[2];
  assign N466 = src1_i[1] ^ src2_i[1];
  assign N467 = src1_i[0] ^ src2_i[0];
  assign N468 = src1_i[63] | src2_i[63];
  assign N469 = src1_i[62] | src2_i[62];
  assign N470 = src1_i[61] | src2_i[61];
  assign N471 = src1_i[60] | src2_i[60];
  assign N472 = src1_i[59] | src2_i[59];
  assign N473 = src1_i[58] | src2_i[58];
  assign N474 = src1_i[57] | src2_i[57];
  assign N475 = src1_i[56] | src2_i[56];
  assign N476 = src1_i[55] | src2_i[55];
  assign N477 = src1_i[54] | src2_i[54];
  assign N478 = src1_i[53] | src2_i[53];
  assign N479 = src1_i[52] | src2_i[52];
  assign N480 = src1_i[51] | src2_i[51];
  assign N481 = src1_i[50] | src2_i[50];
  assign N482 = src1_i[49] | src2_i[49];
  assign N483 = src1_i[48] | src2_i[48];
  assign N484 = src1_i[47] | src2_i[47];
  assign N485 = src1_i[46] | src2_i[46];
  assign N486 = src1_i[45] | src2_i[45];
  assign N487 = src1_i[44] | src2_i[44];
  assign N488 = src1_i[43] | src2_i[43];
  assign N489 = src1_i[42] | src2_i[42];
  assign N490 = src1_i[41] | src2_i[41];
  assign N491 = src1_i[40] | src2_i[40];
  assign N492 = src1_i[39] | src2_i[39];
  assign N493 = src1_i[38] | src2_i[38];
  assign N494 = src1_i[37] | src2_i[37];
  assign N495 = src1_i[36] | src2_i[36];
  assign N496 = src1_i[35] | src2_i[35];
  assign N497 = src1_i[34] | src2_i[34];
  assign N498 = src1_i[33] | src2_i[33];
  assign N499 = src1_i[32] | src2_i[32];
  assign N500 = src1_i[31] | src2_i[31];
  assign N501 = src1_i[30] | src2_i[30];
  assign N502 = src1_i[29] | src2_i[29];
  assign N503 = src1_i[28] | src2_i[28];
  assign N504 = src1_i[27] | src2_i[27];
  assign N505 = src1_i[26] | src2_i[26];
  assign N506 = src1_i[25] | src2_i[25];
  assign N507 = src1_i[24] | src2_i[24];
  assign N508 = src1_i[23] | src2_i[23];
  assign N509 = src1_i[22] | src2_i[22];
  assign N510 = src1_i[21] | src2_i[21];
  assign N511 = src1_i[20] | src2_i[20];
  assign N512 = src1_i[19] | src2_i[19];
  assign N513 = src1_i[18] | src2_i[18];
  assign N514 = src1_i[17] | src2_i[17];
  assign N515 = src1_i[16] | src2_i[16];
  assign N516 = src1_i[15] | src2_i[15];
  assign N517 = src1_i[14] | src2_i[14];
  assign N518 = src1_i[13] | src2_i[13];
  assign N519 = src1_i[12] | src2_i[12];
  assign N520 = src1_i[11] | src2_i[11];
  assign N521 = src1_i[10] | src2_i[10];
  assign N522 = src1_i[9] | src2_i[9];
  assign N523 = src1_i[8] | src2_i[8];
  assign N524 = src1_i[7] | src2_i[7];
  assign N525 = src1_i[6] | src2_i[6];
  assign N526 = src1_i[5] | src2_i[5];
  assign N527 = src1_i[4] | src2_i[4];
  assign N528 = src1_i[3] | src2_i[3];
  assign N529 = src1_i[2] | src2_i[2];
  assign N530 = src1_i[1] | src2_i[1];
  assign N531 = src1_i[0] | src2_i[0];
  assign N532 = src1_i[63] & src2_i[63];
  assign N533 = src1_i[62] & src2_i[62];
  assign N534 = src1_i[61] & src2_i[61];
  assign N535 = src1_i[60] & src2_i[60];
  assign N536 = src1_i[59] & src2_i[59];
  assign N537 = src1_i[58] & src2_i[58];
  assign N538 = src1_i[57] & src2_i[57];
  assign N539 = src1_i[56] & src2_i[56];
  assign N540 = src1_i[55] & src2_i[55];
  assign N541 = src1_i[54] & src2_i[54];
  assign N542 = src1_i[53] & src2_i[53];
  assign N543 = src1_i[52] & src2_i[52];
  assign N544 = src1_i[51] & src2_i[51];
  assign N545 = src1_i[50] & src2_i[50];
  assign N546 = src1_i[49] & src2_i[49];
  assign N547 = src1_i[48] & src2_i[48];
  assign N548 = src1_i[47] & src2_i[47];
  assign N549 = src1_i[46] & src2_i[46];
  assign N550 = src1_i[45] & src2_i[45];
  assign N551 = src1_i[44] & src2_i[44];
  assign N552 = src1_i[43] & src2_i[43];
  assign N553 = src1_i[42] & src2_i[42];
  assign N554 = src1_i[41] & src2_i[41];
  assign N555 = src1_i[40] & src2_i[40];
  assign N556 = src1_i[39] & src2_i[39];
  assign N557 = src1_i[38] & src2_i[38];
  assign N558 = src1_i[37] & src2_i[37];
  assign N559 = src1_i[36] & src2_i[36];
  assign N560 = src1_i[35] & src2_i[35];
  assign N561 = src1_i[34] & src2_i[34];
  assign N562 = src1_i[33] & src2_i[33];
  assign N563 = src1_i[32] & src2_i[32];
  assign N564 = src1_i[31] & src2_i[31];
  assign N565 = src1_i[30] & src2_i[30];
  assign N566 = src1_i[29] & src2_i[29];
  assign N567 = src1_i[28] & src2_i[28];
  assign N568 = src1_i[27] & src2_i[27];
  assign N569 = src1_i[26] & src2_i[26];
  assign N570 = src1_i[25] & src2_i[25];
  assign N571 = src1_i[24] & src2_i[24];
  assign N572 = src1_i[23] & src2_i[23];
  assign N573 = src1_i[22] & src2_i[22];
  assign N574 = src1_i[21] & src2_i[21];
  assign N575 = src1_i[20] & src2_i[20];
  assign N576 = src1_i[19] & src2_i[19];
  assign N577 = src1_i[18] & src2_i[18];
  assign N578 = src1_i[17] & src2_i[17];
  assign N579 = src1_i[16] & src2_i[16];
  assign N580 = src1_i[15] & src2_i[15];
  assign N581 = src1_i[14] & src2_i[14];
  assign N582 = src1_i[13] & src2_i[13];
  assign N583 = src1_i[12] & src2_i[12];
  assign N584 = src1_i[11] & src2_i[11];
  assign N585 = src1_i[10] & src2_i[10];
  assign N586 = src1_i[9] & src2_i[9];
  assign N587 = src1_i[8] & src2_i[8];
  assign N588 = src1_i[7] & src2_i[7];
  assign N589 = src1_i[6] & src2_i[6];
  assign N590 = src1_i[5] & src2_i[5];
  assign N591 = src1_i[4] & src2_i[4];
  assign N592 = src1_i[3] & src2_i[3];
  assign N593 = src1_i[2] & src2_i[2];
  assign N594 = src1_i[1] & src2_i[1];
  assign N595 = src1_i[0] & src2_i[0];
  assign N794 = ~opw_v_i;

endmodule



module bp_be_pipe_int
(
  clk_i,
  reset_i,
  kill_ex1_i,
  decode_i,
  pc_i,
  rs1_i,
  rs2_i,
  imm_i,
  data_o,
  br_tgt_o
);

  input [50:0] decode_i;
  input [63:0] pc_i;
  input [63:0] rs1_i;
  input [63:0] rs2_i;
  input [63:0] imm_i;
  output [63:0] data_o;
  output [63:0] br_tgt_o;
  input clk_i;
  input reset_i;
  input kill_ex1_i;
  wire [63:0] data_o,br_tgt_o,src1,src2,alu_result,baddr,pc_plus4;
  wire N0,N1,N2,N3,N4,N5,N6,N7;

  bp_be_int_alu
  alu
  (
    .src1_i(src1),
    .src2_i(src2),
    .op_i(decode_i[22:19]),
    .opw_v_i(decode_i[23]),
    .result_o(alu_result)
  );

  assign pc_plus4 = pc_i + { 1'b1, 1'b0, 1'b0 };
  assign br_tgt_o = baddr + imm_i;
  assign src1 = (N0)? pc_i :
                (N4)? rs1_i : 1'b0;
  assign N0 = decode_i[3];
  assign src2 = (N1)? imm_i :
                (N5)? rs2_i : 1'b0;
  assign N1 = decode_i[2];
  assign baddr = (N2)? src1 :
                 (N6)? pc_i : 1'b0;
  assign N2 = decode_i[1];
  assign data_o = (N3)? pc_plus4 :
                  (N7)? alu_result : 1'b0;
  assign N3 = decode_i[0];
  assign N4 = ~decode_i[3];
  assign N5 = ~decode_i[2];
  assign N6 = ~decode_i[1];
  assign N7 = ~decode_i[0];

endmodule



module bp_be_pipe_mul
(
  clk_i,
  reset_i,
  kill_ex1_i,
  kill_ex2_i,
  decode_i,
  rs1_i,
  rs2_i,
  data_o
);

  input [50:0] decode_i;
  input [63:0] rs1_i;
  input [63:0] rs2_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input kill_ex1_i;
  input kill_ex2_i;
  wire [63:0] data_o;
  assign data_o[0] = 1'b0;
  assign data_o[1] = 1'b0;
  assign data_o[2] = 1'b0;
  assign data_o[3] = 1'b0;
  assign data_o[4] = 1'b0;
  assign data_o[5] = 1'b0;
  assign data_o[6] = 1'b0;
  assign data_o[7] = 1'b0;
  assign data_o[8] = 1'b0;
  assign data_o[9] = 1'b0;
  assign data_o[10] = 1'b0;
  assign data_o[11] = 1'b0;
  assign data_o[12] = 1'b0;
  assign data_o[13] = 1'b0;
  assign data_o[14] = 1'b0;
  assign data_o[15] = 1'b0;
  assign data_o[16] = 1'b0;
  assign data_o[17] = 1'b0;
  assign data_o[18] = 1'b0;
  assign data_o[19] = 1'b0;
  assign data_o[20] = 1'b0;
  assign data_o[21] = 1'b0;
  assign data_o[22] = 1'b0;
  assign data_o[23] = 1'b0;
  assign data_o[24] = 1'b0;
  assign data_o[25] = 1'b0;
  assign data_o[26] = 1'b0;
  assign data_o[27] = 1'b0;
  assign data_o[28] = 1'b0;
  assign data_o[29] = 1'b0;
  assign data_o[30] = 1'b0;
  assign data_o[31] = 1'b0;
  assign data_o[32] = 1'b0;
  assign data_o[33] = 1'b0;
  assign data_o[34] = 1'b0;
  assign data_o[35] = 1'b0;
  assign data_o[36] = 1'b0;
  assign data_o[37] = 1'b0;
  assign data_o[38] = 1'b0;
  assign data_o[39] = 1'b0;
  assign data_o[40] = 1'b0;
  assign data_o[41] = 1'b0;
  assign data_o[42] = 1'b0;
  assign data_o[43] = 1'b0;
  assign data_o[44] = 1'b0;
  assign data_o[45] = 1'b0;
  assign data_o[46] = 1'b0;
  assign data_o[47] = 1'b0;
  assign data_o[48] = 1'b0;
  assign data_o[49] = 1'b0;
  assign data_o[50] = 1'b0;
  assign data_o[51] = 1'b0;
  assign data_o[52] = 1'b0;
  assign data_o[53] = 1'b0;
  assign data_o[54] = 1'b0;
  assign data_o[55] = 1'b0;
  assign data_o[56] = 1'b0;
  assign data_o[57] = 1'b0;
  assign data_o[58] = 1'b0;
  assign data_o[59] = 1'b0;
  assign data_o[60] = 1'b0;
  assign data_o[61] = 1'b0;
  assign data_o[62] = 1'b0;
  assign data_o[63] = 1'b0;

endmodule



module bsg_shift_reg_width_p115_stages_p2
(
  clk,
  reset_i,
  valid_i,
  data_i,
  valid_o,
  data_o
);

  input [114:0] data_i;
  output [114:0] data_o;
  input clk;
  input reset_i;
  input valid_i;
  output valid_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234;
  reg valid_o,shift_r_0__115_,shift_r_0__114_,shift_r_0__113_,shift_r_0__112_,
  shift_r_0__111_,shift_r_0__110_,shift_r_0__109_,shift_r_0__108_,shift_r_0__107_,
  shift_r_0__106_,shift_r_0__105_,shift_r_0__104_,shift_r_0__103_,shift_r_0__102_,
  shift_r_0__101_,shift_r_0__100_,shift_r_0__99_,shift_r_0__98_,shift_r_0__97_,
  shift_r_0__96_,shift_r_0__95_,shift_r_0__94_,shift_r_0__93_,shift_r_0__92_,shift_r_0__91_,
  shift_r_0__90_,shift_r_0__89_,shift_r_0__88_,shift_r_0__87_,shift_r_0__86_,
  shift_r_0__85_,shift_r_0__84_,shift_r_0__83_,shift_r_0__82_,shift_r_0__81_,
  shift_r_0__80_,shift_r_0__79_,shift_r_0__78_,shift_r_0__77_,shift_r_0__76_,shift_r_0__75_,
  shift_r_0__74_,shift_r_0__73_,shift_r_0__72_,shift_r_0__71_,shift_r_0__70_,
  shift_r_0__69_,shift_r_0__68_,shift_r_0__67_,shift_r_0__66_,shift_r_0__65_,
  shift_r_0__64_,shift_r_0__63_,shift_r_0__62_,shift_r_0__61_,shift_r_0__60_,shift_r_0__59_,
  shift_r_0__58_,shift_r_0__57_,shift_r_0__56_,shift_r_0__55_,shift_r_0__54_,
  shift_r_0__53_,shift_r_0__52_,shift_r_0__51_,shift_r_0__50_,shift_r_0__49_,
  shift_r_0__48_,shift_r_0__47_,shift_r_0__46_,shift_r_0__45_,shift_r_0__44_,shift_r_0__43_,
  shift_r_0__42_,shift_r_0__41_,shift_r_0__40_,shift_r_0__39_,shift_r_0__38_,
  shift_r_0__37_,shift_r_0__36_,shift_r_0__35_,shift_r_0__34_,shift_r_0__33_,
  shift_r_0__32_,shift_r_0__31_,shift_r_0__30_,shift_r_0__29_,shift_r_0__28_,shift_r_0__27_,
  shift_r_0__26_,shift_r_0__25_,shift_r_0__24_,shift_r_0__23_,shift_r_0__22_,
  shift_r_0__21_,shift_r_0__20_,shift_r_0__19_,shift_r_0__18_,shift_r_0__17_,
  shift_r_0__16_,shift_r_0__15_,shift_r_0__14_,shift_r_0__13_,shift_r_0__12_,shift_r_0__11_,
  shift_r_0__10_,shift_r_0__9_,shift_r_0__8_,shift_r_0__7_,shift_r_0__6_,
  shift_r_0__5_,shift_r_0__4_,shift_r_0__3_,shift_r_0__2_,shift_r_0__1_,shift_r_0__0_;
  reg [114:0] data_o;
  assign { N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N1)? { shift_r_0__115_, shift_r_0__114_, shift_r_0__113_, shift_r_0__112_, shift_r_0__111_, shift_r_0__110_, shift_r_0__109_, shift_r_0__108_, shift_r_0__107_, shift_r_0__106_, shift_r_0__105_, shift_r_0__104_, shift_r_0__103_, shift_r_0__102_, shift_r_0__101_, shift_r_0__100_, shift_r_0__99_, shift_r_0__98_, shift_r_0__97_, shift_r_0__96_, shift_r_0__95_, shift_r_0__94_, shift_r_0__93_, shift_r_0__92_, shift_r_0__91_, shift_r_0__90_, shift_r_0__89_, shift_r_0__88_, shift_r_0__87_, shift_r_0__86_, shift_r_0__85_, shift_r_0__84_, shift_r_0__83_, shift_r_0__82_, shift_r_0__81_, shift_r_0__80_, shift_r_0__79_, shift_r_0__78_, shift_r_0__77_, shift_r_0__76_, shift_r_0__75_, shift_r_0__74_, shift_r_0__73_, shift_r_0__72_, shift_r_0__71_, shift_r_0__70_, shift_r_0__69_, shift_r_0__68_, shift_r_0__67_, shift_r_0__66_, shift_r_0__65_, shift_r_0__64_, shift_r_0__63_, shift_r_0__62_, shift_r_0__61_, shift_r_0__60_, shift_r_0__59_, shift_r_0__58_, shift_r_0__57_, shift_r_0__56_, shift_r_0__55_, shift_r_0__54_, shift_r_0__53_, shift_r_0__52_, shift_r_0__51_, shift_r_0__50_, shift_r_0__49_, shift_r_0__48_, shift_r_0__47_, shift_r_0__46_, shift_r_0__45_, shift_r_0__44_, shift_r_0__43_, shift_r_0__42_, shift_r_0__41_, shift_r_0__40_, shift_r_0__39_, shift_r_0__38_, shift_r_0__37_, shift_r_0__36_, shift_r_0__35_, shift_r_0__34_, shift_r_0__33_, shift_r_0__32_, shift_r_0__31_, shift_r_0__30_, shift_r_0__29_, shift_r_0__28_, shift_r_0__27_, shift_r_0__26_, shift_r_0__25_, shift_r_0__24_, shift_r_0__23_, shift_r_0__22_, shift_r_0__21_, shift_r_0__20_, shift_r_0__19_, shift_r_0__18_, shift_r_0__17_, shift_r_0__16_, shift_r_0__15_, shift_r_0__14_, shift_r_0__13_, shift_r_0__12_, shift_r_0__11_, shift_r_0__10_, shift_r_0__9_, shift_r_0__8_, shift_r_0__7_, shift_r_0__6_, shift_r_0__5_, shift_r_0__4_, shift_r_0__3_, shift_r_0__2_, shift_r_0__1_, shift_r_0__0_, valid_i, data_i } : 1'b0;
  assign N0 = reset_i;
  assign N1 = N2;
  assign N2 = ~reset_i;

  always @(posedge clk) begin
    if(1'b1) begin
      valid_o <= N234;
      { data_o[114:0] } <= { N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119 };
      shift_r_0__115_ <= N118;
      shift_r_0__114_ <= N117;
      shift_r_0__113_ <= N116;
      shift_r_0__112_ <= N115;
      shift_r_0__111_ <= N114;
      shift_r_0__110_ <= N113;
      shift_r_0__109_ <= N112;
      shift_r_0__108_ <= N111;
      shift_r_0__107_ <= N110;
      shift_r_0__106_ <= N109;
      shift_r_0__105_ <= N108;
      shift_r_0__104_ <= N107;
      shift_r_0__103_ <= N106;
      shift_r_0__102_ <= N105;
      shift_r_0__101_ <= N104;
      shift_r_0__100_ <= N103;
      shift_r_0__99_ <= N102;
      shift_r_0__98_ <= N101;
      shift_r_0__97_ <= N100;
      shift_r_0__96_ <= N99;
      shift_r_0__95_ <= N98;
      shift_r_0__94_ <= N97;
      shift_r_0__93_ <= N96;
      shift_r_0__92_ <= N95;
      shift_r_0__91_ <= N94;
      shift_r_0__90_ <= N93;
      shift_r_0__89_ <= N92;
      shift_r_0__88_ <= N91;
      shift_r_0__87_ <= N90;
      shift_r_0__86_ <= N89;
      shift_r_0__85_ <= N88;
      shift_r_0__84_ <= N87;
      shift_r_0__83_ <= N86;
      shift_r_0__82_ <= N85;
      shift_r_0__81_ <= N84;
      shift_r_0__80_ <= N83;
      shift_r_0__79_ <= N82;
      shift_r_0__78_ <= N81;
      shift_r_0__77_ <= N80;
      shift_r_0__76_ <= N79;
      shift_r_0__75_ <= N78;
      shift_r_0__74_ <= N77;
      shift_r_0__73_ <= N76;
      shift_r_0__72_ <= N75;
      shift_r_0__71_ <= N74;
      shift_r_0__70_ <= N73;
      shift_r_0__69_ <= N72;
      shift_r_0__68_ <= N71;
      shift_r_0__67_ <= N70;
      shift_r_0__66_ <= N69;
      shift_r_0__65_ <= N68;
      shift_r_0__64_ <= N67;
      shift_r_0__63_ <= N66;
      shift_r_0__62_ <= N65;
      shift_r_0__61_ <= N64;
      shift_r_0__60_ <= N63;
      shift_r_0__59_ <= N62;
      shift_r_0__58_ <= N61;
      shift_r_0__57_ <= N60;
      shift_r_0__56_ <= N59;
      shift_r_0__55_ <= N58;
      shift_r_0__54_ <= N57;
      shift_r_0__53_ <= N56;
      shift_r_0__52_ <= N55;
      shift_r_0__51_ <= N54;
      shift_r_0__50_ <= N53;
      shift_r_0__49_ <= N52;
      shift_r_0__48_ <= N51;
      shift_r_0__47_ <= N50;
      shift_r_0__46_ <= N49;
      shift_r_0__45_ <= N48;
      shift_r_0__44_ <= N47;
      shift_r_0__43_ <= N46;
      shift_r_0__42_ <= N45;
      shift_r_0__41_ <= N44;
      shift_r_0__40_ <= N43;
      shift_r_0__39_ <= N42;
      shift_r_0__38_ <= N41;
      shift_r_0__37_ <= N40;
      shift_r_0__36_ <= N39;
      shift_r_0__35_ <= N38;
      shift_r_0__34_ <= N37;
      shift_r_0__33_ <= N36;
      shift_r_0__32_ <= N35;
      shift_r_0__31_ <= N34;
      shift_r_0__30_ <= N33;
      shift_r_0__29_ <= N32;
      shift_r_0__28_ <= N31;
      shift_r_0__27_ <= N30;
      shift_r_0__26_ <= N29;
      shift_r_0__25_ <= N28;
      shift_r_0__24_ <= N27;
      shift_r_0__23_ <= N26;
      shift_r_0__22_ <= N25;
      shift_r_0__21_ <= N24;
      shift_r_0__20_ <= N23;
      shift_r_0__19_ <= N22;
      shift_r_0__18_ <= N21;
      shift_r_0__17_ <= N20;
      shift_r_0__16_ <= N19;
      shift_r_0__15_ <= N18;
      shift_r_0__14_ <= N17;
      shift_r_0__13_ <= N16;
      shift_r_0__12_ <= N15;
      shift_r_0__11_ <= N14;
      shift_r_0__10_ <= N13;
      shift_r_0__9_ <= N12;
      shift_r_0__8_ <= N11;
      shift_r_0__7_ <= N10;
      shift_r_0__6_ <= N9;
      shift_r_0__5_ <= N8;
      shift_r_0__4_ <= N7;
      shift_r_0__3_ <= N6;
      shift_r_0__2_ <= N5;
      shift_r_0__1_ <= N4;
      shift_r_0__0_ <= N3;
    end
  end


endmodule



module bp_be_pipe_mem_vaddr_width_p39_lce_sets_p64_cce_block_size_in_bytes_p64_core_els_p1
(
  clk_i,
  reset_i,
  kill_ex1_i,
  kill_ex2_i,
  kill_ex3_i,
  decode_i,
  rs1_i,
  rs2_i,
  imm_i,
  mmu_cmd_o,
  mmu_cmd_v_o,
  mmu_cmd_ready_i,
  mmu_resp_i,
  mmu_resp_v_i,
  mmu_resp_ready_o,
  data_o,
  cache_miss_o,
  mhartid_i,
  mcycle_i,
  mtime_i,
  minstret_i,
  mtvec_o,
  mtvec_w_v_o,
  mtvec_i,
  mtval_o,
  mtval_w_v_o,
  mtval_i,
  mepc_o,
  mepc_w_v_o,
  mepc_i,
  mscratch_o,
  mscratch_w_v_o,
  mscratch_i
);

  input [50:0] decode_i;
  input [63:0] rs1_i;
  input [63:0] rs2_i;
  input [63:0] imm_i;
  output [106:0] mmu_cmd_o;
  input [72:0] mmu_resp_i;
  output [63:0] data_o;
  input [0:0] mhartid_i;
  input [63:0] mcycle_i;
  input [63:0] mtime_i;
  input [63:0] minstret_i;
  output [63:0] mtvec_o;
  input [63:0] mtvec_i;
  output [63:0] mtval_o;
  input [63:0] mtval_i;
  output [63:0] mepc_o;
  input [63:0] mepc_i;
  output [63:0] mscratch_o;
  input [63:0] mscratch_i;
  input clk_i;
  input reset_i;
  input kill_ex1_i;
  input kill_ex2_i;
  input kill_ex3_i;
  input mmu_cmd_ready_i;
  input mmu_resp_v_i;
  output mmu_cmd_v_o;
  output mmu_resp_ready_o;
  output cache_miss_o;
  output mtvec_w_v_o;
  output mtval_w_v_o;
  output mepc_w_v_o;
  output mscratch_w_v_o;
  wire [106:0] mmu_cmd_o;
  wire [63:0] data_o,mtvec_o,mtval_o,mepc_o,mscratch_o;
  wire mmu_cmd_v_o,mmu_resp_ready_o,cache_miss_o,mtvec_w_v_o,mtval_w_v_o,mepc_w_v_o,
  mscratch_w_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85;
  wire [50:0] decode_r;
  assign mmu_resp_ready_o = 1'b1;
  assign mmu_cmd_o[106] = decode_i[22];
  assign mmu_cmd_o[105] = decode_i[21];
  assign mmu_cmd_o[104] = decode_i[20];
  assign mmu_cmd_o[103] = decode_i[19];
  assign mmu_cmd_o[63] = rs2_i[63];
  assign mmu_cmd_o[62] = rs2_i[62];
  assign mmu_cmd_o[61] = rs2_i[61];
  assign mmu_cmd_o[60] = rs2_i[60];
  assign mmu_cmd_o[59] = rs2_i[59];
  assign mmu_cmd_o[58] = rs2_i[58];
  assign mmu_cmd_o[57] = rs2_i[57];
  assign mmu_cmd_o[56] = rs2_i[56];
  assign mmu_cmd_o[55] = rs2_i[55];
  assign mmu_cmd_o[54] = rs2_i[54];
  assign mmu_cmd_o[53] = rs2_i[53];
  assign mmu_cmd_o[52] = rs2_i[52];
  assign mmu_cmd_o[51] = rs2_i[51];
  assign mmu_cmd_o[50] = rs2_i[50];
  assign mmu_cmd_o[49] = rs2_i[49];
  assign mmu_cmd_o[48] = rs2_i[48];
  assign mmu_cmd_o[47] = rs2_i[47];
  assign mmu_cmd_o[46] = rs2_i[46];
  assign mmu_cmd_o[45] = rs2_i[45];
  assign mmu_cmd_o[44] = rs2_i[44];
  assign mmu_cmd_o[43] = rs2_i[43];
  assign mmu_cmd_o[42] = rs2_i[42];
  assign mmu_cmd_o[41] = rs2_i[41];
  assign mmu_cmd_o[40] = rs2_i[40];
  assign mmu_cmd_o[39] = rs2_i[39];
  assign mmu_cmd_o[38] = rs2_i[38];
  assign mmu_cmd_o[37] = rs2_i[37];
  assign mmu_cmd_o[36] = rs2_i[36];
  assign mmu_cmd_o[35] = rs2_i[35];
  assign mmu_cmd_o[34] = rs2_i[34];
  assign mmu_cmd_o[33] = rs2_i[33];
  assign mmu_cmd_o[32] = rs2_i[32];
  assign mmu_cmd_o[31] = rs2_i[31];
  assign mmu_cmd_o[30] = rs2_i[30];
  assign mmu_cmd_o[29] = rs2_i[29];
  assign mmu_cmd_o[28] = rs2_i[28];
  assign mmu_cmd_o[27] = rs2_i[27];
  assign mmu_cmd_o[26] = rs2_i[26];
  assign mmu_cmd_o[25] = rs2_i[25];
  assign mmu_cmd_o[24] = rs2_i[24];
  assign mmu_cmd_o[23] = rs2_i[23];
  assign mmu_cmd_o[22] = rs2_i[22];
  assign mmu_cmd_o[21] = rs2_i[21];
  assign mmu_cmd_o[20] = rs2_i[20];
  assign mmu_cmd_o[19] = rs2_i[19];
  assign mmu_cmd_o[18] = rs2_i[18];
  assign mmu_cmd_o[17] = rs2_i[17];
  assign mmu_cmd_o[16] = rs2_i[16];
  assign mmu_cmd_o[15] = rs2_i[15];
  assign mmu_cmd_o[14] = rs2_i[14];
  assign mmu_cmd_o[13] = rs2_i[13];
  assign mmu_cmd_o[12] = rs2_i[12];
  assign mmu_cmd_o[11] = rs2_i[11];
  assign mmu_cmd_o[10] = rs2_i[10];
  assign mmu_cmd_o[9] = rs2_i[9];
  assign mmu_cmd_o[8] = rs2_i[8];
  assign mmu_cmd_o[7] = rs2_i[7];
  assign mmu_cmd_o[6] = rs2_i[6];
  assign mmu_cmd_o[5] = rs2_i[5];
  assign mmu_cmd_o[4] = rs2_i[4];
  assign mmu_cmd_o[3] = rs2_i[3];
  assign mmu_cmd_o[2] = rs2_i[2];
  assign mmu_cmd_o[1] = rs2_i[1];
  assign mmu_cmd_o[0] = rs2_i[0];
  assign cache_miss_o = mmu_resp_i[0];
  assign mscratch_o[63] = mtvec_o[63];
  assign mepc_o[63] = mtvec_o[63];
  assign mtval_o[63] = mtvec_o[63];
  assign mscratch_o[62] = mtvec_o[62];
  assign mepc_o[62] = mtvec_o[62];
  assign mtval_o[62] = mtvec_o[62];
  assign mscratch_o[61] = mtvec_o[61];
  assign mepc_o[61] = mtvec_o[61];
  assign mtval_o[61] = mtvec_o[61];
  assign mscratch_o[60] = mtvec_o[60];
  assign mepc_o[60] = mtvec_o[60];
  assign mtval_o[60] = mtvec_o[60];
  assign mscratch_o[59] = mtvec_o[59];
  assign mepc_o[59] = mtvec_o[59];
  assign mtval_o[59] = mtvec_o[59];
  assign mscratch_o[58] = mtvec_o[58];
  assign mepc_o[58] = mtvec_o[58];
  assign mtval_o[58] = mtvec_o[58];
  assign mscratch_o[57] = mtvec_o[57];
  assign mepc_o[57] = mtvec_o[57];
  assign mtval_o[57] = mtvec_o[57];
  assign mscratch_o[56] = mtvec_o[56];
  assign mepc_o[56] = mtvec_o[56];
  assign mtval_o[56] = mtvec_o[56];
  assign mscratch_o[55] = mtvec_o[55];
  assign mepc_o[55] = mtvec_o[55];
  assign mtval_o[55] = mtvec_o[55];
  assign mscratch_o[54] = mtvec_o[54];
  assign mepc_o[54] = mtvec_o[54];
  assign mtval_o[54] = mtvec_o[54];
  assign mscratch_o[53] = mtvec_o[53];
  assign mepc_o[53] = mtvec_o[53];
  assign mtval_o[53] = mtvec_o[53];
  assign mscratch_o[52] = mtvec_o[52];
  assign mepc_o[52] = mtvec_o[52];
  assign mtval_o[52] = mtvec_o[52];
  assign mscratch_o[51] = mtvec_o[51];
  assign mepc_o[51] = mtvec_o[51];
  assign mtval_o[51] = mtvec_o[51];
  assign mscratch_o[50] = mtvec_o[50];
  assign mepc_o[50] = mtvec_o[50];
  assign mtval_o[50] = mtvec_o[50];
  assign mscratch_o[49] = mtvec_o[49];
  assign mepc_o[49] = mtvec_o[49];
  assign mtval_o[49] = mtvec_o[49];
  assign mscratch_o[48] = mtvec_o[48];
  assign mepc_o[48] = mtvec_o[48];
  assign mtval_o[48] = mtvec_o[48];
  assign mscratch_o[47] = mtvec_o[47];
  assign mepc_o[47] = mtvec_o[47];
  assign mtval_o[47] = mtvec_o[47];
  assign mscratch_o[46] = mtvec_o[46];
  assign mepc_o[46] = mtvec_o[46];
  assign mtval_o[46] = mtvec_o[46];
  assign mscratch_o[45] = mtvec_o[45];
  assign mepc_o[45] = mtvec_o[45];
  assign mtval_o[45] = mtvec_o[45];
  assign mscratch_o[44] = mtvec_o[44];
  assign mepc_o[44] = mtvec_o[44];
  assign mtval_o[44] = mtvec_o[44];
  assign mscratch_o[43] = mtvec_o[43];
  assign mepc_o[43] = mtvec_o[43];
  assign mtval_o[43] = mtvec_o[43];
  assign mscratch_o[42] = mtvec_o[42];
  assign mepc_o[42] = mtvec_o[42];
  assign mtval_o[42] = mtvec_o[42];
  assign mscratch_o[41] = mtvec_o[41];
  assign mepc_o[41] = mtvec_o[41];
  assign mtval_o[41] = mtvec_o[41];
  assign mscratch_o[40] = mtvec_o[40];
  assign mepc_o[40] = mtvec_o[40];
  assign mtval_o[40] = mtvec_o[40];
  assign mscratch_o[39] = mtvec_o[39];
  assign mepc_o[39] = mtvec_o[39];
  assign mtval_o[39] = mtvec_o[39];
  assign mscratch_o[38] = mtvec_o[38];
  assign mepc_o[38] = mtvec_o[38];
  assign mtval_o[38] = mtvec_o[38];
  assign mscratch_o[37] = mtvec_o[37];
  assign mepc_o[37] = mtvec_o[37];
  assign mtval_o[37] = mtvec_o[37];
  assign mscratch_o[36] = mtvec_o[36];
  assign mepc_o[36] = mtvec_o[36];
  assign mtval_o[36] = mtvec_o[36];
  assign mscratch_o[35] = mtvec_o[35];
  assign mepc_o[35] = mtvec_o[35];
  assign mtval_o[35] = mtvec_o[35];
  assign mscratch_o[34] = mtvec_o[34];
  assign mepc_o[34] = mtvec_o[34];
  assign mtval_o[34] = mtvec_o[34];
  assign mscratch_o[33] = mtvec_o[33];
  assign mepc_o[33] = mtvec_o[33];
  assign mtval_o[33] = mtvec_o[33];
  assign mscratch_o[32] = mtvec_o[32];
  assign mepc_o[32] = mtvec_o[32];
  assign mtval_o[32] = mtvec_o[32];
  assign mscratch_o[31] = mtvec_o[31];
  assign mepc_o[31] = mtvec_o[31];
  assign mtval_o[31] = mtvec_o[31];
  assign mscratch_o[30] = mtvec_o[30];
  assign mepc_o[30] = mtvec_o[30];
  assign mtval_o[30] = mtvec_o[30];
  assign mscratch_o[29] = mtvec_o[29];
  assign mepc_o[29] = mtvec_o[29];
  assign mtval_o[29] = mtvec_o[29];
  assign mscratch_o[28] = mtvec_o[28];
  assign mepc_o[28] = mtvec_o[28];
  assign mtval_o[28] = mtvec_o[28];
  assign mscratch_o[27] = mtvec_o[27];
  assign mepc_o[27] = mtvec_o[27];
  assign mtval_o[27] = mtvec_o[27];
  assign mscratch_o[26] = mtvec_o[26];
  assign mepc_o[26] = mtvec_o[26];
  assign mtval_o[26] = mtvec_o[26];
  assign mscratch_o[25] = mtvec_o[25];
  assign mepc_o[25] = mtvec_o[25];
  assign mtval_o[25] = mtvec_o[25];
  assign mscratch_o[24] = mtvec_o[24];
  assign mepc_o[24] = mtvec_o[24];
  assign mtval_o[24] = mtvec_o[24];
  assign mscratch_o[23] = mtvec_o[23];
  assign mepc_o[23] = mtvec_o[23];
  assign mtval_o[23] = mtvec_o[23];
  assign mscratch_o[22] = mtvec_o[22];
  assign mepc_o[22] = mtvec_o[22];
  assign mtval_o[22] = mtvec_o[22];
  assign mscratch_o[21] = mtvec_o[21];
  assign mepc_o[21] = mtvec_o[21];
  assign mtval_o[21] = mtvec_o[21];
  assign mscratch_o[20] = mtvec_o[20];
  assign mepc_o[20] = mtvec_o[20];
  assign mtval_o[20] = mtvec_o[20];
  assign mscratch_o[19] = mtvec_o[19];
  assign mepc_o[19] = mtvec_o[19];
  assign mtval_o[19] = mtvec_o[19];
  assign mscratch_o[18] = mtvec_o[18];
  assign mepc_o[18] = mtvec_o[18];
  assign mtval_o[18] = mtvec_o[18];
  assign mscratch_o[17] = mtvec_o[17];
  assign mepc_o[17] = mtvec_o[17];
  assign mtval_o[17] = mtvec_o[17];
  assign mscratch_o[16] = mtvec_o[16];
  assign mepc_o[16] = mtvec_o[16];
  assign mtval_o[16] = mtvec_o[16];
  assign mscratch_o[15] = mtvec_o[15];
  assign mepc_o[15] = mtvec_o[15];
  assign mtval_o[15] = mtvec_o[15];
  assign mscratch_o[14] = mtvec_o[14];
  assign mepc_o[14] = mtvec_o[14];
  assign mtval_o[14] = mtvec_o[14];
  assign mscratch_o[13] = mtvec_o[13];
  assign mepc_o[13] = mtvec_o[13];
  assign mtval_o[13] = mtvec_o[13];
  assign mscratch_o[12] = mtvec_o[12];
  assign mepc_o[12] = mtvec_o[12];
  assign mtval_o[12] = mtvec_o[12];
  assign mscratch_o[11] = mtvec_o[11];
  assign mepc_o[11] = mtvec_o[11];
  assign mtval_o[11] = mtvec_o[11];
  assign mscratch_o[10] = mtvec_o[10];
  assign mepc_o[10] = mtvec_o[10];
  assign mtval_o[10] = mtvec_o[10];
  assign mscratch_o[9] = mtvec_o[9];
  assign mepc_o[9] = mtvec_o[9];
  assign mtval_o[9] = mtvec_o[9];
  assign mscratch_o[8] = mtvec_o[8];
  assign mepc_o[8] = mtvec_o[8];
  assign mtval_o[8] = mtvec_o[8];
  assign mscratch_o[7] = mtvec_o[7];
  assign mepc_o[7] = mtvec_o[7];
  assign mtval_o[7] = mtvec_o[7];
  assign mscratch_o[6] = mtvec_o[6];
  assign mepc_o[6] = mtvec_o[6];
  assign mtval_o[6] = mtvec_o[6];
  assign mscratch_o[5] = mtvec_o[5];
  assign mepc_o[5] = mtvec_o[5];
  assign mtval_o[5] = mtvec_o[5];
  assign mscratch_o[4] = mtvec_o[4];
  assign mepc_o[4] = mtvec_o[4];
  assign mtval_o[4] = mtvec_o[4];
  assign mscratch_o[3] = mtvec_o[3];
  assign mepc_o[3] = mtvec_o[3];
  assign mtval_o[3] = mtvec_o[3];
  assign mscratch_o[2] = mtvec_o[2];
  assign mepc_o[2] = mtvec_o[2];
  assign mtval_o[2] = mtvec_o[2];
  assign mscratch_o[1] = mtvec_o[1];
  assign mepc_o[1] = mtvec_o[1];
  assign mtval_o[1] = mtvec_o[1];
  assign mscratch_o[0] = mtvec_o[0];
  assign mepc_o[0] = mtvec_o[0];
  assign mtval_o[0] = mtvec_o[0];

  bsg_shift_reg_width_p115_stages_p2
  csr_shift_reg
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .valid_i(1'b1),
    .data_i({ decode_i, rs1_i }),
    .data_o({ decode_r, mtvec_o })
  );

  assign mmu_cmd_o[102:64] = rs1_i[38:0] + imm_i[38:0];
  assign { N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mhartid_i[0:0] } :
                                                                                                                                                                                                                                                                                                                                              (N1)? mcycle_i :
                                                                                                                                                                                                                                                                                                                                              (N2)? mtime_i :
                                                                                                                                                                                                                                                                                                                                              (N3)? minstret_i :
                                                                                                                                                                                                                                                                                                                                              (N4)? mtvec_i :
                                                                                                                                                                                                                                                                                                                                              (N5)? mtval_i :
                                                                                                                                                                                                                                                                                                                                              (N6)? mepc_i :
                                                                                                                                                                                                                                                                                                                                              (N7)? mscratch_i :
                                                                                                                                                                                                                                                                                                                                              (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = decode_r[38];
  assign N1 = decode_r[37];
  assign N2 = decode_r[36];
  assign N3 = decode_r[35];
  assign N4 = decode_r[34];
  assign N5 = decode_r[33];
  assign N6 = decode_r[32];
  assign N7 = decode_r[31];
  assign data_o = (N8)? mmu_resp_i[72:9] :
                  (N9)? { N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19 } : 1'b0;
  assign N8 = mmu_resp_v_i;
  assign N9 = N10;
  assign mmu_cmd_v_o = N83 & N84;
  assign N83 = decode_i[29] | decode_i[30];
  assign N84 = ~kill_ex1_i;
  assign mtvec_w_v_o = decode_r[34] & N85;
  assign N85 = ~kill_ex3_i;
  assign mtval_w_v_o = decode_r[33] & N85;
  assign mepc_w_v_o = decode_r[32] & N85;
  assign mscratch_w_v_o = decode_r[31] & N85;
  assign N10 = ~mmu_resp_v_i;
  assign N11 = decode_r[37] | decode_r[38];
  assign N12 = decode_r[36] | N11;
  assign N13 = decode_r[35] | N12;
  assign N14 = decode_r[34] | N13;
  assign N15 = decode_r[33] | N14;
  assign N16 = decode_r[32] | N15;
  assign N17 = decode_r[31] | N16;
  assign N18 = ~N17;

endmodule



module bp_be_pipe_fp
(
  clk_i,
  reset_i,
  kill_ex1_i,
  kill_ex2_i,
  kill_ex3_i,
  kill_ex4_i,
  decode_i,
  rs1_i,
  rs2_i,
  data_o
);

  input [50:0] decode_i;
  input [63:0] rs1_i;
  input [63:0] rs2_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input kill_ex1_i;
  input kill_ex2_i;
  input kill_ex3_i;
  input kill_ex4_i;
  wire [63:0] data_o;
  assign data_o[0] = 1'b0;
  assign data_o[1] = 1'b0;
  assign data_o[2] = 1'b0;
  assign data_o[3] = 1'b0;
  assign data_o[4] = 1'b0;
  assign data_o[5] = 1'b0;
  assign data_o[6] = 1'b0;
  assign data_o[7] = 1'b0;
  assign data_o[8] = 1'b0;
  assign data_o[9] = 1'b0;
  assign data_o[10] = 1'b0;
  assign data_o[11] = 1'b0;
  assign data_o[12] = 1'b0;
  assign data_o[13] = 1'b0;
  assign data_o[14] = 1'b0;
  assign data_o[15] = 1'b0;
  assign data_o[16] = 1'b0;
  assign data_o[17] = 1'b0;
  assign data_o[18] = 1'b0;
  assign data_o[19] = 1'b0;
  assign data_o[20] = 1'b0;
  assign data_o[21] = 1'b0;
  assign data_o[22] = 1'b0;
  assign data_o[23] = 1'b0;
  assign data_o[24] = 1'b0;
  assign data_o[25] = 1'b0;
  assign data_o[26] = 1'b0;
  assign data_o[27] = 1'b0;
  assign data_o[28] = 1'b0;
  assign data_o[29] = 1'b0;
  assign data_o[30] = 1'b0;
  assign data_o[31] = 1'b0;
  assign data_o[32] = 1'b0;
  assign data_o[33] = 1'b0;
  assign data_o[34] = 1'b0;
  assign data_o[35] = 1'b0;
  assign data_o[36] = 1'b0;
  assign data_o[37] = 1'b0;
  assign data_o[38] = 1'b0;
  assign data_o[39] = 1'b0;
  assign data_o[40] = 1'b0;
  assign data_o[41] = 1'b0;
  assign data_o[42] = 1'b0;
  assign data_o[43] = 1'b0;
  assign data_o[44] = 1'b0;
  assign data_o[45] = 1'b0;
  assign data_o[46] = 1'b0;
  assign data_o[47] = 1'b0;
  assign data_o[48] = 1'b0;
  assign data_o[49] = 1'b0;
  assign data_o[50] = 1'b0;
  assign data_o[51] = 1'b0;
  assign data_o[52] = 1'b0;
  assign data_o[53] = 1'b0;
  assign data_o[54] = 1'b0;
  assign data_o[55] = 1'b0;
  assign data_o[56] = 1'b0;
  assign data_o[57] = 1'b0;
  assign data_o[58] = 1'b0;
  assign data_o[59] = 1'b0;
  assign data_o[60] = 1'b0;
  assign data_o[61] = 1'b0;
  assign data_o[62] = 1'b0;
  assign data_o[63] = 1'b0;

endmodule



module bsg_dff_width_p600
(
  clk_i,
  data_i,
  data_o
);

  input [599:0] data_i;
  output [599:0] data_o;
  input clk_i;
  reg [599:0] data_o;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { data_o[599:0] } <= { data_i[599:0] };
    end
  end


endmodule



module bsg_dff_width_p386
(
  clk_i,
  data_i,
  data_o
);

  input [385:0] data_i;
  output [385:0] data_o;
  input clk_i;
  reg [385:0] data_o;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { data_o[385:0] } <= { data_i[385:0] };
    end
  end


endmodule



module bsg_mux_segmented_segments_p5_segment_width_p64
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [319:0] data0_i;
  input [319:0] data1_i;
  input [4:0] sel_i;
  output [319:0] data_o;
  wire [319:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9;
  assign data_o[63:0] = (N0)? data1_i[63:0] :
                        (N5)? data0_i[63:0] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[127:64] = (N1)? data1_i[127:64] :
                          (N6)? data0_i[127:64] : 1'b0;
  assign N1 = sel_i[1];
  assign data_o[191:128] = (N2)? data1_i[191:128] :
                           (N7)? data0_i[191:128] : 1'b0;
  assign N2 = sel_i[2];
  assign data_o[255:192] = (N3)? data1_i[255:192] :
                           (N8)? data0_i[255:192] : 1'b0;
  assign N3 = sel_i[3];
  assign data_o[319:256] = (N4)? data1_i[319:256] :
                           (N9)? data0_i[319:256] : 1'b0;
  assign N4 = sel_i[4];
  assign N5 = ~sel_i[0];
  assign N6 = ~sel_i[1];
  assign N7 = ~sel_i[2];
  assign N8 = ~sel_i[3];
  assign N9 = ~sel_i[4];

endmodule



module bsg_dff_width_p320
(
  clk_i,
  data_i,
  data_o
);

  input [319:0] data_i;
  output [319:0] data_o;
  input clk_i;
  reg [319:0] data_o;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { data_o[319:0] } <= { data_i[319:0] };
    end
  end


endmodule



module bsg_dff_width_p45
(
  clk_i,
  data_i,
  data_o
);

  input [44:0] data_i;
  output [44:0] data_o;
  input clk_i;
  reg [44:0] data_o;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { data_o[44:0] } <= { data_i[44:0] };
    end
  end


endmodule



module bsg_counter_clear_up_init_val_p0_ptr_width_lp64
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [63:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197;
  reg [63:0] count_o;
  assign { N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6 } = { N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134 } + up_i;
  assign { N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                                                                                                                                                                                                                                                (N1)? { N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6 } : 1'b0;
  assign N0 = reset_i;
  assign N1 = N2;
  assign { N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134 } = count_o * N4;
  assign N2 = ~reset_i;
  assign N3 = N2;
  assign N4 = ~clear_i;
  assign N5 = N3 & N4;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { count_o[63:0] } <= { N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70 };
    end
  end


endmodule



module bp_be_calculator_top_vaddr_width_p39_paddr_width_p22_asid_width_p10_core_els_p1_num_lce_p2_lce_sets_p64_trace_p0_debug_p0_debug_file_pinv
(
  clk_i,
  reset_i,
  proc_cfg_i,
  issue_pkt_i,
  issue_pkt_v_i,
  issue_pkt_ready_o,
  chk_dispatch_v_i,
  chk_roll_i,
  chk_poison_isd_i,
  chk_poison_ex1_i,
  chk_poison_ex2_i,
  chk_poison_ex3_i,
  calc_status_o,
  mmu_cmd_o,
  mmu_cmd_v_o,
  mmu_cmd_ready_i,
  mmu_resp_i,
  mmu_resp_v_i,
  mmu_resp_ready_o,
  mtvec_o,
  mtvec_w_v_o,
  mtvec_i,
  mepc_o,
  mepc_w_v_o,
  mepc_i,
  cmt_rd_w_v_o,
  cmt_rd_addr_o,
  cmt_mem_w_v_o,
  cmt_mem_addr_o,
  cmt_mem_op_o,
  cmt_data_o
);

  input [2:0] proc_cfg_i;
  input [220:0] issue_pkt_i;
  output [306:0] calc_status_o;
  output [106:0] mmu_cmd_o;
  input [72:0] mmu_resp_i;
  output [63:0] mtvec_o;
  input [63:0] mtvec_i;
  output [63:0] mepc_o;
  input [63:0] mepc_i;
  output [4:0] cmt_rd_addr_o;
  output [63:0] cmt_mem_addr_o;
  output [3:0] cmt_mem_op_o;
  output [63:0] cmt_data_o;
  input clk_i;
  input reset_i;
  input issue_pkt_v_i;
  input chk_dispatch_v_i;
  input chk_roll_i;
  input chk_poison_isd_i;
  input chk_poison_ex1_i;
  input chk_poison_ex2_i;
  input chk_poison_ex3_i;
  input mmu_cmd_ready_i;
  input mmu_resp_v_i;
  output issue_pkt_ready_o;
  output mmu_cmd_v_o;
  output mmu_resp_ready_o;
  output mtvec_w_v_o;
  output mepc_w_v_o;
  output cmt_rd_w_v_o;
  output cmt_mem_w_v_o;
  wire [306:0] calc_status_o;
  wire [106:0] mmu_cmd_o;
  wire [63:0] mtvec_o,mepc_o,cmt_mem_addr_o,cmt_data_o,irf_rs1,irf_rs2,frf_rs1,frf_rs2,
  bypass_irs1,bypass_irs2,bypass_frs1,bypass_frs2,bypass_rs1,bypass_rs2,pipe_int_data_lo,
  pipe_mul_data_lo,cycle_cnt_lo,time_cnt_lo,instret_cnt_lo,mtval_lo,mtval_li,
  mscratch_lo,mscratch_li,pipe_mem_data_lo,pipe_fp_data_lo,mtval_mux_lo;
  wire [4:0] cmt_rd_addr_o;
  wire [3:0] cmt_mem_op_o;
  wire issue_pkt_ready_o,mmu_cmd_v_o,mmu_resp_ready_o,mtvec_w_v_o,mepc_w_v_o,
  cmt_rd_w_v_o,cmt_mem_w_v_o,N0,N1,N2,N3,N4,n_0_net_,
  calc_stage_r_4__instr_metadata__itag__7_,calc_stage_r_4__instr_metadata__itag__6_,
  calc_stage_r_4__instr_metadata__itag__5_,calc_stage_r_4__instr_metadata__itag__4_,
  calc_stage_r_4__instr_metadata__itag__3_,calc_stage_r_4__instr_metadata__itag__2_,
  calc_stage_r_4__instr_metadata__itag__1_,calc_stage_r_4__instr_metadata__itag__0_,
  calc_stage_r_4__instr_metadata__pc__63_,calc_stage_r_4__instr_metadata__pc__62_,
  calc_stage_r_4__instr_metadata__pc__61_,calc_stage_r_4__instr_metadata__pc__60_,
  calc_stage_r_4__instr_metadata__pc__59_,calc_stage_r_4__instr_metadata__pc__58_,
  calc_stage_r_4__instr_metadata__pc__57_,calc_stage_r_4__instr_metadata__pc__56_,
  calc_stage_r_4__instr_metadata__pc__55_,calc_stage_r_4__instr_metadata__pc__54_,
  calc_stage_r_4__instr_metadata__pc__53_,calc_stage_r_4__instr_metadata__pc__52_,
  calc_stage_r_4__instr_metadata__pc__51_,calc_stage_r_4__instr_metadata__pc__50_,
  calc_stage_r_4__instr_metadata__pc__49_,calc_stage_r_4__instr_metadata__pc__48_,
  calc_stage_r_4__instr_metadata__pc__47_,calc_stage_r_4__instr_metadata__pc__46_,
  calc_stage_r_4__instr_metadata__pc__45_,calc_stage_r_4__instr_metadata__pc__44_,
  calc_stage_r_4__instr_metadata__pc__43_,calc_stage_r_4__instr_metadata__pc__42_,
  calc_stage_r_4__instr_metadata__pc__41_,calc_stage_r_4__instr_metadata__pc__40_,
  calc_stage_r_4__instr_metadata__pc__39_,calc_stage_r_4__instr_metadata__pc__38_,
  calc_stage_r_4__instr_metadata__pc__37_,calc_stage_r_4__instr_metadata__pc__36_,
  calc_stage_r_4__instr_metadata__pc__35_,calc_stage_r_4__instr_metadata__pc__34_,
  calc_stage_r_4__instr_metadata__pc__33_,calc_stage_r_4__instr_metadata__pc__32_,
  calc_stage_r_4__instr_metadata__pc__31_,calc_stage_r_4__instr_metadata__pc__30_,
  calc_stage_r_4__instr_metadata__pc__29_,calc_stage_r_4__instr_metadata__pc__28_,
  calc_stage_r_4__instr_metadata__pc__27_,calc_stage_r_4__instr_metadata__pc__26_,
  calc_stage_r_4__instr_metadata__pc__25_,calc_stage_r_4__instr_metadata__pc__24_,
  calc_stage_r_4__instr_metadata__pc__23_,calc_stage_r_4__instr_metadata__pc__22_,
  calc_stage_r_4__instr_metadata__pc__21_,calc_stage_r_4__instr_metadata__pc__20_,
  calc_stage_r_4__instr_metadata__pc__19_,calc_stage_r_4__instr_metadata__pc__18_,
  calc_stage_r_4__instr_metadata__pc__17_,calc_stage_r_4__instr_metadata__pc__16_,
  calc_stage_r_4__instr_metadata__pc__15_,calc_stage_r_4__instr_metadata__pc__14_,
  calc_stage_r_4__instr_metadata__pc__13_,calc_stage_r_4__instr_metadata__pc__12_,
  calc_stage_r_4__instr_metadata__pc__11_,calc_stage_r_4__instr_metadata__pc__10_,
  calc_stage_r_4__instr_metadata__pc__9_,calc_stage_r_4__instr_metadata__pc__8_,
  calc_stage_r_4__instr_metadata__pc__7_,calc_stage_r_4__instr_metadata__pc__6_,
  calc_stage_r_4__instr_metadata__pc__5_,calc_stage_r_4__instr_metadata__pc__4_,
  calc_stage_r_4__instr_metadata__pc__3_,calc_stage_r_4__instr_metadata__pc__2_,calc_stage_r_4__instr_metadata__pc__1_,
  calc_stage_r_4__instr_metadata__pc__0_,
  calc_stage_r_4__instr_metadata__fe_exception_not_instr_,calc_stage_r_4__instr_metadata__fe_exception_code__1_,
  calc_stage_r_4__instr_metadata__fe_exception_code__0_,calc_stage_r_4__instr__31_,
  calc_stage_r_4__instr__30_,calc_stage_r_4__instr__29_,calc_stage_r_4__instr__28_,
  calc_stage_r_4__instr__27_,calc_stage_r_4__instr__26_,calc_stage_r_4__instr__25_,
  calc_stage_r_4__instr__24_,calc_stage_r_4__instr__23_,calc_stage_r_4__instr__22_,
  calc_stage_r_4__instr__21_,calc_stage_r_4__instr__20_,calc_stage_r_4__instr__19_,
  calc_stage_r_4__instr__18_,calc_stage_r_4__instr__17_,calc_stage_r_4__instr__16_,
  calc_stage_r_4__instr__15_,calc_stage_r_4__instr__14_,calc_stage_r_4__instr__13_,
  calc_stage_r_4__instr__12_,calc_stage_r_4__instr__11_,calc_stage_r_4__instr__10_,
  calc_stage_r_4__instr__9_,calc_stage_r_4__instr__8_,calc_stage_r_4__instr__7_,
  calc_stage_r_4__instr__6_,calc_stage_r_4__instr__5_,calc_stage_r_4__instr__4_,
  calc_stage_r_4__instr__3_,calc_stage_r_4__instr__2_,calc_stage_r_4__instr__1_,
  calc_stage_r_4__instr__0_,calc_stage_r_4__instr_v_,calc_stage_r_4__pipe_comp_v_,
  calc_stage_r_4__pipe_int_v_,calc_stage_r_4__pipe_mul_v_,calc_stage_r_4__pipe_mem_v_,
  calc_stage_r_4__pipe_fp_v_,calc_stage_r_4__irf_w_v_,calc_stage_r_4__frf_w_v_,
  calc_stage_r_3__instr_metadata__itag__7_,calc_stage_r_3__instr_metadata__itag__6_,
  calc_stage_r_3__instr_metadata__itag__5_,calc_stage_r_3__instr_metadata__itag__4_,
  calc_stage_r_3__instr_metadata__itag__3_,calc_stage_r_3__instr_metadata__itag__2_,
  calc_stage_r_3__instr_metadata__itag__1_,calc_stage_r_3__instr_metadata__itag__0_,
  calc_stage_r_3__instr_metadata__pc__63_,calc_stage_r_3__instr_metadata__pc__62_,
  calc_stage_r_3__instr_metadata__pc__61_,calc_stage_r_3__instr_metadata__pc__60_,
  calc_stage_r_3__instr_metadata__pc__59_,calc_stage_r_3__instr_metadata__pc__58_,
  calc_stage_r_3__instr_metadata__pc__57_,calc_stage_r_3__instr_metadata__pc__56_,
  calc_stage_r_3__instr_metadata__pc__55_,calc_stage_r_3__instr_metadata__pc__54_,
  calc_stage_r_3__instr_metadata__pc__53_,calc_stage_r_3__instr_metadata__pc__52_,
  calc_stage_r_3__instr_metadata__pc__51_,calc_stage_r_3__instr_metadata__pc__50_,
  calc_stage_r_3__instr_metadata__pc__49_,calc_stage_r_3__instr_metadata__pc__48_,
  calc_stage_r_3__instr_metadata__pc__47_,calc_stage_r_3__instr_metadata__pc__46_,
  calc_stage_r_3__instr_metadata__pc__45_,calc_stage_r_3__instr_metadata__pc__44_,
  calc_stage_r_3__instr_metadata__pc__43_,calc_stage_r_3__instr_metadata__pc__42_,
  calc_stage_r_3__instr_metadata__pc__41_,calc_stage_r_3__instr_metadata__pc__40_,
  calc_stage_r_3__instr_metadata__pc__39_,calc_stage_r_3__instr_metadata__pc__38_,
  calc_stage_r_3__instr_metadata__pc__37_,calc_stage_r_3__instr_metadata__pc__36_,
  calc_stage_r_3__instr_metadata__pc__35_,calc_stage_r_3__instr_metadata__pc__34_,
  calc_stage_r_3__instr_metadata__pc__33_,calc_stage_r_3__instr_metadata__pc__32_,
  calc_stage_r_3__instr_metadata__pc__31_,calc_stage_r_3__instr_metadata__pc__30_,
  calc_stage_r_3__instr_metadata__pc__29_,calc_stage_r_3__instr_metadata__pc__28_,
  calc_stage_r_3__instr_metadata__pc__27_,calc_stage_r_3__instr_metadata__pc__26_,
  calc_stage_r_3__instr_metadata__pc__25_,calc_stage_r_3__instr_metadata__pc__24_,
  calc_stage_r_3__instr_metadata__pc__23_,calc_stage_r_3__instr_metadata__pc__22_,
  calc_stage_r_3__instr_metadata__pc__21_,calc_stage_r_3__instr_metadata__pc__20_,
  calc_stage_r_3__instr_metadata__pc__19_,calc_stage_r_3__instr_metadata__pc__18_,
  calc_stage_r_3__instr_metadata__pc__17_,calc_stage_r_3__instr_metadata__pc__16_,
  calc_stage_r_3__instr_metadata__pc__15_,calc_stage_r_3__instr_metadata__pc__14_,
  calc_stage_r_3__instr_metadata__pc__13_,calc_stage_r_3__instr_metadata__pc__12_,
  calc_stage_r_3__instr_metadata__pc__11_,calc_stage_r_3__instr_metadata__pc__10_,
  calc_stage_r_3__instr_metadata__pc__9_,calc_stage_r_3__instr_metadata__pc__8_,
  calc_stage_r_3__instr_metadata__pc__7_,calc_stage_r_3__instr_metadata__pc__6_,
  calc_stage_r_3__instr_metadata__pc__5_,calc_stage_r_3__instr_metadata__pc__4_,
  calc_stage_r_3__instr_metadata__pc__3_,calc_stage_r_3__instr_metadata__pc__2_,
  calc_stage_r_3__instr_metadata__pc__1_,calc_stage_r_3__instr_metadata__pc__0_,
  calc_stage_r_3__instr_metadata__fe_exception_not_instr_,
  calc_stage_r_3__instr_metadata__fe_exception_code__1_,calc_stage_r_3__instr_metadata__fe_exception_code__0_,
  calc_stage_r_3__instr__31_,calc_stage_r_3__instr__30_,calc_stage_r_3__instr__29_,
  calc_stage_r_3__instr__28_,calc_stage_r_3__instr__27_,calc_stage_r_3__instr__26_,
  calc_stage_r_3__instr__25_,calc_stage_r_3__instr__24_,calc_stage_r_3__instr__23_,
  calc_stage_r_3__instr__22_,calc_stage_r_3__instr__21_,calc_stage_r_3__instr__20_,
  calc_stage_r_3__instr__19_,calc_stage_r_3__instr__18_,calc_stage_r_3__instr__17_,
  calc_stage_r_3__instr__16_,calc_stage_r_3__instr__15_,calc_stage_r_3__instr__14_,
  calc_stage_r_3__instr__13_,calc_stage_r_3__instr__12_,
  calc_stage_r_3__instr__11_,calc_stage_r_3__instr__10_,calc_stage_r_3__instr__9_,calc_stage_r_3__instr__8_,
  calc_stage_r_3__instr__7_,calc_stage_r_3__instr__6_,calc_stage_r_3__instr__5_,
  calc_stage_r_3__instr__4_,calc_stage_r_3__instr__3_,calc_stage_r_3__instr__2_,
  calc_stage_r_3__instr__1_,calc_stage_r_3__instr__0_,calc_stage_r_3__instr_v_,
  calc_stage_r_3__pipe_comp_v_,calc_stage_r_3__pipe_int_v_,calc_stage_r_3__pipe_mul_v_,
  calc_stage_r_3__pipe_mem_v_,calc_stage_r_3__pipe_fp_v_,calc_stage_r_3__irf_w_v_,
  calc_stage_r_3__frf_w_v_,calc_stage_r_2__instr_metadata__itag__7_,
  calc_stage_r_2__instr_metadata__itag__6_,calc_stage_r_2__instr_metadata__itag__5_,
  calc_stage_r_2__instr_metadata__itag__4_,calc_stage_r_2__instr_metadata__itag__3_,
  calc_stage_r_2__instr_metadata__itag__2_,calc_stage_r_2__instr_metadata__itag__1_,
  calc_stage_r_2__instr_metadata__itag__0_,
  calc_stage_r_2__instr_metadata__fe_exception_not_instr_,calc_stage_r_2__instr_metadata__fe_exception_code__1_,
  calc_stage_r_2__instr_metadata__fe_exception_code__0_,calc_stage_r_2__instr__31_,
  calc_stage_r_2__instr__30_,calc_stage_r_2__instr__29_,calc_stage_r_2__instr__28_,
  calc_stage_r_2__instr__27_,calc_stage_r_2__instr__26_,calc_stage_r_2__instr__25_,
  calc_stage_r_2__instr__24_,calc_stage_r_2__instr__23_,calc_stage_r_2__instr__22_,
  calc_stage_r_2__instr__21_,calc_stage_r_2__instr__20_,calc_stage_r_2__instr__19_,
  calc_stage_r_2__instr__18_,calc_stage_r_2__instr__17_,calc_stage_r_2__instr__16_,
  calc_stage_r_2__instr__15_,calc_stage_r_2__instr__14_,calc_stage_r_2__instr__13_,
  calc_stage_r_2__instr__12_,calc_stage_r_2__instr__11_,calc_stage_r_2__instr__10_,
  calc_stage_r_2__instr__9_,calc_stage_r_2__instr__8_,calc_stage_r_2__instr__7_,
  calc_stage_r_2__instr__6_,calc_stage_r_2__instr__5_,calc_stage_r_2__instr__4_,
  calc_stage_r_2__instr__3_,calc_stage_r_2__instr__2_,calc_stage_r_2__instr__1_,
  calc_stage_r_2__instr__0_,calc_stage_r_2__instr_v_,calc_stage_r_2__pipe_comp_v_,
  calc_stage_r_2__pipe_int_v_,calc_stage_r_2__pipe_mul_v_,calc_stage_r_2__pipe_mem_v_,
  calc_stage_r_2__pipe_fp_v_,calc_stage_r_2__irf_w_v_,calc_stage_r_2__frf_w_v_,
  calc_stage_r_1__instr_metadata__itag__7_,calc_stage_r_1__instr_metadata__itag__6_,
  calc_stage_r_1__instr_metadata__itag__5_,calc_stage_r_1__instr_metadata__itag__4_,
  calc_stage_r_1__instr_metadata__itag__3_,calc_stage_r_1__instr_metadata__itag__2_,
  calc_stage_r_1__instr_metadata__itag__1_,calc_stage_r_1__instr_metadata__itag__0_,
  calc_stage_r_1__instr_metadata__pc__63_,calc_stage_r_1__instr_metadata__pc__62_,
  calc_stage_r_1__instr_metadata__pc__61_,calc_stage_r_1__instr_metadata__pc__60_,
  calc_stage_r_1__instr_metadata__pc__59_,calc_stage_r_1__instr_metadata__pc__58_,
  calc_stage_r_1__instr_metadata__pc__57_,calc_stage_r_1__instr_metadata__pc__56_,
  calc_stage_r_1__instr_metadata__pc__55_,calc_stage_r_1__instr_metadata__pc__54_,
  calc_stage_r_1__instr_metadata__pc__53_,calc_stage_r_1__instr_metadata__pc__52_,
  calc_stage_r_1__instr_metadata__pc__51_,calc_stage_r_1__instr_metadata__pc__50_,
  calc_stage_r_1__instr_metadata__pc__49_,calc_stage_r_1__instr_metadata__pc__48_,
  calc_stage_r_1__instr_metadata__pc__47_,calc_stage_r_1__instr_metadata__pc__46_,
  calc_stage_r_1__instr_metadata__pc__45_,calc_stage_r_1__instr_metadata__pc__44_,
  calc_stage_r_1__instr_metadata__pc__43_,calc_stage_r_1__instr_metadata__pc__42_,
  calc_stage_r_1__instr_metadata__pc__41_,calc_stage_r_1__instr_metadata__pc__40_,
  calc_stage_r_1__instr_metadata__pc__39_,calc_stage_r_1__instr_metadata__pc__38_,
  calc_stage_r_1__instr_metadata__pc__37_,calc_stage_r_1__instr_metadata__pc__36_,
  calc_stage_r_1__instr_metadata__pc__35_,calc_stage_r_1__instr_metadata__pc__34_,
  calc_stage_r_1__instr_metadata__pc__33_,calc_stage_r_1__instr_metadata__pc__32_,
  calc_stage_r_1__instr_metadata__pc__31_,calc_stage_r_1__instr_metadata__pc__30_,
  calc_stage_r_1__instr_metadata__pc__29_,calc_stage_r_1__instr_metadata__pc__28_,
  calc_stage_r_1__instr_metadata__pc__27_,calc_stage_r_1__instr_metadata__pc__26_,
  calc_stage_r_1__instr_metadata__pc__25_,calc_stage_r_1__instr_metadata__pc__24_,
  calc_stage_r_1__instr_metadata__pc__23_,calc_stage_r_1__instr_metadata__pc__22_,
  calc_stage_r_1__instr_metadata__pc__21_,calc_stage_r_1__instr_metadata__pc__20_,
  calc_stage_r_1__instr_metadata__pc__19_,calc_stage_r_1__instr_metadata__pc__18_,
  calc_stage_r_1__instr_metadata__pc__17_,calc_stage_r_1__instr_metadata__pc__16_,
  calc_stage_r_1__instr_metadata__pc__15_,calc_stage_r_1__instr_metadata__pc__14_,
  calc_stage_r_1__instr_metadata__pc__13_,calc_stage_r_1__instr_metadata__pc__12_,
  calc_stage_r_1__instr_metadata__pc__11_,calc_stage_r_1__instr_metadata__pc__10_,
  calc_stage_r_1__instr_metadata__pc__9_,calc_stage_r_1__instr_metadata__pc__8_,
  calc_stage_r_1__instr_metadata__pc__7_,calc_stage_r_1__instr_metadata__pc__6_,
  calc_stage_r_1__instr_metadata__pc__5_,calc_stage_r_1__instr_metadata__pc__4_,
  calc_stage_r_1__instr_metadata__pc__3_,calc_stage_r_1__instr_metadata__pc__2_,
  calc_stage_r_1__instr_metadata__pc__1_,calc_stage_r_1__instr_metadata__pc__0_,
  calc_stage_r_1__instr_metadata__fe_exception_not_instr_,
  calc_stage_r_1__instr_metadata__fe_exception_code__1_,calc_stage_r_1__instr_metadata__fe_exception_code__0_,
  calc_stage_r_1__instr__31_,calc_stage_r_1__instr__30_,calc_stage_r_1__instr__29_,
  calc_stage_r_1__instr__28_,calc_stage_r_1__instr__27_,calc_stage_r_1__instr__26_,
  calc_stage_r_1__instr__25_,calc_stage_r_1__instr__24_,calc_stage_r_1__instr__23_,
  calc_stage_r_1__instr__22_,calc_stage_r_1__instr__21_,calc_stage_r_1__instr__20_,
  calc_stage_r_1__instr__19_,calc_stage_r_1__instr__18_,calc_stage_r_1__instr__17_,
  calc_stage_r_1__instr__16_,calc_stage_r_1__instr__15_,calc_stage_r_1__instr__14_,
  calc_stage_r_1__instr__13_,calc_stage_r_1__instr__12_,calc_stage_r_1__instr__11_,
  calc_stage_r_1__instr__10_,calc_stage_r_1__instr__9_,calc_stage_r_1__instr__8_,
  calc_stage_r_1__instr__7_,calc_stage_r_1__instr__6_,calc_stage_r_1__instr__5_,
  calc_stage_r_1__instr__4_,calc_stage_r_1__instr__3_,calc_stage_r_1__instr__2_,
  calc_stage_r_1__instr__1_,calc_stage_r_1__instr__0_,calc_stage_r_1__instr_v_,
  calc_stage_r_1__pipe_comp_v_,calc_stage_r_1__pipe_int_v_,calc_stage_r_1__pipe_mul_v_,
  calc_stage_r_1__pipe_mem_v_,calc_stage_r_1__pipe_fp_v_,calc_stage_r_1__irf_w_v_,
  calc_stage_r_1__frf_w_v_,calc_stage_r_0__instr_metadata__itag__7_,
  calc_stage_r_0__instr_metadata__itag__6_,calc_stage_r_0__instr_metadata__itag__5_,
  calc_stage_r_0__instr_metadata__itag__4_,calc_stage_r_0__instr_metadata__itag__3_,
  calc_stage_r_0__instr_metadata__itag__2_,calc_stage_r_0__instr_metadata__itag__1_,
  calc_stage_r_0__instr_metadata__itag__0_,calc_stage_r_0__instr_metadata__pc__63_,
  calc_stage_r_0__instr_metadata__pc__62_,calc_stage_r_0__instr_metadata__pc__61_,
  calc_stage_r_0__instr_metadata__pc__60_,calc_stage_r_0__instr_metadata__pc__59_,
  calc_stage_r_0__instr_metadata__pc__58_,calc_stage_r_0__instr_metadata__pc__57_,
  calc_stage_r_0__instr_metadata__pc__56_,calc_stage_r_0__instr_metadata__pc__55_,
  calc_stage_r_0__instr_metadata__pc__54_,calc_stage_r_0__instr_metadata__pc__53_,
  calc_stage_r_0__instr_metadata__pc__52_,calc_stage_r_0__instr_metadata__pc__51_,
  calc_stage_r_0__instr_metadata__pc__50_,calc_stage_r_0__instr_metadata__pc__49_,
  calc_stage_r_0__instr_metadata__pc__48_,calc_stage_r_0__instr_metadata__pc__47_,
  calc_stage_r_0__instr_metadata__pc__46_,calc_stage_r_0__instr_metadata__pc__45_,
  calc_stage_r_0__instr_metadata__pc__44_,calc_stage_r_0__instr_metadata__pc__43_,
  calc_stage_r_0__instr_metadata__pc__42_,calc_stage_r_0__instr_metadata__pc__41_,
  calc_stage_r_0__instr_metadata__pc__40_,calc_stage_r_0__instr_metadata__pc__39_,
  calc_stage_r_0__instr_metadata__pc__38_,calc_stage_r_0__instr_metadata__pc__37_,
  calc_stage_r_0__instr_metadata__pc__36_,calc_stage_r_0__instr_metadata__pc__35_,
  calc_stage_r_0__instr_metadata__pc__34_,calc_stage_r_0__instr_metadata__pc__33_,
  calc_stage_r_0__instr_metadata__pc__32_,calc_stage_r_0__instr_metadata__pc__31_,
  calc_stage_r_0__instr_metadata__pc__30_,calc_stage_r_0__instr_metadata__pc__29_,
  calc_stage_r_0__instr_metadata__pc__28_,calc_stage_r_0__instr_metadata__pc__27_,
  calc_stage_r_0__instr_metadata__pc__26_,calc_stage_r_0__instr_metadata__pc__25_,
  calc_stage_r_0__instr_metadata__pc__24_,calc_stage_r_0__instr_metadata__pc__23_,
  calc_stage_r_0__instr_metadata__pc__22_,calc_stage_r_0__instr_metadata__pc__21_,
  calc_stage_r_0__instr_metadata__pc__20_,calc_stage_r_0__instr_metadata__pc__19_,
  calc_stage_r_0__instr_metadata__pc__18_,calc_stage_r_0__instr_metadata__pc__17_,
  calc_stage_r_0__instr_metadata__pc__16_,calc_stage_r_0__instr_metadata__pc__15_,
  calc_stage_r_0__instr_metadata__pc__14_,calc_stage_r_0__instr_metadata__pc__13_,
  calc_stage_r_0__instr_metadata__pc__12_,calc_stage_r_0__instr_metadata__pc__11_,
  calc_stage_r_0__instr_metadata__pc__10_,calc_stage_r_0__instr_metadata__pc__9_,
  calc_stage_r_0__instr_metadata__pc__8_,calc_stage_r_0__instr_metadata__pc__7_,
  calc_stage_r_0__instr_metadata__pc__6_,calc_stage_r_0__instr_metadata__pc__5_,
  calc_stage_r_0__instr_metadata__pc__4_,calc_stage_r_0__instr_metadata__pc__3_,
  calc_stage_r_0__instr_metadata__pc__2_,calc_stage_r_0__instr_metadata__pc__1_,
  calc_stage_r_0__instr_metadata__pc__0_,calc_stage_r_0__instr_metadata__fe_exception_not_instr_,
  calc_stage_r_0__instr_metadata__fe_exception_code__1_,
  calc_stage_r_0__instr_metadata__fe_exception_code__0_,calc_stage_r_0__instr__31_,calc_stage_r_0__instr__30_,
  calc_stage_r_0__instr__29_,calc_stage_r_0__instr__28_,calc_stage_r_0__instr__27_,
  calc_stage_r_0__instr__26_,calc_stage_r_0__instr__25_,calc_stage_r_0__instr__24_,
  calc_stage_r_0__instr__23_,calc_stage_r_0__instr__22_,calc_stage_r_0__instr__21_,
  calc_stage_r_0__instr__20_,calc_stage_r_0__instr__19_,calc_stage_r_0__instr__18_,
  calc_stage_r_0__instr__17_,calc_stage_r_0__instr__16_,calc_stage_r_0__instr__15_,
  calc_stage_r_0__instr__14_,calc_stage_r_0__instr__13_,calc_stage_r_0__instr__12_,
  calc_stage_r_0__instr__11_,calc_stage_r_0__instr__10_,calc_stage_r_0__instr__9_,
  calc_stage_r_0__instr__8_,calc_stage_r_0__instr__7_,calc_stage_r_0__instr__6_,
  calc_stage_r_0__instr__5_,calc_stage_r_0__instr__4_,calc_stage_r_0__instr__3_,
  calc_stage_r_0__instr__2_,calc_stage_r_0__instr__1_,calc_stage_r_0__instr__0_,
  calc_stage_r_0__instr_v_,calc_stage_r_0__pipe_comp_v_,calc_stage_r_0__pipe_int_v_,
  calc_stage_r_0__pipe_mul_v_,calc_stage_r_0__pipe_mem_v_,calc_stage_r_0__pipe_fp_v_,
  calc_stage_r_0__irf_w_v_,calc_stage_r_0__frf_w_v_,exc_stage_r_4__poison_v_,
  exc_stage_r_4__roll_v_,exc_stage_r_4__illegal_instr_v_,exc_stage_r_4__ret_instr_v_,
  exc_stage_r_4__csr_instr_v_,exc_stage_r_4__tlb_miss_v_,exc_stage_r_4__load_fault_v_,
  exc_stage_r_4__store_fault_v_,exc_stage_r_4__cache_miss_v_,exc_stage_r_3__roll_v_,
  exc_stage_r_3__illegal_instr_v_,exc_stage_r_3__ret_instr_v_,
  exc_stage_r_3__csr_instr_v_,exc_stage_r_3__tlb_miss_v_,exc_stage_r_3__load_fault_v_,
  exc_stage_r_3__store_fault_v_,exc_stage_r_3__cache_miss_v_,exc_stage_r_2__poison_v_,
  exc_stage_r_2__roll_v_,exc_stage_r_2__illegal_instr_v_,exc_stage_r_2__ret_instr_v_,
  exc_stage_r_2__csr_instr_v_,exc_stage_r_2__tlb_miss_v_,exc_stage_r_2__load_fault_v_,
  exc_stage_r_2__store_fault_v_,exc_stage_r_2__cache_miss_v_,exc_stage_r_1__poison_v_,
  exc_stage_r_1__roll_v_,exc_stage_r_1__illegal_instr_v_,
  exc_stage_r_1__ret_instr_v_,exc_stage_r_1__csr_instr_v_,exc_stage_r_1__tlb_miss_v_,
  exc_stage_r_1__load_fault_v_,exc_stage_r_1__store_fault_v_,exc_stage_r_1__cache_miss_v_,
  exc_stage_r_0__poison_v_,exc_stage_r_0__roll_v_,exc_stage_r_0__illegal_instr_v_,
  exc_stage_r_0__ret_instr_v_,exc_stage_r_0__csr_instr_v_,exc_stage_r_0__tlb_miss_v_,
  exc_stage_r_0__load_fault_v_,exc_stage_r_0__store_fault_v_,exc_stage_r_0__cache_miss_v_,
  n_6_net_,n_12_net_,issue_pkt_r_instr_metadata__itag__7_,
  issue_pkt_r_instr_metadata__itag__6_,issue_pkt_r_instr_metadata__itag__5_,
  issue_pkt_r_instr_metadata__itag__4_,issue_pkt_r_instr_metadata__itag__3_,issue_pkt_r_instr_metadata__itag__2_,
  issue_pkt_r_instr_metadata__itag__1_,issue_pkt_r_instr_metadata__itag__0_,
  issue_pkt_r_instr_metadata__pc__63_,issue_pkt_r_instr_metadata__pc__62_,
  issue_pkt_r_instr_metadata__pc__61_,issue_pkt_r_instr_metadata__pc__60_,
  issue_pkt_r_instr_metadata__pc__59_,issue_pkt_r_instr_metadata__pc__58_,
  issue_pkt_r_instr_metadata__pc__57_,issue_pkt_r_instr_metadata__pc__56_,issue_pkt_r_instr_metadata__pc__55_,
  issue_pkt_r_instr_metadata__pc__54_,issue_pkt_r_instr_metadata__pc__53_,
  issue_pkt_r_instr_metadata__pc__52_,issue_pkt_r_instr_metadata__pc__51_,
  issue_pkt_r_instr_metadata__pc__50_,issue_pkt_r_instr_metadata__pc__49_,
  issue_pkt_r_instr_metadata__pc__48_,issue_pkt_r_instr_metadata__pc__47_,issue_pkt_r_instr_metadata__pc__46_,
  issue_pkt_r_instr_metadata__pc__45_,issue_pkt_r_instr_metadata__pc__44_,
  issue_pkt_r_instr_metadata__pc__43_,issue_pkt_r_instr_metadata__pc__42_,
  issue_pkt_r_instr_metadata__pc__41_,issue_pkt_r_instr_metadata__pc__40_,
  issue_pkt_r_instr_metadata__pc__39_,issue_pkt_r_instr_metadata__pc__38_,
  issue_pkt_r_instr_metadata__pc__37_,issue_pkt_r_instr_metadata__pc__36_,issue_pkt_r_instr_metadata__pc__35_,
  issue_pkt_r_instr_metadata__pc__34_,issue_pkt_r_instr_metadata__pc__33_,
  issue_pkt_r_instr_metadata__pc__32_,issue_pkt_r_instr_metadata__pc__31_,
  issue_pkt_r_instr_metadata__pc__30_,issue_pkt_r_instr_metadata__pc__29_,
  issue_pkt_r_instr_metadata__pc__28_,issue_pkt_r_instr_metadata__pc__27_,issue_pkt_r_instr_metadata__pc__26_,
  issue_pkt_r_instr_metadata__pc__25_,issue_pkt_r_instr_metadata__pc__24_,
  issue_pkt_r_instr_metadata__pc__23_,issue_pkt_r_instr_metadata__pc__22_,
  issue_pkt_r_instr_metadata__pc__21_,issue_pkt_r_instr_metadata__pc__20_,
  issue_pkt_r_instr_metadata__pc__19_,issue_pkt_r_instr_metadata__pc__18_,
  issue_pkt_r_instr_metadata__pc__17_,issue_pkt_r_instr_metadata__pc__16_,issue_pkt_r_instr_metadata__pc__15_,
  issue_pkt_r_instr_metadata__pc__14_,issue_pkt_r_instr_metadata__pc__13_,
  issue_pkt_r_instr_metadata__pc__12_,issue_pkt_r_instr_metadata__pc__11_,
  issue_pkt_r_instr_metadata__pc__10_,issue_pkt_r_instr_metadata__pc__9_,
  issue_pkt_r_instr_metadata__pc__8_,issue_pkt_r_instr_metadata__pc__7_,issue_pkt_r_instr_metadata__pc__6_,
  issue_pkt_r_instr_metadata__pc__5_,issue_pkt_r_instr_metadata__pc__4_,
  issue_pkt_r_instr_metadata__pc__3_,issue_pkt_r_instr_metadata__pc__2_,
  issue_pkt_r_instr_metadata__pc__1_,issue_pkt_r_instr_metadata__pc__0_,
  issue_pkt_r_instr_metadata__fe_exception_not_instr_,issue_pkt_r_instr_metadata__fe_exception_code__1_,
  issue_pkt_r_instr_metadata__fe_exception_code__0_,issue_pkt_r_branch_metadata_fwd__35_,
  issue_pkt_r_branch_metadata_fwd__34_,issue_pkt_r_branch_metadata_fwd__33_,
  issue_pkt_r_branch_metadata_fwd__32_,issue_pkt_r_branch_metadata_fwd__31_,
  issue_pkt_r_branch_metadata_fwd__30_,issue_pkt_r_branch_metadata_fwd__29_,
  issue_pkt_r_branch_metadata_fwd__28_,issue_pkt_r_branch_metadata_fwd__27_,
  issue_pkt_r_branch_metadata_fwd__26_,issue_pkt_r_branch_metadata_fwd__25_,
  issue_pkt_r_branch_metadata_fwd__24_,issue_pkt_r_branch_metadata_fwd__23_,issue_pkt_r_branch_metadata_fwd__22_,
  issue_pkt_r_branch_metadata_fwd__21_,issue_pkt_r_branch_metadata_fwd__20_,
  issue_pkt_r_branch_metadata_fwd__19_,issue_pkt_r_branch_metadata_fwd__18_,
  issue_pkt_r_branch_metadata_fwd__17_,issue_pkt_r_branch_metadata_fwd__16_,
  issue_pkt_r_branch_metadata_fwd__15_,issue_pkt_r_branch_metadata_fwd__14_,
  issue_pkt_r_branch_metadata_fwd__13_,issue_pkt_r_branch_metadata_fwd__12_,
  issue_pkt_r_branch_metadata_fwd__11_,issue_pkt_r_branch_metadata_fwd__10_,issue_pkt_r_branch_metadata_fwd__9_,
  issue_pkt_r_branch_metadata_fwd__8_,issue_pkt_r_branch_metadata_fwd__7_,
  issue_pkt_r_branch_metadata_fwd__6_,issue_pkt_r_branch_metadata_fwd__5_,
  issue_pkt_r_branch_metadata_fwd__4_,issue_pkt_r_branch_metadata_fwd__3_,
  issue_pkt_r_branch_metadata_fwd__2_,issue_pkt_r_branch_metadata_fwd__1_,issue_pkt_r_branch_metadata_fwd__0_,
  issue_pkt_r_instr__31_,issue_pkt_r_instr__30_,issue_pkt_r_instr__29_,
  issue_pkt_r_instr__28_,issue_pkt_r_instr__27_,issue_pkt_r_instr__26_,issue_pkt_r_instr__25_,
  issue_pkt_r_instr__24_,issue_pkt_r_instr__23_,issue_pkt_r_instr__22_,
  issue_pkt_r_instr__21_,issue_pkt_r_instr__20_,issue_pkt_r_instr__19_,
  issue_pkt_r_instr__18_,issue_pkt_r_instr__17_,issue_pkt_r_instr__16_,issue_pkt_r_instr__15_,
  issue_pkt_r_instr__14_,issue_pkt_r_instr__13_,issue_pkt_r_instr__12_,
  issue_pkt_r_instr__11_,issue_pkt_r_instr__10_,issue_pkt_r_instr__9_,issue_pkt_r_instr__8_,
  issue_pkt_r_instr__7_,issue_pkt_r_instr__6_,issue_pkt_r_instr__5_,issue_pkt_r_instr__4_,
  issue_pkt_r_instr__3_,issue_pkt_r_instr__2_,issue_pkt_r_instr__1_,
  issue_pkt_r_instr__0_,issue_pkt_r_imm__63_,issue_pkt_r_imm__62_,issue_pkt_r_imm__61_,
  issue_pkt_r_imm__60_,issue_pkt_r_imm__59_,issue_pkt_r_imm__58_,issue_pkt_r_imm__57_,
  issue_pkt_r_imm__56_,issue_pkt_r_imm__55_,issue_pkt_r_imm__54_,issue_pkt_r_imm__53_,
  issue_pkt_r_imm__52_,issue_pkt_r_imm__51_,issue_pkt_r_imm__50_,issue_pkt_r_imm__49_,
  issue_pkt_r_imm__48_,issue_pkt_r_imm__47_,issue_pkt_r_imm__46_,
  issue_pkt_r_imm__45_,issue_pkt_r_imm__44_,issue_pkt_r_imm__43_,issue_pkt_r_imm__42_,
  issue_pkt_r_imm__41_,issue_pkt_r_imm__40_,issue_pkt_r_imm__39_,issue_pkt_r_imm__38_,
  issue_pkt_r_imm__37_,issue_pkt_r_imm__36_,issue_pkt_r_imm__35_,issue_pkt_r_imm__34_,
  issue_pkt_r_imm__33_,issue_pkt_r_imm__32_,issue_pkt_r_imm__31_,issue_pkt_r_imm__30_,
  issue_pkt_r_imm__29_,issue_pkt_r_imm__28_,issue_pkt_r_imm__27_,
  issue_pkt_r_imm__26_,issue_pkt_r_imm__25_,issue_pkt_r_imm__24_,issue_pkt_r_imm__23_,
  issue_pkt_r_imm__22_,issue_pkt_r_imm__21_,issue_pkt_r_imm__20_,issue_pkt_r_imm__19_,
  issue_pkt_r_imm__18_,issue_pkt_r_imm__17_,issue_pkt_r_imm__16_,issue_pkt_r_imm__15_,
  issue_pkt_r_imm__14_,issue_pkt_r_imm__13_,issue_pkt_r_imm__12_,issue_pkt_r_imm__11_,
  issue_pkt_r_imm__10_,issue_pkt_r_imm__9_,issue_pkt_r_imm__8_,issue_pkt_r_imm__7_,
  issue_pkt_r_imm__6_,issue_pkt_r_imm__5_,issue_pkt_r_imm__4_,issue_pkt_r_imm__3_,
  issue_pkt_r_imm__2_,issue_pkt_r_imm__1_,issue_pkt_r_imm__0_,illegal_instr_isd,
  n_28_net_,dispatch_pkt_r_instr_metadata__itag__7_,
  dispatch_pkt_r_instr_metadata__itag__6_,dispatch_pkt_r_instr_metadata__itag__5_,
  dispatch_pkt_r_instr_metadata__itag__4_,dispatch_pkt_r_instr_metadata__itag__3_,
  dispatch_pkt_r_instr_metadata__itag__2_,dispatch_pkt_r_instr_metadata__itag__1_,
  dispatch_pkt_r_instr_metadata__itag__0_,dispatch_pkt_r_instr_metadata__fe_exception_not_instr_,
  dispatch_pkt_r_instr_metadata__fe_exception_code__1_,
  dispatch_pkt_r_instr_metadata__fe_exception_code__0_,dispatch_pkt_r_instr__31_,dispatch_pkt_r_instr__30_,
  dispatch_pkt_r_instr__29_,dispatch_pkt_r_instr__28_,dispatch_pkt_r_instr__27_,
  dispatch_pkt_r_instr__26_,dispatch_pkt_r_instr__25_,dispatch_pkt_r_instr__24_,
  dispatch_pkt_r_instr__23_,dispatch_pkt_r_instr__22_,dispatch_pkt_r_instr__21_,dispatch_pkt_r_instr__20_,
  dispatch_pkt_r_instr__19_,dispatch_pkt_r_instr__18_,dispatch_pkt_r_instr__17_,
  dispatch_pkt_r_instr__16_,dispatch_pkt_r_instr__15_,dispatch_pkt_r_instr__14_,
  dispatch_pkt_r_instr__13_,dispatch_pkt_r_instr__12_,dispatch_pkt_r_instr__11_,
  dispatch_pkt_r_instr__10_,dispatch_pkt_r_instr__9_,dispatch_pkt_r_instr__8_,
  dispatch_pkt_r_instr__7_,dispatch_pkt_r_instr__6_,dispatch_pkt_r_instr__5_,
  dispatch_pkt_r_instr__4_,dispatch_pkt_r_instr__3_,dispatch_pkt_r_instr__2_,
  dispatch_pkt_r_instr__1_,dispatch_pkt_r_instr__0_,dispatch_pkt_r_decode__fe_nop_v_,
  dispatch_pkt_r_decode__be_nop_v_,dispatch_pkt_r_decode__me_nop_v_,
  dispatch_pkt_r_decode__pipe_comp_v_,dispatch_pkt_r_decode__pipe_mul_v_,dispatch_pkt_r_decode__pipe_mem_v_,
  dispatch_pkt_r_decode__pipe_fp_v_,dispatch_pkt_r_decode__irf_w_v_,
  dispatch_pkt_r_decode__frf_w_v_,dispatch_pkt_r_decode__csr_instr_v_,
  dispatch_pkt_r_decode__mhartid_r_v_,dispatch_pkt_r_decode__mcycle_r_v_,dispatch_pkt_r_decode__mtime_r_v_,
  dispatch_pkt_r_decode__minstret_r_v_,dispatch_pkt_r_decode__mtvec_rw_v_,
  dispatch_pkt_r_decode__mtval_rw_v_,dispatch_pkt_r_decode__mepc_rw_v_,
  dispatch_pkt_r_decode__mscratch_rw_v_,dispatch_pkt_r_decode__dcache_w_v_,
  dispatch_pkt_r_decode__dcache_r_v_,dispatch_pkt_r_decode__fp_not_int_v_,dispatch_pkt_r_decode__ret_v_,
  dispatch_pkt_r_decode__amo_v_,dispatch_pkt_r_decode__jmp_v_,dispatch_pkt_r_decode__br_v_,
  dispatch_pkt_r_decode__opw_v_,dispatch_pkt_r_decode__fu_op__fu_op__3_,
  dispatch_pkt_r_decode__fu_op__fu_op__2_,dispatch_pkt_r_decode__fu_op__fu_op__1_,
  dispatch_pkt_r_decode__fu_op__fu_op__0_,dispatch_pkt_r_decode__rs1_addr__4_,
  dispatch_pkt_r_decode__rs1_addr__3_,dispatch_pkt_r_decode__rs1_addr__2_,
  dispatch_pkt_r_decode__rs1_addr__1_,dispatch_pkt_r_decode__rs1_addr__0_,
  dispatch_pkt_r_decode__rs2_addr__4_,dispatch_pkt_r_decode__rs2_addr__3_,dispatch_pkt_r_decode__rs2_addr__2_,
  dispatch_pkt_r_decode__rs2_addr__1_,dispatch_pkt_r_decode__rs2_addr__0_,
  dispatch_pkt_r_decode__rd_addr__4_,dispatch_pkt_r_decode__rd_addr__3_,
  dispatch_pkt_r_decode__rd_addr__2_,dispatch_pkt_r_decode__rd_addr__1_,
  dispatch_pkt_r_decode__rd_addr__0_,dispatch_pkt_r_decode__src1_sel_,dispatch_pkt_r_decode__src2_sel_,
  dispatch_pkt_r_decode__baddr_sel_,dispatch_pkt_r_decode__result_sel_,
  dispatch_pkt_r_rs1__63_,dispatch_pkt_r_rs1__62_,dispatch_pkt_r_rs1__61_,dispatch_pkt_r_rs1__60_,
  dispatch_pkt_r_rs1__59_,dispatch_pkt_r_rs1__58_,dispatch_pkt_r_rs1__57_,
  dispatch_pkt_r_rs1__56_,dispatch_pkt_r_rs1__55_,dispatch_pkt_r_rs1__54_,
  dispatch_pkt_r_rs1__53_,dispatch_pkt_r_rs1__52_,dispatch_pkt_r_rs1__51_,dispatch_pkt_r_rs1__50_,
  dispatch_pkt_r_rs1__49_,dispatch_pkt_r_rs1__48_,dispatch_pkt_r_rs1__47_,
  dispatch_pkt_r_rs1__46_,dispatch_pkt_r_rs1__45_,dispatch_pkt_r_rs1__44_,
  dispatch_pkt_r_rs1__43_,dispatch_pkt_r_rs1__42_,dispatch_pkt_r_rs1__41_,dispatch_pkt_r_rs1__40_,
  dispatch_pkt_r_rs1__39_,dispatch_pkt_r_rs1__38_,dispatch_pkt_r_rs1__37_,
  dispatch_pkt_r_rs1__36_,dispatch_pkt_r_rs1__35_,dispatch_pkt_r_rs1__34_,
  dispatch_pkt_r_rs1__33_,dispatch_pkt_r_rs1__32_,dispatch_pkt_r_rs1__31_,dispatch_pkt_r_rs1__30_,
  dispatch_pkt_r_rs1__29_,dispatch_pkt_r_rs1__28_,dispatch_pkt_r_rs1__27_,
  dispatch_pkt_r_rs1__26_,dispatch_pkt_r_rs1__25_,dispatch_pkt_r_rs1__24_,
  dispatch_pkt_r_rs1__23_,dispatch_pkt_r_rs1__22_,dispatch_pkt_r_rs1__21_,dispatch_pkt_r_rs1__20_,
  dispatch_pkt_r_rs1__19_,dispatch_pkt_r_rs1__18_,dispatch_pkt_r_rs1__17_,
  dispatch_pkt_r_rs1__16_,dispatch_pkt_r_rs1__15_,dispatch_pkt_r_rs1__14_,
  dispatch_pkt_r_rs1__13_,dispatch_pkt_r_rs1__12_,dispatch_pkt_r_rs1__11_,dispatch_pkt_r_rs1__10_,
  dispatch_pkt_r_rs1__9_,dispatch_pkt_r_rs1__8_,dispatch_pkt_r_rs1__7_,
  dispatch_pkt_r_rs1__6_,dispatch_pkt_r_rs1__5_,dispatch_pkt_r_rs1__4_,dispatch_pkt_r_rs1__3_,
  dispatch_pkt_r_rs1__2_,dispatch_pkt_r_rs1__1_,dispatch_pkt_r_rs1__0_,
  dispatch_pkt_r_rs2__63_,dispatch_pkt_r_rs2__62_,dispatch_pkt_r_rs2__61_,
  dispatch_pkt_r_rs2__60_,dispatch_pkt_r_rs2__59_,dispatch_pkt_r_rs2__58_,dispatch_pkt_r_rs2__57_,
  dispatch_pkt_r_rs2__56_,dispatch_pkt_r_rs2__55_,dispatch_pkt_r_rs2__54_,
  dispatch_pkt_r_rs2__53_,dispatch_pkt_r_rs2__52_,dispatch_pkt_r_rs2__51_,
  dispatch_pkt_r_rs2__50_,dispatch_pkt_r_rs2__49_,dispatch_pkt_r_rs2__48_,dispatch_pkt_r_rs2__47_,
  dispatch_pkt_r_rs2__46_,dispatch_pkt_r_rs2__45_,dispatch_pkt_r_rs2__44_,
  dispatch_pkt_r_rs2__43_,dispatch_pkt_r_rs2__42_,dispatch_pkt_r_rs2__41_,
  dispatch_pkt_r_rs2__40_,dispatch_pkt_r_rs2__39_,dispatch_pkt_r_rs2__38_,dispatch_pkt_r_rs2__37_,
  dispatch_pkt_r_rs2__36_,dispatch_pkt_r_rs2__35_,dispatch_pkt_r_rs2__34_,
  dispatch_pkt_r_rs2__33_,dispatch_pkt_r_rs2__32_,dispatch_pkt_r_rs2__31_,
  dispatch_pkt_r_rs2__30_,dispatch_pkt_r_rs2__29_,dispatch_pkt_r_rs2__28_,dispatch_pkt_r_rs2__27_,
  dispatch_pkt_r_rs2__26_,dispatch_pkt_r_rs2__25_,dispatch_pkt_r_rs2__24_,
  dispatch_pkt_r_rs2__23_,dispatch_pkt_r_rs2__22_,dispatch_pkt_r_rs2__21_,
  dispatch_pkt_r_rs2__20_,dispatch_pkt_r_rs2__19_,dispatch_pkt_r_rs2__18_,dispatch_pkt_r_rs2__17_,
  dispatch_pkt_r_rs2__16_,dispatch_pkt_r_rs2__15_,dispatch_pkt_r_rs2__14_,
  dispatch_pkt_r_rs2__13_,dispatch_pkt_r_rs2__12_,dispatch_pkt_r_rs2__11_,
  dispatch_pkt_r_rs2__10_,dispatch_pkt_r_rs2__9_,dispatch_pkt_r_rs2__8_,dispatch_pkt_r_rs2__7_,
  dispatch_pkt_r_rs2__6_,dispatch_pkt_r_rs2__5_,dispatch_pkt_r_rs2__4_,
  dispatch_pkt_r_rs2__3_,dispatch_pkt_r_rs2__2_,dispatch_pkt_r_rs2__1_,dispatch_pkt_r_rs2__0_,
  dispatch_pkt_r_imm__63_,dispatch_pkt_r_imm__62_,dispatch_pkt_r_imm__61_,
  dispatch_pkt_r_imm__60_,dispatch_pkt_r_imm__59_,dispatch_pkt_r_imm__58_,dispatch_pkt_r_imm__57_,
  dispatch_pkt_r_imm__56_,dispatch_pkt_r_imm__55_,dispatch_pkt_r_imm__54_,
  dispatch_pkt_r_imm__53_,dispatch_pkt_r_imm__52_,dispatch_pkt_r_imm__51_,
  dispatch_pkt_r_imm__50_,dispatch_pkt_r_imm__49_,dispatch_pkt_r_imm__48_,dispatch_pkt_r_imm__47_,
  dispatch_pkt_r_imm__46_,dispatch_pkt_r_imm__45_,dispatch_pkt_r_imm__44_,
  dispatch_pkt_r_imm__43_,dispatch_pkt_r_imm__42_,dispatch_pkt_r_imm__41_,
  dispatch_pkt_r_imm__40_,dispatch_pkt_r_imm__39_,dispatch_pkt_r_imm__38_,dispatch_pkt_r_imm__37_,
  dispatch_pkt_r_imm__36_,dispatch_pkt_r_imm__35_,dispatch_pkt_r_imm__34_,
  dispatch_pkt_r_imm__33_,dispatch_pkt_r_imm__32_,dispatch_pkt_r_imm__31_,
  dispatch_pkt_r_imm__30_,dispatch_pkt_r_imm__29_,dispatch_pkt_r_imm__28_,dispatch_pkt_r_imm__27_,
  dispatch_pkt_r_imm__26_,dispatch_pkt_r_imm__25_,dispatch_pkt_r_imm__24_,
  dispatch_pkt_r_imm__23_,dispatch_pkt_r_imm__22_,dispatch_pkt_r_imm__21_,
  dispatch_pkt_r_imm__20_,dispatch_pkt_r_imm__19_,dispatch_pkt_r_imm__18_,dispatch_pkt_r_imm__17_,
  dispatch_pkt_r_imm__16_,dispatch_pkt_r_imm__15_,dispatch_pkt_r_imm__14_,
  dispatch_pkt_r_imm__13_,dispatch_pkt_r_imm__12_,dispatch_pkt_r_imm__11_,
  dispatch_pkt_r_imm__10_,dispatch_pkt_r_imm__9_,dispatch_pkt_r_imm__8_,dispatch_pkt_r_imm__7_,
  dispatch_pkt_r_imm__6_,dispatch_pkt_r_imm__5_,dispatch_pkt_r_imm__4_,
  dispatch_pkt_r_imm__3_,dispatch_pkt_r_imm__2_,dispatch_pkt_r_imm__1_,dispatch_pkt_r_imm__0_,
  exc_stage_n_4__poison_v_,exc_stage_n_3__poison_v_,exc_stage_n_3__roll_v_,
  exc_stage_n_3__cache_miss_v_,exc_stage_n_2__poison_v_,exc_stage_n_2__roll_v_,
  exc_stage_n_1__poison_v_,exc_stage_n_1__roll_v_,exc_stage_n_0__illegal_instr_v_,
  exc_stage_n_0__ret_instr_v_,exc_stage_n_0__csr_instr_v_,mtval_w_v_lo,mscratch_w_v_lo,
  fe_nop_v,be_nop_v,me_nop_v,n_63_net_,n_64_net_,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,
  N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,
  N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,
  N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,
  N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,
  N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,
  N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,
  N129,N130,N131,N132,N133,N134,N135,N136,N137,N138;
  wire [319:0] comp_stage_r,comp_stage_n;
  wire [50:0] decoded;
  wire [4:1] comp_stage_n_slice_iwb_v,comp_stage_n_slice_fwb_v;
  wire [385:0] dispatch_pkt;
  assign cmt_data_o[0] = 1'b0;
  assign cmt_data_o[1] = 1'b0;
  assign cmt_data_o[2] = 1'b0;
  assign cmt_data_o[3] = 1'b0;
  assign cmt_data_o[4] = 1'b0;
  assign cmt_data_o[5] = 1'b0;
  assign cmt_data_o[6] = 1'b0;
  assign cmt_data_o[7] = 1'b0;
  assign cmt_data_o[8] = 1'b0;
  assign cmt_data_o[9] = 1'b0;
  assign cmt_data_o[10] = 1'b0;
  assign cmt_data_o[11] = 1'b0;
  assign cmt_data_o[12] = 1'b0;
  assign cmt_data_o[13] = 1'b0;
  assign cmt_data_o[14] = 1'b0;
  assign cmt_data_o[15] = 1'b0;
  assign cmt_data_o[16] = 1'b0;
  assign cmt_data_o[17] = 1'b0;
  assign cmt_data_o[18] = 1'b0;
  assign cmt_data_o[19] = 1'b0;
  assign cmt_data_o[20] = 1'b0;
  assign cmt_data_o[21] = 1'b0;
  assign cmt_data_o[22] = 1'b0;
  assign cmt_data_o[23] = 1'b0;
  assign cmt_data_o[24] = 1'b0;
  assign cmt_data_o[25] = 1'b0;
  assign cmt_data_o[26] = 1'b0;
  assign cmt_data_o[27] = 1'b0;
  assign cmt_data_o[28] = 1'b0;
  assign cmt_data_o[29] = 1'b0;
  assign cmt_data_o[30] = 1'b0;
  assign cmt_data_o[31] = 1'b0;
  assign cmt_data_o[32] = 1'b0;
  assign cmt_data_o[33] = 1'b0;
  assign cmt_data_o[34] = 1'b0;
  assign cmt_data_o[35] = 1'b0;
  assign cmt_data_o[36] = 1'b0;
  assign cmt_data_o[37] = 1'b0;
  assign cmt_data_o[38] = 1'b0;
  assign cmt_data_o[39] = 1'b0;
  assign cmt_data_o[40] = 1'b0;
  assign cmt_data_o[41] = 1'b0;
  assign cmt_data_o[42] = 1'b0;
  assign cmt_data_o[43] = 1'b0;
  assign cmt_data_o[44] = 1'b0;
  assign cmt_data_o[45] = 1'b0;
  assign cmt_data_o[46] = 1'b0;
  assign cmt_data_o[47] = 1'b0;
  assign cmt_data_o[48] = 1'b0;
  assign cmt_data_o[49] = 1'b0;
  assign cmt_data_o[50] = 1'b0;
  assign cmt_data_o[51] = 1'b0;
  assign cmt_data_o[52] = 1'b0;
  assign cmt_data_o[53] = 1'b0;
  assign cmt_data_o[54] = 1'b0;
  assign cmt_data_o[55] = 1'b0;
  assign cmt_data_o[56] = 1'b0;
  assign cmt_data_o[57] = 1'b0;
  assign cmt_data_o[58] = 1'b0;
  assign cmt_data_o[59] = 1'b0;
  assign cmt_data_o[60] = 1'b0;
  assign cmt_data_o[61] = 1'b0;
  assign cmt_data_o[62] = 1'b0;
  assign cmt_data_o[63] = 1'b0;
  assign cmt_mem_op_o[0] = 1'b0;
  assign cmt_mem_op_o[1] = 1'b0;
  assign cmt_mem_op_o[2] = 1'b0;
  assign cmt_mem_op_o[3] = 1'b0;
  assign cmt_mem_addr_o[0] = 1'b0;
  assign cmt_mem_addr_o[1] = 1'b0;
  assign cmt_mem_addr_o[2] = 1'b0;
  assign cmt_mem_addr_o[3] = 1'b0;
  assign cmt_mem_addr_o[4] = 1'b0;
  assign cmt_mem_addr_o[5] = 1'b0;
  assign cmt_mem_addr_o[6] = 1'b0;
  assign cmt_mem_addr_o[7] = 1'b0;
  assign cmt_mem_addr_o[8] = 1'b0;
  assign cmt_mem_addr_o[9] = 1'b0;
  assign cmt_mem_addr_o[10] = 1'b0;
  assign cmt_mem_addr_o[11] = 1'b0;
  assign cmt_mem_addr_o[12] = 1'b0;
  assign cmt_mem_addr_o[13] = 1'b0;
  assign cmt_mem_addr_o[14] = 1'b0;
  assign cmt_mem_addr_o[15] = 1'b0;
  assign cmt_mem_addr_o[16] = 1'b0;
  assign cmt_mem_addr_o[17] = 1'b0;
  assign cmt_mem_addr_o[18] = 1'b0;
  assign cmt_mem_addr_o[19] = 1'b0;
  assign cmt_mem_addr_o[20] = 1'b0;
  assign cmt_mem_addr_o[21] = 1'b0;
  assign cmt_mem_addr_o[22] = 1'b0;
  assign cmt_mem_addr_o[23] = 1'b0;
  assign cmt_mem_addr_o[24] = 1'b0;
  assign cmt_mem_addr_o[25] = 1'b0;
  assign cmt_mem_addr_o[26] = 1'b0;
  assign cmt_mem_addr_o[27] = 1'b0;
  assign cmt_mem_addr_o[28] = 1'b0;
  assign cmt_mem_addr_o[29] = 1'b0;
  assign cmt_mem_addr_o[30] = 1'b0;
  assign cmt_mem_addr_o[31] = 1'b0;
  assign cmt_mem_addr_o[32] = 1'b0;
  assign cmt_mem_addr_o[33] = 1'b0;
  assign cmt_mem_addr_o[34] = 1'b0;
  assign cmt_mem_addr_o[35] = 1'b0;
  assign cmt_mem_addr_o[36] = 1'b0;
  assign cmt_mem_addr_o[37] = 1'b0;
  assign cmt_mem_addr_o[38] = 1'b0;
  assign cmt_mem_addr_o[39] = 1'b0;
  assign cmt_mem_addr_o[40] = 1'b0;
  assign cmt_mem_addr_o[41] = 1'b0;
  assign cmt_mem_addr_o[42] = 1'b0;
  assign cmt_mem_addr_o[43] = 1'b0;
  assign cmt_mem_addr_o[44] = 1'b0;
  assign cmt_mem_addr_o[45] = 1'b0;
  assign cmt_mem_addr_o[46] = 1'b0;
  assign cmt_mem_addr_o[47] = 1'b0;
  assign cmt_mem_addr_o[48] = 1'b0;
  assign cmt_mem_addr_o[49] = 1'b0;
  assign cmt_mem_addr_o[50] = 1'b0;
  assign cmt_mem_addr_o[51] = 1'b0;
  assign cmt_mem_addr_o[52] = 1'b0;
  assign cmt_mem_addr_o[53] = 1'b0;
  assign cmt_mem_addr_o[54] = 1'b0;
  assign cmt_mem_addr_o[55] = 1'b0;
  assign cmt_mem_addr_o[56] = 1'b0;
  assign cmt_mem_addr_o[57] = 1'b0;
  assign cmt_mem_addr_o[58] = 1'b0;
  assign cmt_mem_addr_o[59] = 1'b0;
  assign cmt_mem_addr_o[60] = 1'b0;
  assign cmt_mem_addr_o[61] = 1'b0;
  assign cmt_mem_addr_o[62] = 1'b0;
  assign cmt_mem_addr_o[63] = 1'b0;
  assign cmt_mem_w_v_o = 1'b0;
  assign cmt_rd_addr_o[0] = 1'b0;
  assign cmt_rd_addr_o[1] = 1'b0;
  assign cmt_rd_addr_o[2] = 1'b0;
  assign cmt_rd_addr_o[3] = 1'b0;
  assign cmt_rd_addr_o[4] = 1'b0;
  assign cmt_rd_w_v_o = 1'b0;

  bp_be_regfile
  int_regfile
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .issue_v_i(issue_pkt_v_i),
    .dispatch_v_i(chk_dispatch_v_i),
    .rd_w_v_i(n_0_net_),
    .rd_addr_i(calc_status_o[106:102]),
    .rd_data_i(comp_stage_r[255:192]),
    .rs1_r_v_i(issue_pkt_i[77]),
    .rs1_addr_i(issue_pkt_i[73:69]),
    .rs1_data_o(irf_rs1),
    .rs2_r_v_i(issue_pkt_i[76]),
    .rs2_addr_i(issue_pkt_i[68:64]),
    .rs2_data_o(irf_rs2)
  );


  bp_be_regfile_harden_p0
  float_regfile
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .issue_v_i(issue_pkt_v_i),
    .dispatch_v_i(chk_dispatch_v_i),
    .rd_w_v_i(n_6_net_),
    .rd_addr_i(calc_status_o[117:113]),
    .rd_data_i(comp_stage_r[319:256]),
    .rs1_r_v_i(issue_pkt_i[75]),
    .rs1_addr_i(issue_pkt_i[73:69]),
    .rs1_data_o(frf_rs1),
    .rs2_r_v_i(issue_pkt_i[74]),
    .rs2_addr_i(issue_pkt_i[68:64]),
    .rs2_data_o(frf_rs2)
  );


  bsg_dff_reset_en_width_p222
  issue_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(n_12_net_),
    .data_i({ issue_pkt_v_i, issue_pkt_i }),
    .data_o({ calc_status_o[306:306], issue_pkt_r_instr_metadata__itag__7_, issue_pkt_r_instr_metadata__itag__6_, issue_pkt_r_instr_metadata__itag__5_, issue_pkt_r_instr_metadata__itag__4_, issue_pkt_r_instr_metadata__itag__3_, issue_pkt_r_instr_metadata__itag__2_, issue_pkt_r_instr_metadata__itag__1_, issue_pkt_r_instr_metadata__itag__0_, issue_pkt_r_instr_metadata__pc__63_, issue_pkt_r_instr_metadata__pc__62_, issue_pkt_r_instr_metadata__pc__61_, issue_pkt_r_instr_metadata__pc__60_, issue_pkt_r_instr_metadata__pc__59_, issue_pkt_r_instr_metadata__pc__58_, issue_pkt_r_instr_metadata__pc__57_, issue_pkt_r_instr_metadata__pc__56_, issue_pkt_r_instr_metadata__pc__55_, issue_pkt_r_instr_metadata__pc__54_, issue_pkt_r_instr_metadata__pc__53_, issue_pkt_r_instr_metadata__pc__52_, issue_pkt_r_instr_metadata__pc__51_, issue_pkt_r_instr_metadata__pc__50_, issue_pkt_r_instr_metadata__pc__49_, issue_pkt_r_instr_metadata__pc__48_, issue_pkt_r_instr_metadata__pc__47_, issue_pkt_r_instr_metadata__pc__46_, issue_pkt_r_instr_metadata__pc__45_, issue_pkt_r_instr_metadata__pc__44_, issue_pkt_r_instr_metadata__pc__43_, issue_pkt_r_instr_metadata__pc__42_, issue_pkt_r_instr_metadata__pc__41_, issue_pkt_r_instr_metadata__pc__40_, issue_pkt_r_instr_metadata__pc__39_, issue_pkt_r_instr_metadata__pc__38_, issue_pkt_r_instr_metadata__pc__37_, issue_pkt_r_instr_metadata__pc__36_, issue_pkt_r_instr_metadata__pc__35_, issue_pkt_r_instr_metadata__pc__34_, issue_pkt_r_instr_metadata__pc__33_, issue_pkt_r_instr_metadata__pc__32_, issue_pkt_r_instr_metadata__pc__31_, issue_pkt_r_instr_metadata__pc__30_, issue_pkt_r_instr_metadata__pc__29_, issue_pkt_r_instr_metadata__pc__28_, issue_pkt_r_instr_metadata__pc__27_, issue_pkt_r_instr_metadata__pc__26_, issue_pkt_r_instr_metadata__pc__25_, issue_pkt_r_instr_metadata__pc__24_, issue_pkt_r_instr_metadata__pc__23_, issue_pkt_r_instr_metadata__pc__22_, issue_pkt_r_instr_metadata__pc__21_, issue_pkt_r_instr_metadata__pc__20_, issue_pkt_r_instr_metadata__pc__19_, issue_pkt_r_instr_metadata__pc__18_, issue_pkt_r_instr_metadata__pc__17_, issue_pkt_r_instr_metadata__pc__16_, issue_pkt_r_instr_metadata__pc__15_, issue_pkt_r_instr_metadata__pc__14_, issue_pkt_r_instr_metadata__pc__13_, issue_pkt_r_instr_metadata__pc__12_, issue_pkt_r_instr_metadata__pc__11_, issue_pkt_r_instr_metadata__pc__10_, issue_pkt_r_instr_metadata__pc__9_, issue_pkt_r_instr_metadata__pc__8_, issue_pkt_r_instr_metadata__pc__7_, issue_pkt_r_instr_metadata__pc__6_, issue_pkt_r_instr_metadata__pc__5_, issue_pkt_r_instr_metadata__pc__4_, issue_pkt_r_instr_metadata__pc__3_, issue_pkt_r_instr_metadata__pc__2_, issue_pkt_r_instr_metadata__pc__1_, issue_pkt_r_instr_metadata__pc__0_, issue_pkt_r_instr_metadata__fe_exception_not_instr_, issue_pkt_r_instr_metadata__fe_exception_code__1_, issue_pkt_r_instr_metadata__fe_exception_code__0_, issue_pkt_r_branch_metadata_fwd__35_, issue_pkt_r_branch_metadata_fwd__34_, issue_pkt_r_branch_metadata_fwd__33_, issue_pkt_r_branch_metadata_fwd__32_, issue_pkt_r_branch_metadata_fwd__31_, issue_pkt_r_branch_metadata_fwd__30_, issue_pkt_r_branch_metadata_fwd__29_, issue_pkt_r_branch_metadata_fwd__28_, issue_pkt_r_branch_metadata_fwd__27_, issue_pkt_r_branch_metadata_fwd__26_, issue_pkt_r_branch_metadata_fwd__25_, issue_pkt_r_branch_metadata_fwd__24_, issue_pkt_r_branch_metadata_fwd__23_, issue_pkt_r_branch_metadata_fwd__22_, issue_pkt_r_branch_metadata_fwd__21_, issue_pkt_r_branch_metadata_fwd__20_, issue_pkt_r_branch_metadata_fwd__19_, issue_pkt_r_branch_metadata_fwd__18_, issue_pkt_r_branch_metadata_fwd__17_, issue_pkt_r_branch_metadata_fwd__16_, issue_pkt_r_branch_metadata_fwd__15_, issue_pkt_r_branch_metadata_fwd__14_, issue_pkt_r_branch_metadata_fwd__13_, issue_pkt_r_branch_metadata_fwd__12_, issue_pkt_r_branch_metadata_fwd__11_, issue_pkt_r_branch_metadata_fwd__10_, issue_pkt_r_branch_metadata_fwd__9_, issue_pkt_r_branch_metadata_fwd__8_, issue_pkt_r_branch_metadata_fwd__7_, issue_pkt_r_branch_metadata_fwd__6_, issue_pkt_r_branch_metadata_fwd__5_, issue_pkt_r_branch_metadata_fwd__4_, issue_pkt_r_branch_metadata_fwd__3_, issue_pkt_r_branch_metadata_fwd__2_, issue_pkt_r_branch_metadata_fwd__1_, issue_pkt_r_branch_metadata_fwd__0_, issue_pkt_r_instr__31_, issue_pkt_r_instr__30_, issue_pkt_r_instr__29_, issue_pkt_r_instr__28_, issue_pkt_r_instr__27_, issue_pkt_r_instr__26_, issue_pkt_r_instr__25_, issue_pkt_r_instr__24_, issue_pkt_r_instr__23_, issue_pkt_r_instr__22_, issue_pkt_r_instr__21_, issue_pkt_r_instr__20_, issue_pkt_r_instr__19_, issue_pkt_r_instr__18_, issue_pkt_r_instr__17_, issue_pkt_r_instr__16_, issue_pkt_r_instr__15_, issue_pkt_r_instr__14_, issue_pkt_r_instr__13_, issue_pkt_r_instr__12_, issue_pkt_r_instr__11_, issue_pkt_r_instr__10_, issue_pkt_r_instr__9_, issue_pkt_r_instr__8_, issue_pkt_r_instr__7_, issue_pkt_r_instr__6_, issue_pkt_r_instr__5_, issue_pkt_r_instr__4_, issue_pkt_r_instr__3_, issue_pkt_r_instr__2_, issue_pkt_r_instr__1_, issue_pkt_r_instr__0_, calc_status_o[305:305], calc_status_o[298:298], calc_status_o[304:304], calc_status_o[297:297], calc_status_o[303:299], calc_status_o[296:292], issue_pkt_r_imm__63_, issue_pkt_r_imm__62_, issue_pkt_r_imm__61_, issue_pkt_r_imm__60_, issue_pkt_r_imm__59_, issue_pkt_r_imm__58_, issue_pkt_r_imm__57_, issue_pkt_r_imm__56_, issue_pkt_r_imm__55_, issue_pkt_r_imm__54_, issue_pkt_r_imm__53_, issue_pkt_r_imm__52_, issue_pkt_r_imm__51_, issue_pkt_r_imm__50_, issue_pkt_r_imm__49_, issue_pkt_r_imm__48_, issue_pkt_r_imm__47_, issue_pkt_r_imm__46_, issue_pkt_r_imm__45_, issue_pkt_r_imm__44_, issue_pkt_r_imm__43_, issue_pkt_r_imm__42_, issue_pkt_r_imm__41_, issue_pkt_r_imm__40_, issue_pkt_r_imm__39_, issue_pkt_r_imm__38_, issue_pkt_r_imm__37_, issue_pkt_r_imm__36_, issue_pkt_r_imm__35_, issue_pkt_r_imm__34_, issue_pkt_r_imm__33_, issue_pkt_r_imm__32_, issue_pkt_r_imm__31_, issue_pkt_r_imm__30_, issue_pkt_r_imm__29_, issue_pkt_r_imm__28_, issue_pkt_r_imm__27_, issue_pkt_r_imm__26_, issue_pkt_r_imm__25_, issue_pkt_r_imm__24_, issue_pkt_r_imm__23_, issue_pkt_r_imm__22_, issue_pkt_r_imm__21_, issue_pkt_r_imm__20_, issue_pkt_r_imm__19_, issue_pkt_r_imm__18_, issue_pkt_r_imm__17_, issue_pkt_r_imm__16_, issue_pkt_r_imm__15_, issue_pkt_r_imm__14_, issue_pkt_r_imm__13_, issue_pkt_r_imm__12_, issue_pkt_r_imm__11_, issue_pkt_r_imm__10_, issue_pkt_r_imm__9_, issue_pkt_r_imm__8_, issue_pkt_r_imm__7_, issue_pkt_r_imm__6_, issue_pkt_r_imm__5_, issue_pkt_r_imm__4_, issue_pkt_r_imm__3_, issue_pkt_r_imm__2_, issue_pkt_r_imm__1_, issue_pkt_r_imm__0_ })
  );


  bp_be_instr_decoder
  instr_decoder
  (
    .instr_i({ issue_pkt_r_instr__31_, issue_pkt_r_instr__30_, issue_pkt_r_instr__29_, issue_pkt_r_instr__28_, issue_pkt_r_instr__27_, issue_pkt_r_instr__26_, issue_pkt_r_instr__25_, issue_pkt_r_instr__24_, issue_pkt_r_instr__23_, issue_pkt_r_instr__22_, issue_pkt_r_instr__21_, issue_pkt_r_instr__20_, issue_pkt_r_instr__19_, issue_pkt_r_instr__18_, issue_pkt_r_instr__17_, issue_pkt_r_instr__16_, issue_pkt_r_instr__15_, issue_pkt_r_instr__14_, issue_pkt_r_instr__13_, issue_pkt_r_instr__12_, issue_pkt_r_instr__11_, issue_pkt_r_instr__10_, issue_pkt_r_instr__9_, issue_pkt_r_instr__8_, issue_pkt_r_instr__7_, issue_pkt_r_instr__6_, issue_pkt_r_instr__5_, issue_pkt_r_instr__4_, issue_pkt_r_instr__3_, issue_pkt_r_instr__2_, issue_pkt_r_instr__1_, issue_pkt_r_instr__0_ }),
    .decode_o(decoded),
    .illegal_instr_o(illegal_instr_isd),
    .ret_instr_o(exc_stage_n_0__ret_instr_v_),
    .csr_instr_o(exc_stage_n_0__csr_instr_v_)
  );


  bp_be_bypass_fwd_els_p4
  int_bypass
  (
    .id_rs1_v_i(calc_status_o[305]),
    .id_rs1_addr_i(decoded[18:14]),
    .id_rs1_i(irf_rs1),
    .id_rs2_v_i(calc_status_o[298]),
    .id_rs2_addr_i(decoded[13:9]),
    .id_rs2_i(irf_rs2),
    .fwd_rd_v_i(comp_stage_n_slice_iwb_v),
    .fwd_rd_addr_i({ calc_status_o[106:102], calc_status_o[95:91], calc_status_o[84:80], calc_status_o[73:69] }),
    .fwd_rd_i(comp_stage_n[319:64]),
    .bypass_rs1_o(bypass_irs1),
    .bypass_rs2_o(bypass_irs2)
  );


  bp_be_bypass_fwd_els_p4
  fp_bypass
  (
    .id_rs1_v_i(calc_status_o[304]),
    .id_rs1_addr_i(decoded[18:14]),
    .id_rs1_i(frf_rs1),
    .id_rs2_v_i(calc_status_o[297]),
    .id_rs2_addr_i(decoded[13:9]),
    .id_rs2_i(frf_rs2),
    .fwd_rd_v_i(comp_stage_n_slice_fwb_v),
    .fwd_rd_addr_i({ calc_status_o[106:102], calc_status_o[95:91], calc_status_o[84:80], calc_status_o[73:69] }),
    .fwd_rd_i(comp_stage_n[319:64]),
    .bypass_rs1_o(bypass_frs1),
    .bypass_rs2_o(bypass_frs2)
  );


  bsg_mux_width_p64_els_p2
  bypass_xrs1_mux
  (
    .data_i({ bypass_frs1, bypass_irs1 }),
    .sel_i(calc_status_o[304]),
    .data_o(bypass_rs1)
  );


  bsg_mux_width_p64_els_p2
  bypass_xrs2_mux
  (
    .data_i({ bypass_frs2, bypass_irs2 }),
    .sel_i(calc_status_o[297]),
    .data_o(bypass_rs2)
  );


  bp_be_pipe_int
  pipe_int
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .kill_ex1_i(n_28_net_),
    .decode_i({ calc_status_o[188:188], dispatch_pkt_r_decode__fe_nop_v_, dispatch_pkt_r_decode__be_nop_v_, dispatch_pkt_r_decode__me_nop_v_, dispatch_pkt_r_decode__pipe_comp_v_, calc_status_o[291:291], dispatch_pkt_r_decode__pipe_mul_v_, dispatch_pkt_r_decode__pipe_mem_v_, dispatch_pkt_r_decode__pipe_fp_v_, dispatch_pkt_r_decode__irf_w_v_, dispatch_pkt_r_decode__frf_w_v_, dispatch_pkt_r_decode__csr_instr_v_, dispatch_pkt_r_decode__mhartid_r_v_, dispatch_pkt_r_decode__mcycle_r_v_, dispatch_pkt_r_decode__mtime_r_v_, dispatch_pkt_r_decode__minstret_r_v_, dispatch_pkt_r_decode__mtvec_rw_v_, dispatch_pkt_r_decode__mtval_rw_v_, dispatch_pkt_r_decode__mepc_rw_v_, dispatch_pkt_r_decode__mscratch_rw_v_, dispatch_pkt_r_decode__dcache_w_v_, dispatch_pkt_r_decode__dcache_r_v_, dispatch_pkt_r_decode__fp_not_int_v_, dispatch_pkt_r_decode__ret_v_, dispatch_pkt_r_decode__amo_v_, dispatch_pkt_r_decode__jmp_v_, dispatch_pkt_r_decode__br_v_, dispatch_pkt_r_decode__opw_v_, dispatch_pkt_r_decode__fu_op__fu_op__3_, dispatch_pkt_r_decode__fu_op__fu_op__2_, dispatch_pkt_r_decode__fu_op__fu_op__1_, dispatch_pkt_r_decode__fu_op__fu_op__0_, dispatch_pkt_r_decode__rs1_addr__4_, dispatch_pkt_r_decode__rs1_addr__3_, dispatch_pkt_r_decode__rs1_addr__2_, dispatch_pkt_r_decode__rs1_addr__1_, dispatch_pkt_r_decode__rs1_addr__0_, dispatch_pkt_r_decode__rs2_addr__4_, dispatch_pkt_r_decode__rs2_addr__3_, dispatch_pkt_r_decode__rs2_addr__2_, dispatch_pkt_r_decode__rs2_addr__1_, dispatch_pkt_r_decode__rs2_addr__0_, dispatch_pkt_r_decode__rd_addr__4_, dispatch_pkt_r_decode__rd_addr__3_, dispatch_pkt_r_decode__rd_addr__2_, dispatch_pkt_r_decode__rd_addr__1_, dispatch_pkt_r_decode__rd_addr__0_, dispatch_pkt_r_decode__src1_sel_, dispatch_pkt_r_decode__src2_sel_, dispatch_pkt_r_decode__baddr_sel_, dispatch_pkt_r_decode__result_sel_ }),
    .pc_i(calc_status_o[187:124]),
    .rs1_i({ dispatch_pkt_r_rs1__63_, dispatch_pkt_r_rs1__62_, dispatch_pkt_r_rs1__61_, dispatch_pkt_r_rs1__60_, dispatch_pkt_r_rs1__59_, dispatch_pkt_r_rs1__58_, dispatch_pkt_r_rs1__57_, dispatch_pkt_r_rs1__56_, dispatch_pkt_r_rs1__55_, dispatch_pkt_r_rs1__54_, dispatch_pkt_r_rs1__53_, dispatch_pkt_r_rs1__52_, dispatch_pkt_r_rs1__51_, dispatch_pkt_r_rs1__50_, dispatch_pkt_r_rs1__49_, dispatch_pkt_r_rs1__48_, dispatch_pkt_r_rs1__47_, dispatch_pkt_r_rs1__46_, dispatch_pkt_r_rs1__45_, dispatch_pkt_r_rs1__44_, dispatch_pkt_r_rs1__43_, dispatch_pkt_r_rs1__42_, dispatch_pkt_r_rs1__41_, dispatch_pkt_r_rs1__40_, dispatch_pkt_r_rs1__39_, dispatch_pkt_r_rs1__38_, dispatch_pkt_r_rs1__37_, dispatch_pkt_r_rs1__36_, dispatch_pkt_r_rs1__35_, dispatch_pkt_r_rs1__34_, dispatch_pkt_r_rs1__33_, dispatch_pkt_r_rs1__32_, dispatch_pkt_r_rs1__31_, dispatch_pkt_r_rs1__30_, dispatch_pkt_r_rs1__29_, dispatch_pkt_r_rs1__28_, dispatch_pkt_r_rs1__27_, dispatch_pkt_r_rs1__26_, dispatch_pkt_r_rs1__25_, dispatch_pkt_r_rs1__24_, dispatch_pkt_r_rs1__23_, dispatch_pkt_r_rs1__22_, dispatch_pkt_r_rs1__21_, dispatch_pkt_r_rs1__20_, dispatch_pkt_r_rs1__19_, dispatch_pkt_r_rs1__18_, dispatch_pkt_r_rs1__17_, dispatch_pkt_r_rs1__16_, dispatch_pkt_r_rs1__15_, dispatch_pkt_r_rs1__14_, dispatch_pkt_r_rs1__13_, dispatch_pkt_r_rs1__12_, dispatch_pkt_r_rs1__11_, dispatch_pkt_r_rs1__10_, dispatch_pkt_r_rs1__9_, dispatch_pkt_r_rs1__8_, dispatch_pkt_r_rs1__7_, dispatch_pkt_r_rs1__6_, dispatch_pkt_r_rs1__5_, dispatch_pkt_r_rs1__4_, dispatch_pkt_r_rs1__3_, dispatch_pkt_r_rs1__2_, dispatch_pkt_r_rs1__1_, dispatch_pkt_r_rs1__0_ }),
    .rs2_i({ dispatch_pkt_r_rs2__63_, dispatch_pkt_r_rs2__62_, dispatch_pkt_r_rs2__61_, dispatch_pkt_r_rs2__60_, dispatch_pkt_r_rs2__59_, dispatch_pkt_r_rs2__58_, dispatch_pkt_r_rs2__57_, dispatch_pkt_r_rs2__56_, dispatch_pkt_r_rs2__55_, dispatch_pkt_r_rs2__54_, dispatch_pkt_r_rs2__53_, dispatch_pkt_r_rs2__52_, dispatch_pkt_r_rs2__51_, dispatch_pkt_r_rs2__50_, dispatch_pkt_r_rs2__49_, dispatch_pkt_r_rs2__48_, dispatch_pkt_r_rs2__47_, dispatch_pkt_r_rs2__46_, dispatch_pkt_r_rs2__45_, dispatch_pkt_r_rs2__44_, dispatch_pkt_r_rs2__43_, dispatch_pkt_r_rs2__42_, dispatch_pkt_r_rs2__41_, dispatch_pkt_r_rs2__40_, dispatch_pkt_r_rs2__39_, dispatch_pkt_r_rs2__38_, dispatch_pkt_r_rs2__37_, dispatch_pkt_r_rs2__36_, dispatch_pkt_r_rs2__35_, dispatch_pkt_r_rs2__34_, dispatch_pkt_r_rs2__33_, dispatch_pkt_r_rs2__32_, dispatch_pkt_r_rs2__31_, dispatch_pkt_r_rs2__30_, dispatch_pkt_r_rs2__29_, dispatch_pkt_r_rs2__28_, dispatch_pkt_r_rs2__27_, dispatch_pkt_r_rs2__26_, dispatch_pkt_r_rs2__25_, dispatch_pkt_r_rs2__24_, dispatch_pkt_r_rs2__23_, dispatch_pkt_r_rs2__22_, dispatch_pkt_r_rs2__21_, dispatch_pkt_r_rs2__20_, dispatch_pkt_r_rs2__19_, dispatch_pkt_r_rs2__18_, dispatch_pkt_r_rs2__17_, dispatch_pkt_r_rs2__16_, dispatch_pkt_r_rs2__15_, dispatch_pkt_r_rs2__14_, dispatch_pkt_r_rs2__13_, dispatch_pkt_r_rs2__12_, dispatch_pkt_r_rs2__11_, dispatch_pkt_r_rs2__10_, dispatch_pkt_r_rs2__9_, dispatch_pkt_r_rs2__8_, dispatch_pkt_r_rs2__7_, dispatch_pkt_r_rs2__6_, dispatch_pkt_r_rs2__5_, dispatch_pkt_r_rs2__4_, dispatch_pkt_r_rs2__3_, dispatch_pkt_r_rs2__2_, dispatch_pkt_r_rs2__1_, dispatch_pkt_r_rs2__0_ }),
    .imm_i({ dispatch_pkt_r_imm__63_, dispatch_pkt_r_imm__62_, dispatch_pkt_r_imm__61_, dispatch_pkt_r_imm__60_, dispatch_pkt_r_imm__59_, dispatch_pkt_r_imm__58_, dispatch_pkt_r_imm__57_, dispatch_pkt_r_imm__56_, dispatch_pkt_r_imm__55_, dispatch_pkt_r_imm__54_, dispatch_pkt_r_imm__53_, dispatch_pkt_r_imm__52_, dispatch_pkt_r_imm__51_, dispatch_pkt_r_imm__50_, dispatch_pkt_r_imm__49_, dispatch_pkt_r_imm__48_, dispatch_pkt_r_imm__47_, dispatch_pkt_r_imm__46_, dispatch_pkt_r_imm__45_, dispatch_pkt_r_imm__44_, dispatch_pkt_r_imm__43_, dispatch_pkt_r_imm__42_, dispatch_pkt_r_imm__41_, dispatch_pkt_r_imm__40_, dispatch_pkt_r_imm__39_, dispatch_pkt_r_imm__38_, dispatch_pkt_r_imm__37_, dispatch_pkt_r_imm__36_, dispatch_pkt_r_imm__35_, dispatch_pkt_r_imm__34_, dispatch_pkt_r_imm__33_, dispatch_pkt_r_imm__32_, dispatch_pkt_r_imm__31_, dispatch_pkt_r_imm__30_, dispatch_pkt_r_imm__29_, dispatch_pkt_r_imm__28_, dispatch_pkt_r_imm__27_, dispatch_pkt_r_imm__26_, dispatch_pkt_r_imm__25_, dispatch_pkt_r_imm__24_, dispatch_pkt_r_imm__23_, dispatch_pkt_r_imm__22_, dispatch_pkt_r_imm__21_, dispatch_pkt_r_imm__20_, dispatch_pkt_r_imm__19_, dispatch_pkt_r_imm__18_, dispatch_pkt_r_imm__17_, dispatch_pkt_r_imm__16_, dispatch_pkt_r_imm__15_, dispatch_pkt_r_imm__14_, dispatch_pkt_r_imm__13_, dispatch_pkt_r_imm__12_, dispatch_pkt_r_imm__11_, dispatch_pkt_r_imm__10_, dispatch_pkt_r_imm__9_, dispatch_pkt_r_imm__8_, dispatch_pkt_r_imm__7_, dispatch_pkt_r_imm__6_, dispatch_pkt_r_imm__5_, dispatch_pkt_r_imm__4_, dispatch_pkt_r_imm__3_, dispatch_pkt_r_imm__2_, dispatch_pkt_r_imm__1_, dispatch_pkt_r_imm__0_ }),
    .data_o(pipe_int_data_lo),
    .br_tgt_o(calc_status_o[290:227])
  );


  bp_be_pipe_mul
  pipe_mul
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .kill_ex1_i(exc_stage_n_1__poison_v_),
    .kill_ex2_i(exc_stage_n_2__poison_v_),
    .decode_i({ calc_status_o[188:188], dispatch_pkt_r_decode__fe_nop_v_, dispatch_pkt_r_decode__be_nop_v_, dispatch_pkt_r_decode__me_nop_v_, dispatch_pkt_r_decode__pipe_comp_v_, calc_status_o[291:291], dispatch_pkt_r_decode__pipe_mul_v_, dispatch_pkt_r_decode__pipe_mem_v_, dispatch_pkt_r_decode__pipe_fp_v_, dispatch_pkt_r_decode__irf_w_v_, dispatch_pkt_r_decode__frf_w_v_, dispatch_pkt_r_decode__csr_instr_v_, dispatch_pkt_r_decode__mhartid_r_v_, dispatch_pkt_r_decode__mcycle_r_v_, dispatch_pkt_r_decode__mtime_r_v_, dispatch_pkt_r_decode__minstret_r_v_, dispatch_pkt_r_decode__mtvec_rw_v_, dispatch_pkt_r_decode__mtval_rw_v_, dispatch_pkt_r_decode__mepc_rw_v_, dispatch_pkt_r_decode__mscratch_rw_v_, dispatch_pkt_r_decode__dcache_w_v_, dispatch_pkt_r_decode__dcache_r_v_, dispatch_pkt_r_decode__fp_not_int_v_, dispatch_pkt_r_decode__ret_v_, dispatch_pkt_r_decode__amo_v_, dispatch_pkt_r_decode__jmp_v_, dispatch_pkt_r_decode__br_v_, dispatch_pkt_r_decode__opw_v_, dispatch_pkt_r_decode__fu_op__fu_op__3_, dispatch_pkt_r_decode__fu_op__fu_op__2_, dispatch_pkt_r_decode__fu_op__fu_op__1_, dispatch_pkt_r_decode__fu_op__fu_op__0_, dispatch_pkt_r_decode__rs1_addr__4_, dispatch_pkt_r_decode__rs1_addr__3_, dispatch_pkt_r_decode__rs1_addr__2_, dispatch_pkt_r_decode__rs1_addr__1_, dispatch_pkt_r_decode__rs1_addr__0_, dispatch_pkt_r_decode__rs2_addr__4_, dispatch_pkt_r_decode__rs2_addr__3_, dispatch_pkt_r_decode__rs2_addr__2_, dispatch_pkt_r_decode__rs2_addr__1_, dispatch_pkt_r_decode__rs2_addr__0_, dispatch_pkt_r_decode__rd_addr__4_, dispatch_pkt_r_decode__rd_addr__3_, dispatch_pkt_r_decode__rd_addr__2_, dispatch_pkt_r_decode__rd_addr__1_, dispatch_pkt_r_decode__rd_addr__0_, dispatch_pkt_r_decode__src1_sel_, dispatch_pkt_r_decode__src2_sel_, dispatch_pkt_r_decode__baddr_sel_, dispatch_pkt_r_decode__result_sel_ }),
    .rs1_i({ dispatch_pkt_r_rs1__63_, dispatch_pkt_r_rs1__62_, dispatch_pkt_r_rs1__61_, dispatch_pkt_r_rs1__60_, dispatch_pkt_r_rs1__59_, dispatch_pkt_r_rs1__58_, dispatch_pkt_r_rs1__57_, dispatch_pkt_r_rs1__56_, dispatch_pkt_r_rs1__55_, dispatch_pkt_r_rs1__54_, dispatch_pkt_r_rs1__53_, dispatch_pkt_r_rs1__52_, dispatch_pkt_r_rs1__51_, dispatch_pkt_r_rs1__50_, dispatch_pkt_r_rs1__49_, dispatch_pkt_r_rs1__48_, dispatch_pkt_r_rs1__47_, dispatch_pkt_r_rs1__46_, dispatch_pkt_r_rs1__45_, dispatch_pkt_r_rs1__44_, dispatch_pkt_r_rs1__43_, dispatch_pkt_r_rs1__42_, dispatch_pkt_r_rs1__41_, dispatch_pkt_r_rs1__40_, dispatch_pkt_r_rs1__39_, dispatch_pkt_r_rs1__38_, dispatch_pkt_r_rs1__37_, dispatch_pkt_r_rs1__36_, dispatch_pkt_r_rs1__35_, dispatch_pkt_r_rs1__34_, dispatch_pkt_r_rs1__33_, dispatch_pkt_r_rs1__32_, dispatch_pkt_r_rs1__31_, dispatch_pkt_r_rs1__30_, dispatch_pkt_r_rs1__29_, dispatch_pkt_r_rs1__28_, dispatch_pkt_r_rs1__27_, dispatch_pkt_r_rs1__26_, dispatch_pkt_r_rs1__25_, dispatch_pkt_r_rs1__24_, dispatch_pkt_r_rs1__23_, dispatch_pkt_r_rs1__22_, dispatch_pkt_r_rs1__21_, dispatch_pkt_r_rs1__20_, dispatch_pkt_r_rs1__19_, dispatch_pkt_r_rs1__18_, dispatch_pkt_r_rs1__17_, dispatch_pkt_r_rs1__16_, dispatch_pkt_r_rs1__15_, dispatch_pkt_r_rs1__14_, dispatch_pkt_r_rs1__13_, dispatch_pkt_r_rs1__12_, dispatch_pkt_r_rs1__11_, dispatch_pkt_r_rs1__10_, dispatch_pkt_r_rs1__9_, dispatch_pkt_r_rs1__8_, dispatch_pkt_r_rs1__7_, dispatch_pkt_r_rs1__6_, dispatch_pkt_r_rs1__5_, dispatch_pkt_r_rs1__4_, dispatch_pkt_r_rs1__3_, dispatch_pkt_r_rs1__2_, dispatch_pkt_r_rs1__1_, dispatch_pkt_r_rs1__0_ }),
    .rs2_i({ dispatch_pkt_r_rs2__63_, dispatch_pkt_r_rs2__62_, dispatch_pkt_r_rs2__61_, dispatch_pkt_r_rs2__60_, dispatch_pkt_r_rs2__59_, dispatch_pkt_r_rs2__58_, dispatch_pkt_r_rs2__57_, dispatch_pkt_r_rs2__56_, dispatch_pkt_r_rs2__55_, dispatch_pkt_r_rs2__54_, dispatch_pkt_r_rs2__53_, dispatch_pkt_r_rs2__52_, dispatch_pkt_r_rs2__51_, dispatch_pkt_r_rs2__50_, dispatch_pkt_r_rs2__49_, dispatch_pkt_r_rs2__48_, dispatch_pkt_r_rs2__47_, dispatch_pkt_r_rs2__46_, dispatch_pkt_r_rs2__45_, dispatch_pkt_r_rs2__44_, dispatch_pkt_r_rs2__43_, dispatch_pkt_r_rs2__42_, dispatch_pkt_r_rs2__41_, dispatch_pkt_r_rs2__40_, dispatch_pkt_r_rs2__39_, dispatch_pkt_r_rs2__38_, dispatch_pkt_r_rs2__37_, dispatch_pkt_r_rs2__36_, dispatch_pkt_r_rs2__35_, dispatch_pkt_r_rs2__34_, dispatch_pkt_r_rs2__33_, dispatch_pkt_r_rs2__32_, dispatch_pkt_r_rs2__31_, dispatch_pkt_r_rs2__30_, dispatch_pkt_r_rs2__29_, dispatch_pkt_r_rs2__28_, dispatch_pkt_r_rs2__27_, dispatch_pkt_r_rs2__26_, dispatch_pkt_r_rs2__25_, dispatch_pkt_r_rs2__24_, dispatch_pkt_r_rs2__23_, dispatch_pkt_r_rs2__22_, dispatch_pkt_r_rs2__21_, dispatch_pkt_r_rs2__20_, dispatch_pkt_r_rs2__19_, dispatch_pkt_r_rs2__18_, dispatch_pkt_r_rs2__17_, dispatch_pkt_r_rs2__16_, dispatch_pkt_r_rs2__15_, dispatch_pkt_r_rs2__14_, dispatch_pkt_r_rs2__13_, dispatch_pkt_r_rs2__12_, dispatch_pkt_r_rs2__11_, dispatch_pkt_r_rs2__10_, dispatch_pkt_r_rs2__9_, dispatch_pkt_r_rs2__8_, dispatch_pkt_r_rs2__7_, dispatch_pkt_r_rs2__6_, dispatch_pkt_r_rs2__5_, dispatch_pkt_r_rs2__4_, dispatch_pkt_r_rs2__3_, dispatch_pkt_r_rs2__2_, dispatch_pkt_r_rs2__1_, dispatch_pkt_r_rs2__0_ }),
    .data_o(pipe_mul_data_lo)
  );


  bp_be_pipe_mem_vaddr_width_p39_lce_sets_p64_cce_block_size_in_bytes_p64_core_els_p1
  pipe_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .kill_ex1_i(exc_stage_n_1__poison_v_),
    .kill_ex2_i(exc_stage_n_2__poison_v_),
    .kill_ex3_i(exc_stage_n_3__poison_v_),
    .decode_i({ calc_status_o[188:188], dispatch_pkt_r_decode__fe_nop_v_, dispatch_pkt_r_decode__be_nop_v_, dispatch_pkt_r_decode__me_nop_v_, dispatch_pkt_r_decode__pipe_comp_v_, calc_status_o[291:291], dispatch_pkt_r_decode__pipe_mul_v_, dispatch_pkt_r_decode__pipe_mem_v_, dispatch_pkt_r_decode__pipe_fp_v_, dispatch_pkt_r_decode__irf_w_v_, dispatch_pkt_r_decode__frf_w_v_, dispatch_pkt_r_decode__csr_instr_v_, dispatch_pkt_r_decode__mhartid_r_v_, dispatch_pkt_r_decode__mcycle_r_v_, dispatch_pkt_r_decode__mtime_r_v_, dispatch_pkt_r_decode__minstret_r_v_, dispatch_pkt_r_decode__mtvec_rw_v_, dispatch_pkt_r_decode__mtval_rw_v_, dispatch_pkt_r_decode__mepc_rw_v_, dispatch_pkt_r_decode__mscratch_rw_v_, dispatch_pkt_r_decode__dcache_w_v_, dispatch_pkt_r_decode__dcache_r_v_, dispatch_pkt_r_decode__fp_not_int_v_, dispatch_pkt_r_decode__ret_v_, dispatch_pkt_r_decode__amo_v_, dispatch_pkt_r_decode__jmp_v_, dispatch_pkt_r_decode__br_v_, dispatch_pkt_r_decode__opw_v_, dispatch_pkt_r_decode__fu_op__fu_op__3_, dispatch_pkt_r_decode__fu_op__fu_op__2_, dispatch_pkt_r_decode__fu_op__fu_op__1_, dispatch_pkt_r_decode__fu_op__fu_op__0_, dispatch_pkt_r_decode__rs1_addr__4_, dispatch_pkt_r_decode__rs1_addr__3_, dispatch_pkt_r_decode__rs1_addr__2_, dispatch_pkt_r_decode__rs1_addr__1_, dispatch_pkt_r_decode__rs1_addr__0_, dispatch_pkt_r_decode__rs2_addr__4_, dispatch_pkt_r_decode__rs2_addr__3_, dispatch_pkt_r_decode__rs2_addr__2_, dispatch_pkt_r_decode__rs2_addr__1_, dispatch_pkt_r_decode__rs2_addr__0_, dispatch_pkt_r_decode__rd_addr__4_, dispatch_pkt_r_decode__rd_addr__3_, dispatch_pkt_r_decode__rd_addr__2_, dispatch_pkt_r_decode__rd_addr__1_, dispatch_pkt_r_decode__rd_addr__0_, dispatch_pkt_r_decode__src1_sel_, dispatch_pkt_r_decode__src2_sel_, dispatch_pkt_r_decode__baddr_sel_, dispatch_pkt_r_decode__result_sel_ }),
    .rs1_i({ dispatch_pkt_r_rs1__63_, dispatch_pkt_r_rs1__62_, dispatch_pkt_r_rs1__61_, dispatch_pkt_r_rs1__60_, dispatch_pkt_r_rs1__59_, dispatch_pkt_r_rs1__58_, dispatch_pkt_r_rs1__57_, dispatch_pkt_r_rs1__56_, dispatch_pkt_r_rs1__55_, dispatch_pkt_r_rs1__54_, dispatch_pkt_r_rs1__53_, dispatch_pkt_r_rs1__52_, dispatch_pkt_r_rs1__51_, dispatch_pkt_r_rs1__50_, dispatch_pkt_r_rs1__49_, dispatch_pkt_r_rs1__48_, dispatch_pkt_r_rs1__47_, dispatch_pkt_r_rs1__46_, dispatch_pkt_r_rs1__45_, dispatch_pkt_r_rs1__44_, dispatch_pkt_r_rs1__43_, dispatch_pkt_r_rs1__42_, dispatch_pkt_r_rs1__41_, dispatch_pkt_r_rs1__40_, dispatch_pkt_r_rs1__39_, dispatch_pkt_r_rs1__38_, dispatch_pkt_r_rs1__37_, dispatch_pkt_r_rs1__36_, dispatch_pkt_r_rs1__35_, dispatch_pkt_r_rs1__34_, dispatch_pkt_r_rs1__33_, dispatch_pkt_r_rs1__32_, dispatch_pkt_r_rs1__31_, dispatch_pkt_r_rs1__30_, dispatch_pkt_r_rs1__29_, dispatch_pkt_r_rs1__28_, dispatch_pkt_r_rs1__27_, dispatch_pkt_r_rs1__26_, dispatch_pkt_r_rs1__25_, dispatch_pkt_r_rs1__24_, dispatch_pkt_r_rs1__23_, dispatch_pkt_r_rs1__22_, dispatch_pkt_r_rs1__21_, dispatch_pkt_r_rs1__20_, dispatch_pkt_r_rs1__19_, dispatch_pkt_r_rs1__18_, dispatch_pkt_r_rs1__17_, dispatch_pkt_r_rs1__16_, dispatch_pkt_r_rs1__15_, dispatch_pkt_r_rs1__14_, dispatch_pkt_r_rs1__13_, dispatch_pkt_r_rs1__12_, dispatch_pkt_r_rs1__11_, dispatch_pkt_r_rs1__10_, dispatch_pkt_r_rs1__9_, dispatch_pkt_r_rs1__8_, dispatch_pkt_r_rs1__7_, dispatch_pkt_r_rs1__6_, dispatch_pkt_r_rs1__5_, dispatch_pkt_r_rs1__4_, dispatch_pkt_r_rs1__3_, dispatch_pkt_r_rs1__2_, dispatch_pkt_r_rs1__1_, dispatch_pkt_r_rs1__0_ }),
    .rs2_i({ dispatch_pkt_r_rs2__63_, dispatch_pkt_r_rs2__62_, dispatch_pkt_r_rs2__61_, dispatch_pkt_r_rs2__60_, dispatch_pkt_r_rs2__59_, dispatch_pkt_r_rs2__58_, dispatch_pkt_r_rs2__57_, dispatch_pkt_r_rs2__56_, dispatch_pkt_r_rs2__55_, dispatch_pkt_r_rs2__54_, dispatch_pkt_r_rs2__53_, dispatch_pkt_r_rs2__52_, dispatch_pkt_r_rs2__51_, dispatch_pkt_r_rs2__50_, dispatch_pkt_r_rs2__49_, dispatch_pkt_r_rs2__48_, dispatch_pkt_r_rs2__47_, dispatch_pkt_r_rs2__46_, dispatch_pkt_r_rs2__45_, dispatch_pkt_r_rs2__44_, dispatch_pkt_r_rs2__43_, dispatch_pkt_r_rs2__42_, dispatch_pkt_r_rs2__41_, dispatch_pkt_r_rs2__40_, dispatch_pkt_r_rs2__39_, dispatch_pkt_r_rs2__38_, dispatch_pkt_r_rs2__37_, dispatch_pkt_r_rs2__36_, dispatch_pkt_r_rs2__35_, dispatch_pkt_r_rs2__34_, dispatch_pkt_r_rs2__33_, dispatch_pkt_r_rs2__32_, dispatch_pkt_r_rs2__31_, dispatch_pkt_r_rs2__30_, dispatch_pkt_r_rs2__29_, dispatch_pkt_r_rs2__28_, dispatch_pkt_r_rs2__27_, dispatch_pkt_r_rs2__26_, dispatch_pkt_r_rs2__25_, dispatch_pkt_r_rs2__24_, dispatch_pkt_r_rs2__23_, dispatch_pkt_r_rs2__22_, dispatch_pkt_r_rs2__21_, dispatch_pkt_r_rs2__20_, dispatch_pkt_r_rs2__19_, dispatch_pkt_r_rs2__18_, dispatch_pkt_r_rs2__17_, dispatch_pkt_r_rs2__16_, dispatch_pkt_r_rs2__15_, dispatch_pkt_r_rs2__14_, dispatch_pkt_r_rs2__13_, dispatch_pkt_r_rs2__12_, dispatch_pkt_r_rs2__11_, dispatch_pkt_r_rs2__10_, dispatch_pkt_r_rs2__9_, dispatch_pkt_r_rs2__8_, dispatch_pkt_r_rs2__7_, dispatch_pkt_r_rs2__6_, dispatch_pkt_r_rs2__5_, dispatch_pkt_r_rs2__4_, dispatch_pkt_r_rs2__3_, dispatch_pkt_r_rs2__2_, dispatch_pkt_r_rs2__1_, dispatch_pkt_r_rs2__0_ }),
    .imm_i({ dispatch_pkt_r_imm__63_, dispatch_pkt_r_imm__62_, dispatch_pkt_r_imm__61_, dispatch_pkt_r_imm__60_, dispatch_pkt_r_imm__59_, dispatch_pkt_r_imm__58_, dispatch_pkt_r_imm__57_, dispatch_pkt_r_imm__56_, dispatch_pkt_r_imm__55_, dispatch_pkt_r_imm__54_, dispatch_pkt_r_imm__53_, dispatch_pkt_r_imm__52_, dispatch_pkt_r_imm__51_, dispatch_pkt_r_imm__50_, dispatch_pkt_r_imm__49_, dispatch_pkt_r_imm__48_, dispatch_pkt_r_imm__47_, dispatch_pkt_r_imm__46_, dispatch_pkt_r_imm__45_, dispatch_pkt_r_imm__44_, dispatch_pkt_r_imm__43_, dispatch_pkt_r_imm__42_, dispatch_pkt_r_imm__41_, dispatch_pkt_r_imm__40_, dispatch_pkt_r_imm__39_, dispatch_pkt_r_imm__38_, dispatch_pkt_r_imm__37_, dispatch_pkt_r_imm__36_, dispatch_pkt_r_imm__35_, dispatch_pkt_r_imm__34_, dispatch_pkt_r_imm__33_, dispatch_pkt_r_imm__32_, dispatch_pkt_r_imm__31_, dispatch_pkt_r_imm__30_, dispatch_pkt_r_imm__29_, dispatch_pkt_r_imm__28_, dispatch_pkt_r_imm__27_, dispatch_pkt_r_imm__26_, dispatch_pkt_r_imm__25_, dispatch_pkt_r_imm__24_, dispatch_pkt_r_imm__23_, dispatch_pkt_r_imm__22_, dispatch_pkt_r_imm__21_, dispatch_pkt_r_imm__20_, dispatch_pkt_r_imm__19_, dispatch_pkt_r_imm__18_, dispatch_pkt_r_imm__17_, dispatch_pkt_r_imm__16_, dispatch_pkt_r_imm__15_, dispatch_pkt_r_imm__14_, dispatch_pkt_r_imm__13_, dispatch_pkt_r_imm__12_, dispatch_pkt_r_imm__11_, dispatch_pkt_r_imm__10_, dispatch_pkt_r_imm__9_, dispatch_pkt_r_imm__8_, dispatch_pkt_r_imm__7_, dispatch_pkt_r_imm__6_, dispatch_pkt_r_imm__5_, dispatch_pkt_r_imm__4_, dispatch_pkt_r_imm__3_, dispatch_pkt_r_imm__2_, dispatch_pkt_r_imm__1_, dispatch_pkt_r_imm__0_ }),
    .mmu_cmd_o(mmu_cmd_o),
    .mmu_cmd_v_o(mmu_cmd_v_o),
    .mmu_cmd_ready_i(mmu_cmd_ready_i),
    .mmu_resp_i(mmu_resp_i),
    .mmu_resp_v_i(mmu_resp_v_i),
    .mmu_resp_ready_o(mmu_resp_ready_o),
    .data_o(pipe_mem_data_lo),
    .cache_miss_o(exc_stage_n_3__cache_miss_v_),
    .mhartid_i(proc_cfg_i[2]),
    .mcycle_i(cycle_cnt_lo),
    .mtime_i(time_cnt_lo),
    .minstret_i(instret_cnt_lo),
    .mtvec_o(mtvec_o),
    .mtvec_w_v_o(mtvec_w_v_o),
    .mtvec_i(mtvec_i),
    .mtval_o(mtval_lo),
    .mtval_w_v_o(mtval_w_v_lo),
    .mtval_i(mtval_li),
    .mepc_o(mepc_o),
    .mepc_w_v_o(mepc_w_v_o),
    .mepc_i(mepc_i),
    .mscratch_o(mscratch_lo),
    .mscratch_w_v_o(mscratch_w_v_lo),
    .mscratch_i(mscratch_li)
  );


  bp_be_pipe_fp
  pipe_fp
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .kill_ex1_i(exc_stage_n_1__poison_v_),
    .kill_ex2_i(exc_stage_n_2__poison_v_),
    .kill_ex3_i(exc_stage_n_3__poison_v_),
    .kill_ex4_i(exc_stage_n_4__poison_v_),
    .decode_i({ calc_status_o[188:188], dispatch_pkt_r_decode__fe_nop_v_, dispatch_pkt_r_decode__be_nop_v_, dispatch_pkt_r_decode__me_nop_v_, dispatch_pkt_r_decode__pipe_comp_v_, calc_status_o[291:291], dispatch_pkt_r_decode__pipe_mul_v_, dispatch_pkt_r_decode__pipe_mem_v_, dispatch_pkt_r_decode__pipe_fp_v_, dispatch_pkt_r_decode__irf_w_v_, dispatch_pkt_r_decode__frf_w_v_, dispatch_pkt_r_decode__csr_instr_v_, dispatch_pkt_r_decode__mhartid_r_v_, dispatch_pkt_r_decode__mcycle_r_v_, dispatch_pkt_r_decode__mtime_r_v_, dispatch_pkt_r_decode__minstret_r_v_, dispatch_pkt_r_decode__mtvec_rw_v_, dispatch_pkt_r_decode__mtval_rw_v_, dispatch_pkt_r_decode__mepc_rw_v_, dispatch_pkt_r_decode__mscratch_rw_v_, dispatch_pkt_r_decode__dcache_w_v_, dispatch_pkt_r_decode__dcache_r_v_, dispatch_pkt_r_decode__fp_not_int_v_, dispatch_pkt_r_decode__ret_v_, dispatch_pkt_r_decode__amo_v_, dispatch_pkt_r_decode__jmp_v_, dispatch_pkt_r_decode__br_v_, dispatch_pkt_r_decode__opw_v_, dispatch_pkt_r_decode__fu_op__fu_op__3_, dispatch_pkt_r_decode__fu_op__fu_op__2_, dispatch_pkt_r_decode__fu_op__fu_op__1_, dispatch_pkt_r_decode__fu_op__fu_op__0_, dispatch_pkt_r_decode__rs1_addr__4_, dispatch_pkt_r_decode__rs1_addr__3_, dispatch_pkt_r_decode__rs1_addr__2_, dispatch_pkt_r_decode__rs1_addr__1_, dispatch_pkt_r_decode__rs1_addr__0_, dispatch_pkt_r_decode__rs2_addr__4_, dispatch_pkt_r_decode__rs2_addr__3_, dispatch_pkt_r_decode__rs2_addr__2_, dispatch_pkt_r_decode__rs2_addr__1_, dispatch_pkt_r_decode__rs2_addr__0_, dispatch_pkt_r_decode__rd_addr__4_, dispatch_pkt_r_decode__rd_addr__3_, dispatch_pkt_r_decode__rd_addr__2_, dispatch_pkt_r_decode__rd_addr__1_, dispatch_pkt_r_decode__rd_addr__0_, dispatch_pkt_r_decode__src1_sel_, dispatch_pkt_r_decode__src2_sel_, dispatch_pkt_r_decode__baddr_sel_, dispatch_pkt_r_decode__result_sel_ }),
    .rs1_i({ dispatch_pkt_r_rs1__63_, dispatch_pkt_r_rs1__62_, dispatch_pkt_r_rs1__61_, dispatch_pkt_r_rs1__60_, dispatch_pkt_r_rs1__59_, dispatch_pkt_r_rs1__58_, dispatch_pkt_r_rs1__57_, dispatch_pkt_r_rs1__56_, dispatch_pkt_r_rs1__55_, dispatch_pkt_r_rs1__54_, dispatch_pkt_r_rs1__53_, dispatch_pkt_r_rs1__52_, dispatch_pkt_r_rs1__51_, dispatch_pkt_r_rs1__50_, dispatch_pkt_r_rs1__49_, dispatch_pkt_r_rs1__48_, dispatch_pkt_r_rs1__47_, dispatch_pkt_r_rs1__46_, dispatch_pkt_r_rs1__45_, dispatch_pkt_r_rs1__44_, dispatch_pkt_r_rs1__43_, dispatch_pkt_r_rs1__42_, dispatch_pkt_r_rs1__41_, dispatch_pkt_r_rs1__40_, dispatch_pkt_r_rs1__39_, dispatch_pkt_r_rs1__38_, dispatch_pkt_r_rs1__37_, dispatch_pkt_r_rs1__36_, dispatch_pkt_r_rs1__35_, dispatch_pkt_r_rs1__34_, dispatch_pkt_r_rs1__33_, dispatch_pkt_r_rs1__32_, dispatch_pkt_r_rs1__31_, dispatch_pkt_r_rs1__30_, dispatch_pkt_r_rs1__29_, dispatch_pkt_r_rs1__28_, dispatch_pkt_r_rs1__27_, dispatch_pkt_r_rs1__26_, dispatch_pkt_r_rs1__25_, dispatch_pkt_r_rs1__24_, dispatch_pkt_r_rs1__23_, dispatch_pkt_r_rs1__22_, dispatch_pkt_r_rs1__21_, dispatch_pkt_r_rs1__20_, dispatch_pkt_r_rs1__19_, dispatch_pkt_r_rs1__18_, dispatch_pkt_r_rs1__17_, dispatch_pkt_r_rs1__16_, dispatch_pkt_r_rs1__15_, dispatch_pkt_r_rs1__14_, dispatch_pkt_r_rs1__13_, dispatch_pkt_r_rs1__12_, dispatch_pkt_r_rs1__11_, dispatch_pkt_r_rs1__10_, dispatch_pkt_r_rs1__9_, dispatch_pkt_r_rs1__8_, dispatch_pkt_r_rs1__7_, dispatch_pkt_r_rs1__6_, dispatch_pkt_r_rs1__5_, dispatch_pkt_r_rs1__4_, dispatch_pkt_r_rs1__3_, dispatch_pkt_r_rs1__2_, dispatch_pkt_r_rs1__1_, dispatch_pkt_r_rs1__0_ }),
    .rs2_i({ dispatch_pkt_r_rs2__63_, dispatch_pkt_r_rs2__62_, dispatch_pkt_r_rs2__61_, dispatch_pkt_r_rs2__60_, dispatch_pkt_r_rs2__59_, dispatch_pkt_r_rs2__58_, dispatch_pkt_r_rs2__57_, dispatch_pkt_r_rs2__56_, dispatch_pkt_r_rs2__55_, dispatch_pkt_r_rs2__54_, dispatch_pkt_r_rs2__53_, dispatch_pkt_r_rs2__52_, dispatch_pkt_r_rs2__51_, dispatch_pkt_r_rs2__50_, dispatch_pkt_r_rs2__49_, dispatch_pkt_r_rs2__48_, dispatch_pkt_r_rs2__47_, dispatch_pkt_r_rs2__46_, dispatch_pkt_r_rs2__45_, dispatch_pkt_r_rs2__44_, dispatch_pkt_r_rs2__43_, dispatch_pkt_r_rs2__42_, dispatch_pkt_r_rs2__41_, dispatch_pkt_r_rs2__40_, dispatch_pkt_r_rs2__39_, dispatch_pkt_r_rs2__38_, dispatch_pkt_r_rs2__37_, dispatch_pkt_r_rs2__36_, dispatch_pkt_r_rs2__35_, dispatch_pkt_r_rs2__34_, dispatch_pkt_r_rs2__33_, dispatch_pkt_r_rs2__32_, dispatch_pkt_r_rs2__31_, dispatch_pkt_r_rs2__30_, dispatch_pkt_r_rs2__29_, dispatch_pkt_r_rs2__28_, dispatch_pkt_r_rs2__27_, dispatch_pkt_r_rs2__26_, dispatch_pkt_r_rs2__25_, dispatch_pkt_r_rs2__24_, dispatch_pkt_r_rs2__23_, dispatch_pkt_r_rs2__22_, dispatch_pkt_r_rs2__21_, dispatch_pkt_r_rs2__20_, dispatch_pkt_r_rs2__19_, dispatch_pkt_r_rs2__18_, dispatch_pkt_r_rs2__17_, dispatch_pkt_r_rs2__16_, dispatch_pkt_r_rs2__15_, dispatch_pkt_r_rs2__14_, dispatch_pkt_r_rs2__13_, dispatch_pkt_r_rs2__12_, dispatch_pkt_r_rs2__11_, dispatch_pkt_r_rs2__10_, dispatch_pkt_r_rs2__9_, dispatch_pkt_r_rs2__8_, dispatch_pkt_r_rs2__7_, dispatch_pkt_r_rs2__6_, dispatch_pkt_r_rs2__5_, dispatch_pkt_r_rs2__4_, dispatch_pkt_r_rs2__3_, dispatch_pkt_r_rs2__2_, dispatch_pkt_r_rs2__1_, dispatch_pkt_r_rs2__0_ }),
    .data_o(pipe_fp_data_lo)
  );


  bsg_dff_width_p600
  calc_stage_reg
  (
    .clk_i(clk_i),
    .data_i({ calc_stage_r_3__instr_metadata__itag__7_, calc_stage_r_3__instr_metadata__itag__6_, calc_stage_r_3__instr_metadata__itag__5_, calc_stage_r_3__instr_metadata__itag__4_, calc_stage_r_3__instr_metadata__itag__3_, calc_stage_r_3__instr_metadata__itag__2_, calc_stage_r_3__instr_metadata__itag__1_, calc_stage_r_3__instr_metadata__itag__0_, calc_stage_r_3__instr_metadata__pc__63_, calc_stage_r_3__instr_metadata__pc__62_, calc_stage_r_3__instr_metadata__pc__61_, calc_stage_r_3__instr_metadata__pc__60_, calc_stage_r_3__instr_metadata__pc__59_, calc_stage_r_3__instr_metadata__pc__58_, calc_stage_r_3__instr_metadata__pc__57_, calc_stage_r_3__instr_metadata__pc__56_, calc_stage_r_3__instr_metadata__pc__55_, calc_stage_r_3__instr_metadata__pc__54_, calc_stage_r_3__instr_metadata__pc__53_, calc_stage_r_3__instr_metadata__pc__52_, calc_stage_r_3__instr_metadata__pc__51_, calc_stage_r_3__instr_metadata__pc__50_, calc_stage_r_3__instr_metadata__pc__49_, calc_stage_r_3__instr_metadata__pc__48_, calc_stage_r_3__instr_metadata__pc__47_, calc_stage_r_3__instr_metadata__pc__46_, calc_stage_r_3__instr_metadata__pc__45_, calc_stage_r_3__instr_metadata__pc__44_, calc_stage_r_3__instr_metadata__pc__43_, calc_stage_r_3__instr_metadata__pc__42_, calc_stage_r_3__instr_metadata__pc__41_, calc_stage_r_3__instr_metadata__pc__40_, calc_stage_r_3__instr_metadata__pc__39_, calc_stage_r_3__instr_metadata__pc__38_, calc_stage_r_3__instr_metadata__pc__37_, calc_stage_r_3__instr_metadata__pc__36_, calc_stage_r_3__instr_metadata__pc__35_, calc_stage_r_3__instr_metadata__pc__34_, calc_stage_r_3__instr_metadata__pc__33_, calc_stage_r_3__instr_metadata__pc__32_, calc_stage_r_3__instr_metadata__pc__31_, calc_stage_r_3__instr_metadata__pc__30_, calc_stage_r_3__instr_metadata__pc__29_, calc_stage_r_3__instr_metadata__pc__28_, calc_stage_r_3__instr_metadata__pc__27_, calc_stage_r_3__instr_metadata__pc__26_, calc_stage_r_3__instr_metadata__pc__25_, calc_stage_r_3__instr_metadata__pc__24_, calc_stage_r_3__instr_metadata__pc__23_, calc_stage_r_3__instr_metadata__pc__22_, calc_stage_r_3__instr_metadata__pc__21_, calc_stage_r_3__instr_metadata__pc__20_, calc_stage_r_3__instr_metadata__pc__19_, calc_stage_r_3__instr_metadata__pc__18_, calc_stage_r_3__instr_metadata__pc__17_, calc_stage_r_3__instr_metadata__pc__16_, calc_stage_r_3__instr_metadata__pc__15_, calc_stage_r_3__instr_metadata__pc__14_, calc_stage_r_3__instr_metadata__pc__13_, calc_stage_r_3__instr_metadata__pc__12_, calc_stage_r_3__instr_metadata__pc__11_, calc_stage_r_3__instr_metadata__pc__10_, calc_stage_r_3__instr_metadata__pc__9_, calc_stage_r_3__instr_metadata__pc__8_, calc_stage_r_3__instr_metadata__pc__7_, calc_stage_r_3__instr_metadata__pc__6_, calc_stage_r_3__instr_metadata__pc__5_, calc_stage_r_3__instr_metadata__pc__4_, calc_stage_r_3__instr_metadata__pc__3_, calc_stage_r_3__instr_metadata__pc__2_, calc_stage_r_3__instr_metadata__pc__1_, calc_stage_r_3__instr_metadata__pc__0_, calc_stage_r_3__instr_metadata__fe_exception_not_instr_, calc_stage_r_3__instr_metadata__fe_exception_code__1_, calc_stage_r_3__instr_metadata__fe_exception_code__0_, calc_stage_r_3__instr__31_, calc_stage_r_3__instr__30_, calc_stage_r_3__instr__29_, calc_stage_r_3__instr__28_, calc_stage_r_3__instr__27_, calc_stage_r_3__instr__26_, calc_stage_r_3__instr__25_, calc_stage_r_3__instr__24_, calc_stage_r_3__instr__23_, calc_stage_r_3__instr__22_, calc_stage_r_3__instr__21_, calc_stage_r_3__instr__20_, calc_stage_r_3__instr__19_, calc_stage_r_3__instr__18_, calc_stage_r_3__instr__17_, calc_stage_r_3__instr__16_, calc_stage_r_3__instr__15_, calc_stage_r_3__instr__14_, calc_stage_r_3__instr__13_, calc_stage_r_3__instr__12_, calc_stage_r_3__instr__11_, calc_stage_r_3__instr__10_, calc_stage_r_3__instr__9_, calc_stage_r_3__instr__8_, calc_stage_r_3__instr__7_, calc_stage_r_3__instr__6_, calc_stage_r_3__instr__5_, calc_stage_r_3__instr__4_, calc_stage_r_3__instr__3_, calc_stage_r_3__instr__2_, calc_stage_r_3__instr__1_, calc_stage_r_3__instr__0_, calc_stage_r_3__instr_v_, calc_stage_r_3__pipe_comp_v_, calc_stage_r_3__pipe_int_v_, calc_stage_r_3__pipe_mul_v_, calc_stage_r_3__pipe_mem_v_, calc_stage_r_3__pipe_fp_v_, calc_stage_r_3__irf_w_v_, calc_stage_r_3__frf_w_v_, calc_status_o[106:102], calc_stage_r_2__instr_metadata__itag__7_, calc_stage_r_2__instr_metadata__itag__6_, calc_stage_r_2__instr_metadata__itag__5_, calc_stage_r_2__instr_metadata__itag__4_, calc_stage_r_2__instr_metadata__itag__3_, calc_stage_r_2__instr_metadata__itag__2_, calc_stage_r_2__instr_metadata__itag__1_, calc_stage_r_2__instr_metadata__itag__0_, calc_status_o[67:4], calc_stage_r_2__instr_metadata__fe_exception_not_instr_, calc_stage_r_2__instr_metadata__fe_exception_code__1_, calc_stage_r_2__instr_metadata__fe_exception_code__0_, calc_stage_r_2__instr__31_, calc_stage_r_2__instr__30_, calc_stage_r_2__instr__29_, calc_stage_r_2__instr__28_, calc_stage_r_2__instr__27_, calc_stage_r_2__instr__26_, calc_stage_r_2__instr__25_, calc_stage_r_2__instr__24_, calc_stage_r_2__instr__23_, calc_stage_r_2__instr__22_, calc_stage_r_2__instr__21_, calc_stage_r_2__instr__20_, calc_stage_r_2__instr__19_, calc_stage_r_2__instr__18_, calc_stage_r_2__instr__17_, calc_stage_r_2__instr__16_, calc_stage_r_2__instr__15_, calc_stage_r_2__instr__14_, calc_stage_r_2__instr__13_, calc_stage_r_2__instr__12_, calc_stage_r_2__instr__11_, calc_stage_r_2__instr__10_, calc_stage_r_2__instr__9_, calc_stage_r_2__instr__8_, calc_stage_r_2__instr__7_, calc_stage_r_2__instr__6_, calc_stage_r_2__instr__5_, calc_stage_r_2__instr__4_, calc_stage_r_2__instr__3_, calc_stage_r_2__instr__2_, calc_stage_r_2__instr__1_, calc_stage_r_2__instr__0_, calc_stage_r_2__instr_v_, calc_stage_r_2__pipe_comp_v_, calc_stage_r_2__pipe_int_v_, calc_stage_r_2__pipe_mul_v_, calc_stage_r_2__pipe_mem_v_, calc_stage_r_2__pipe_fp_v_, calc_stage_r_2__irf_w_v_, calc_stage_r_2__frf_w_v_, calc_status_o[95:91], calc_stage_r_1__instr_metadata__itag__7_, calc_stage_r_1__instr_metadata__itag__6_, calc_stage_r_1__instr_metadata__itag__5_, calc_stage_r_1__instr_metadata__itag__4_, calc_stage_r_1__instr_metadata__itag__3_, calc_stage_r_1__instr_metadata__itag__2_, calc_stage_r_1__instr_metadata__itag__1_, calc_stage_r_1__instr_metadata__itag__0_, calc_stage_r_1__instr_metadata__pc__63_, calc_stage_r_1__instr_metadata__pc__62_, calc_stage_r_1__instr_metadata__pc__61_, calc_stage_r_1__instr_metadata__pc__60_, calc_stage_r_1__instr_metadata__pc__59_, calc_stage_r_1__instr_metadata__pc__58_, calc_stage_r_1__instr_metadata__pc__57_, calc_stage_r_1__instr_metadata__pc__56_, calc_stage_r_1__instr_metadata__pc__55_, calc_stage_r_1__instr_metadata__pc__54_, calc_stage_r_1__instr_metadata__pc__53_, calc_stage_r_1__instr_metadata__pc__52_, calc_stage_r_1__instr_metadata__pc__51_, calc_stage_r_1__instr_metadata__pc__50_, calc_stage_r_1__instr_metadata__pc__49_, calc_stage_r_1__instr_metadata__pc__48_, calc_stage_r_1__instr_metadata__pc__47_, calc_stage_r_1__instr_metadata__pc__46_, calc_stage_r_1__instr_metadata__pc__45_, calc_stage_r_1__instr_metadata__pc__44_, calc_stage_r_1__instr_metadata__pc__43_, calc_stage_r_1__instr_metadata__pc__42_, calc_stage_r_1__instr_metadata__pc__41_, calc_stage_r_1__instr_metadata__pc__40_, calc_stage_r_1__instr_metadata__pc__39_, calc_stage_r_1__instr_metadata__pc__38_, calc_stage_r_1__instr_metadata__pc__37_, calc_stage_r_1__instr_metadata__pc__36_, calc_stage_r_1__instr_metadata__pc__35_, calc_stage_r_1__instr_metadata__pc__34_, calc_stage_r_1__instr_metadata__pc__33_, calc_stage_r_1__instr_metadata__pc__32_, calc_stage_r_1__instr_metadata__pc__31_, calc_stage_r_1__instr_metadata__pc__30_, calc_stage_r_1__instr_metadata__pc__29_, calc_stage_r_1__instr_metadata__pc__28_, calc_stage_r_1__instr_metadata__pc__27_, calc_stage_r_1__instr_metadata__pc__26_, calc_stage_r_1__instr_metadata__pc__25_, calc_stage_r_1__instr_metadata__pc__24_, calc_stage_r_1__instr_metadata__pc__23_, calc_stage_r_1__instr_metadata__pc__22_, calc_stage_r_1__instr_metadata__pc__21_, calc_stage_r_1__instr_metadata__pc__20_, calc_stage_r_1__instr_metadata__pc__19_, calc_stage_r_1__instr_metadata__pc__18_, calc_stage_r_1__instr_metadata__pc__17_, calc_stage_r_1__instr_metadata__pc__16_, calc_stage_r_1__instr_metadata__pc__15_, calc_stage_r_1__instr_metadata__pc__14_, calc_stage_r_1__instr_metadata__pc__13_, calc_stage_r_1__instr_metadata__pc__12_, calc_stage_r_1__instr_metadata__pc__11_, calc_stage_r_1__instr_metadata__pc__10_, calc_stage_r_1__instr_metadata__pc__9_, calc_stage_r_1__instr_metadata__pc__8_, calc_stage_r_1__instr_metadata__pc__7_, calc_stage_r_1__instr_metadata__pc__6_, calc_stage_r_1__instr_metadata__pc__5_, calc_stage_r_1__instr_metadata__pc__4_, calc_stage_r_1__instr_metadata__pc__3_, calc_stage_r_1__instr_metadata__pc__2_, calc_stage_r_1__instr_metadata__pc__1_, calc_stage_r_1__instr_metadata__pc__0_, calc_stage_r_1__instr_metadata__fe_exception_not_instr_, calc_stage_r_1__instr_metadata__fe_exception_code__1_, calc_stage_r_1__instr_metadata__fe_exception_code__0_, calc_stage_r_1__instr__31_, calc_stage_r_1__instr__30_, calc_stage_r_1__instr__29_, calc_stage_r_1__instr__28_, calc_stage_r_1__instr__27_, calc_stage_r_1__instr__26_, calc_stage_r_1__instr__25_, calc_stage_r_1__instr__24_, calc_stage_r_1__instr__23_, calc_stage_r_1__instr__22_, calc_stage_r_1__instr__21_, calc_stage_r_1__instr__20_, calc_stage_r_1__instr__19_, calc_stage_r_1__instr__18_, calc_stage_r_1__instr__17_, calc_stage_r_1__instr__16_, calc_stage_r_1__instr__15_, calc_stage_r_1__instr__14_, calc_stage_r_1__instr__13_, calc_stage_r_1__instr__12_, calc_stage_r_1__instr__11_, calc_stage_r_1__instr__10_, calc_stage_r_1__instr__9_, calc_stage_r_1__instr__8_, calc_stage_r_1__instr__7_, calc_stage_r_1__instr__6_, calc_stage_r_1__instr__5_, calc_stage_r_1__instr__4_, calc_stage_r_1__instr__3_, calc_stage_r_1__instr__2_, calc_stage_r_1__instr__1_, calc_stage_r_1__instr__0_, calc_stage_r_1__instr_v_, calc_stage_r_1__pipe_comp_v_, calc_stage_r_1__pipe_int_v_, calc_stage_r_1__pipe_mul_v_, calc_stage_r_1__pipe_mem_v_, calc_stage_r_1__pipe_fp_v_, calc_stage_r_1__irf_w_v_, calc_stage_r_1__frf_w_v_, calc_status_o[84:80], calc_stage_r_0__instr_metadata__itag__7_, calc_stage_r_0__instr_metadata__itag__6_, calc_stage_r_0__instr_metadata__itag__5_, calc_stage_r_0__instr_metadata__itag__4_, calc_stage_r_0__instr_metadata__itag__3_, calc_stage_r_0__instr_metadata__itag__2_, calc_stage_r_0__instr_metadata__itag__1_, calc_stage_r_0__instr_metadata__itag__0_, calc_stage_r_0__instr_metadata__pc__63_, calc_stage_r_0__instr_metadata__pc__62_, calc_stage_r_0__instr_metadata__pc__61_, calc_stage_r_0__instr_metadata__pc__60_, calc_stage_r_0__instr_metadata__pc__59_, calc_stage_r_0__instr_metadata__pc__58_, calc_stage_r_0__instr_metadata__pc__57_, calc_stage_r_0__instr_metadata__pc__56_, calc_stage_r_0__instr_metadata__pc__55_, calc_stage_r_0__instr_metadata__pc__54_, calc_stage_r_0__instr_metadata__pc__53_, calc_stage_r_0__instr_metadata__pc__52_, calc_stage_r_0__instr_metadata__pc__51_, calc_stage_r_0__instr_metadata__pc__50_, calc_stage_r_0__instr_metadata__pc__49_, calc_stage_r_0__instr_metadata__pc__48_, calc_stage_r_0__instr_metadata__pc__47_, calc_stage_r_0__instr_metadata__pc__46_, calc_stage_r_0__instr_metadata__pc__45_, calc_stage_r_0__instr_metadata__pc__44_, calc_stage_r_0__instr_metadata__pc__43_, calc_stage_r_0__instr_metadata__pc__42_, calc_stage_r_0__instr_metadata__pc__41_, calc_stage_r_0__instr_metadata__pc__40_, calc_stage_r_0__instr_metadata__pc__39_, calc_stage_r_0__instr_metadata__pc__38_, calc_stage_r_0__instr_metadata__pc__37_, calc_stage_r_0__instr_metadata__pc__36_, calc_stage_r_0__instr_metadata__pc__35_, calc_stage_r_0__instr_metadata__pc__34_, calc_stage_r_0__instr_metadata__pc__33_, calc_stage_r_0__instr_metadata__pc__32_, calc_stage_r_0__instr_metadata__pc__31_, calc_stage_r_0__instr_metadata__pc__30_, calc_stage_r_0__instr_metadata__pc__29_, calc_stage_r_0__instr_metadata__pc__28_, calc_stage_r_0__instr_metadata__pc__27_, calc_stage_r_0__instr_metadata__pc__26_, calc_stage_r_0__instr_metadata__pc__25_, calc_stage_r_0__instr_metadata__pc__24_, calc_stage_r_0__instr_metadata__pc__23_, calc_stage_r_0__instr_metadata__pc__22_, calc_stage_r_0__instr_metadata__pc__21_, calc_stage_r_0__instr_metadata__pc__20_, calc_stage_r_0__instr_metadata__pc__19_, calc_stage_r_0__instr_metadata__pc__18_, calc_stage_r_0__instr_metadata__pc__17_, calc_stage_r_0__instr_metadata__pc__16_, calc_stage_r_0__instr_metadata__pc__15_, calc_stage_r_0__instr_metadata__pc__14_, calc_stage_r_0__instr_metadata__pc__13_, calc_stage_r_0__instr_metadata__pc__12_, calc_stage_r_0__instr_metadata__pc__11_, calc_stage_r_0__instr_metadata__pc__10_, calc_stage_r_0__instr_metadata__pc__9_, calc_stage_r_0__instr_metadata__pc__8_, calc_stage_r_0__instr_metadata__pc__7_, calc_stage_r_0__instr_metadata__pc__6_, calc_stage_r_0__instr_metadata__pc__5_, calc_stage_r_0__instr_metadata__pc__4_, calc_stage_r_0__instr_metadata__pc__3_, calc_stage_r_0__instr_metadata__pc__2_, calc_stage_r_0__instr_metadata__pc__1_, calc_stage_r_0__instr_metadata__pc__0_, calc_stage_r_0__instr_metadata__fe_exception_not_instr_, calc_stage_r_0__instr_metadata__fe_exception_code__1_, calc_stage_r_0__instr_metadata__fe_exception_code__0_, calc_stage_r_0__instr__31_, calc_stage_r_0__instr__30_, calc_stage_r_0__instr__29_, calc_stage_r_0__instr__28_, calc_stage_r_0__instr__27_, calc_stage_r_0__instr__26_, calc_stage_r_0__instr__25_, calc_stage_r_0__instr__24_, calc_stage_r_0__instr__23_, calc_stage_r_0__instr__22_, calc_stage_r_0__instr__21_, calc_stage_r_0__instr__20_, calc_stage_r_0__instr__19_, calc_stage_r_0__instr__18_, calc_stage_r_0__instr__17_, calc_stage_r_0__instr__16_, calc_stage_r_0__instr__15_, calc_stage_r_0__instr__14_, calc_stage_r_0__instr__13_, calc_stage_r_0__instr__12_, calc_stage_r_0__instr__11_, calc_stage_r_0__instr__10_, calc_stage_r_0__instr__9_, calc_stage_r_0__instr__8_, calc_stage_r_0__instr__7_, calc_stage_r_0__instr__6_, calc_stage_r_0__instr__5_, calc_stage_r_0__instr__4_, calc_stage_r_0__instr__3_, calc_stage_r_0__instr__2_, calc_stage_r_0__instr__1_, calc_stage_r_0__instr__0_, calc_stage_r_0__instr_v_, calc_stage_r_0__pipe_comp_v_, calc_stage_r_0__pipe_int_v_, calc_stage_r_0__pipe_mul_v_, calc_stage_r_0__pipe_mem_v_, calc_stage_r_0__pipe_fp_v_, calc_stage_r_0__irf_w_v_, calc_stage_r_0__frf_w_v_, calc_status_o[73:69], dispatch_pkt[385:311], dispatch_pkt[274:242], dispatch_pkt[238:232], dispatch_pkt[200:196] }),
    .data_o({ calc_stage_r_4__instr_metadata__itag__7_, calc_stage_r_4__instr_metadata__itag__6_, calc_stage_r_4__instr_metadata__itag__5_, calc_stage_r_4__instr_metadata__itag__4_, calc_stage_r_4__instr_metadata__itag__3_, calc_stage_r_4__instr_metadata__itag__2_, calc_stage_r_4__instr_metadata__itag__1_, calc_stage_r_4__instr_metadata__itag__0_, calc_stage_r_4__instr_metadata__pc__63_, calc_stage_r_4__instr_metadata__pc__62_, calc_stage_r_4__instr_metadata__pc__61_, calc_stage_r_4__instr_metadata__pc__60_, calc_stage_r_4__instr_metadata__pc__59_, calc_stage_r_4__instr_metadata__pc__58_, calc_stage_r_4__instr_metadata__pc__57_, calc_stage_r_4__instr_metadata__pc__56_, calc_stage_r_4__instr_metadata__pc__55_, calc_stage_r_4__instr_metadata__pc__54_, calc_stage_r_4__instr_metadata__pc__53_, calc_stage_r_4__instr_metadata__pc__52_, calc_stage_r_4__instr_metadata__pc__51_, calc_stage_r_4__instr_metadata__pc__50_, calc_stage_r_4__instr_metadata__pc__49_, calc_stage_r_4__instr_metadata__pc__48_, calc_stage_r_4__instr_metadata__pc__47_, calc_stage_r_4__instr_metadata__pc__46_, calc_stage_r_4__instr_metadata__pc__45_, calc_stage_r_4__instr_metadata__pc__44_, calc_stage_r_4__instr_metadata__pc__43_, calc_stage_r_4__instr_metadata__pc__42_, calc_stage_r_4__instr_metadata__pc__41_, calc_stage_r_4__instr_metadata__pc__40_, calc_stage_r_4__instr_metadata__pc__39_, calc_stage_r_4__instr_metadata__pc__38_, calc_stage_r_4__instr_metadata__pc__37_, calc_stage_r_4__instr_metadata__pc__36_, calc_stage_r_4__instr_metadata__pc__35_, calc_stage_r_4__instr_metadata__pc__34_, calc_stage_r_4__instr_metadata__pc__33_, calc_stage_r_4__instr_metadata__pc__32_, calc_stage_r_4__instr_metadata__pc__31_, calc_stage_r_4__instr_metadata__pc__30_, calc_stage_r_4__instr_metadata__pc__29_, calc_stage_r_4__instr_metadata__pc__28_, calc_stage_r_4__instr_metadata__pc__27_, calc_stage_r_4__instr_metadata__pc__26_, calc_stage_r_4__instr_metadata__pc__25_, calc_stage_r_4__instr_metadata__pc__24_, calc_stage_r_4__instr_metadata__pc__23_, calc_stage_r_4__instr_metadata__pc__22_, calc_stage_r_4__instr_metadata__pc__21_, calc_stage_r_4__instr_metadata__pc__20_, calc_stage_r_4__instr_metadata__pc__19_, calc_stage_r_4__instr_metadata__pc__18_, calc_stage_r_4__instr_metadata__pc__17_, calc_stage_r_4__instr_metadata__pc__16_, calc_stage_r_4__instr_metadata__pc__15_, calc_stage_r_4__instr_metadata__pc__14_, calc_stage_r_4__instr_metadata__pc__13_, calc_stage_r_4__instr_metadata__pc__12_, calc_stage_r_4__instr_metadata__pc__11_, calc_stage_r_4__instr_metadata__pc__10_, calc_stage_r_4__instr_metadata__pc__9_, calc_stage_r_4__instr_metadata__pc__8_, calc_stage_r_4__instr_metadata__pc__7_, calc_stage_r_4__instr_metadata__pc__6_, calc_stage_r_4__instr_metadata__pc__5_, calc_stage_r_4__instr_metadata__pc__4_, calc_stage_r_4__instr_metadata__pc__3_, calc_stage_r_4__instr_metadata__pc__2_, calc_stage_r_4__instr_metadata__pc__1_, calc_stage_r_4__instr_metadata__pc__0_, calc_stage_r_4__instr_metadata__fe_exception_not_instr_, calc_stage_r_4__instr_metadata__fe_exception_code__1_, calc_stage_r_4__instr_metadata__fe_exception_code__0_, calc_stage_r_4__instr__31_, calc_stage_r_4__instr__30_, calc_stage_r_4__instr__29_, calc_stage_r_4__instr__28_, calc_stage_r_4__instr__27_, calc_stage_r_4__instr__26_, calc_stage_r_4__instr__25_, calc_stage_r_4__instr__24_, calc_stage_r_4__instr__23_, calc_stage_r_4__instr__22_, calc_stage_r_4__instr__21_, calc_stage_r_4__instr__20_, calc_stage_r_4__instr__19_, calc_stage_r_4__instr__18_, calc_stage_r_4__instr__17_, calc_stage_r_4__instr__16_, calc_stage_r_4__instr__15_, calc_stage_r_4__instr__14_, calc_stage_r_4__instr__13_, calc_stage_r_4__instr__12_, calc_stage_r_4__instr__11_, calc_stage_r_4__instr__10_, calc_stage_r_4__instr__9_, calc_stage_r_4__instr__8_, calc_stage_r_4__instr__7_, calc_stage_r_4__instr__6_, calc_stage_r_4__instr__5_, calc_stage_r_4__instr__4_, calc_stage_r_4__instr__3_, calc_stage_r_4__instr__2_, calc_stage_r_4__instr__1_, calc_stage_r_4__instr__0_, calc_stage_r_4__instr_v_, calc_stage_r_4__pipe_comp_v_, calc_stage_r_4__pipe_int_v_, calc_stage_r_4__pipe_mul_v_, calc_stage_r_4__pipe_mem_v_, calc_stage_r_4__pipe_fp_v_, calc_stage_r_4__irf_w_v_, calc_stage_r_4__frf_w_v_, calc_status_o[117:113], calc_stage_r_3__instr_metadata__itag__7_, calc_stage_r_3__instr_metadata__itag__6_, calc_stage_r_3__instr_metadata__itag__5_, calc_stage_r_3__instr_metadata__itag__4_, calc_stage_r_3__instr_metadata__itag__3_, calc_stage_r_3__instr_metadata__itag__2_, calc_stage_r_3__instr_metadata__itag__1_, calc_stage_r_3__instr_metadata__itag__0_, calc_stage_r_3__instr_metadata__pc__63_, calc_stage_r_3__instr_metadata__pc__62_, calc_stage_r_3__instr_metadata__pc__61_, calc_stage_r_3__instr_metadata__pc__60_, calc_stage_r_3__instr_metadata__pc__59_, calc_stage_r_3__instr_metadata__pc__58_, calc_stage_r_3__instr_metadata__pc__57_, calc_stage_r_3__instr_metadata__pc__56_, calc_stage_r_3__instr_metadata__pc__55_, calc_stage_r_3__instr_metadata__pc__54_, calc_stage_r_3__instr_metadata__pc__53_, calc_stage_r_3__instr_metadata__pc__52_, calc_stage_r_3__instr_metadata__pc__51_, calc_stage_r_3__instr_metadata__pc__50_, calc_stage_r_3__instr_metadata__pc__49_, calc_stage_r_3__instr_metadata__pc__48_, calc_stage_r_3__instr_metadata__pc__47_, calc_stage_r_3__instr_metadata__pc__46_, calc_stage_r_3__instr_metadata__pc__45_, calc_stage_r_3__instr_metadata__pc__44_, calc_stage_r_3__instr_metadata__pc__43_, calc_stage_r_3__instr_metadata__pc__42_, calc_stage_r_3__instr_metadata__pc__41_, calc_stage_r_3__instr_metadata__pc__40_, calc_stage_r_3__instr_metadata__pc__39_, calc_stage_r_3__instr_metadata__pc__38_, calc_stage_r_3__instr_metadata__pc__37_, calc_stage_r_3__instr_metadata__pc__36_, calc_stage_r_3__instr_metadata__pc__35_, calc_stage_r_3__instr_metadata__pc__34_, calc_stage_r_3__instr_metadata__pc__33_, calc_stage_r_3__instr_metadata__pc__32_, calc_stage_r_3__instr_metadata__pc__31_, calc_stage_r_3__instr_metadata__pc__30_, calc_stage_r_3__instr_metadata__pc__29_, calc_stage_r_3__instr_metadata__pc__28_, calc_stage_r_3__instr_metadata__pc__27_, calc_stage_r_3__instr_metadata__pc__26_, calc_stage_r_3__instr_metadata__pc__25_, calc_stage_r_3__instr_metadata__pc__24_, calc_stage_r_3__instr_metadata__pc__23_, calc_stage_r_3__instr_metadata__pc__22_, calc_stage_r_3__instr_metadata__pc__21_, calc_stage_r_3__instr_metadata__pc__20_, calc_stage_r_3__instr_metadata__pc__19_, calc_stage_r_3__instr_metadata__pc__18_, calc_stage_r_3__instr_metadata__pc__17_, calc_stage_r_3__instr_metadata__pc__16_, calc_stage_r_3__instr_metadata__pc__15_, calc_stage_r_3__instr_metadata__pc__14_, calc_stage_r_3__instr_metadata__pc__13_, calc_stage_r_3__instr_metadata__pc__12_, calc_stage_r_3__instr_metadata__pc__11_, calc_stage_r_3__instr_metadata__pc__10_, calc_stage_r_3__instr_metadata__pc__9_, calc_stage_r_3__instr_metadata__pc__8_, calc_stage_r_3__instr_metadata__pc__7_, calc_stage_r_3__instr_metadata__pc__6_, calc_stage_r_3__instr_metadata__pc__5_, calc_stage_r_3__instr_metadata__pc__4_, calc_stage_r_3__instr_metadata__pc__3_, calc_stage_r_3__instr_metadata__pc__2_, calc_stage_r_3__instr_metadata__pc__1_, calc_stage_r_3__instr_metadata__pc__0_, calc_stage_r_3__instr_metadata__fe_exception_not_instr_, calc_stage_r_3__instr_metadata__fe_exception_code__1_, calc_stage_r_3__instr_metadata__fe_exception_code__0_, calc_stage_r_3__instr__31_, calc_stage_r_3__instr__30_, calc_stage_r_3__instr__29_, calc_stage_r_3__instr__28_, calc_stage_r_3__instr__27_, calc_stage_r_3__instr__26_, calc_stage_r_3__instr__25_, calc_stage_r_3__instr__24_, calc_stage_r_3__instr__23_, calc_stage_r_3__instr__22_, calc_stage_r_3__instr__21_, calc_stage_r_3__instr__20_, calc_stage_r_3__instr__19_, calc_stage_r_3__instr__18_, calc_stage_r_3__instr__17_, calc_stage_r_3__instr__16_, calc_stage_r_3__instr__15_, calc_stage_r_3__instr__14_, calc_stage_r_3__instr__13_, calc_stage_r_3__instr__12_, calc_stage_r_3__instr__11_, calc_stage_r_3__instr__10_, calc_stage_r_3__instr__9_, calc_stage_r_3__instr__8_, calc_stage_r_3__instr__7_, calc_stage_r_3__instr__6_, calc_stage_r_3__instr__5_, calc_stage_r_3__instr__4_, calc_stage_r_3__instr__3_, calc_stage_r_3__instr__2_, calc_stage_r_3__instr__1_, calc_stage_r_3__instr__0_, calc_stage_r_3__instr_v_, calc_stage_r_3__pipe_comp_v_, calc_stage_r_3__pipe_int_v_, calc_stage_r_3__pipe_mul_v_, calc_stage_r_3__pipe_mem_v_, calc_stage_r_3__pipe_fp_v_, calc_stage_r_3__irf_w_v_, calc_stage_r_3__frf_w_v_, calc_status_o[106:102], calc_stage_r_2__instr_metadata__itag__7_, calc_stage_r_2__instr_metadata__itag__6_, calc_stage_r_2__instr_metadata__itag__5_, calc_stage_r_2__instr_metadata__itag__4_, calc_stage_r_2__instr_metadata__itag__3_, calc_stage_r_2__instr_metadata__itag__2_, calc_stage_r_2__instr_metadata__itag__1_, calc_stage_r_2__instr_metadata__itag__0_, calc_status_o[67:4], calc_stage_r_2__instr_metadata__fe_exception_not_instr_, calc_stage_r_2__instr_metadata__fe_exception_code__1_, calc_stage_r_2__instr_metadata__fe_exception_code__0_, calc_stage_r_2__instr__31_, calc_stage_r_2__instr__30_, calc_stage_r_2__instr__29_, calc_stage_r_2__instr__28_, calc_stage_r_2__instr__27_, calc_stage_r_2__instr__26_, calc_stage_r_2__instr__25_, calc_stage_r_2__instr__24_, calc_stage_r_2__instr__23_, calc_stage_r_2__instr__22_, calc_stage_r_2__instr__21_, calc_stage_r_2__instr__20_, calc_stage_r_2__instr__19_, calc_stage_r_2__instr__18_, calc_stage_r_2__instr__17_, calc_stage_r_2__instr__16_, calc_stage_r_2__instr__15_, calc_stage_r_2__instr__14_, calc_stage_r_2__instr__13_, calc_stage_r_2__instr__12_, calc_stage_r_2__instr__11_, calc_stage_r_2__instr__10_, calc_stage_r_2__instr__9_, calc_stage_r_2__instr__8_, calc_stage_r_2__instr__7_, calc_stage_r_2__instr__6_, calc_stage_r_2__instr__5_, calc_stage_r_2__instr__4_, calc_stage_r_2__instr__3_, calc_stage_r_2__instr__2_, calc_stage_r_2__instr__1_, calc_stage_r_2__instr__0_, calc_stage_r_2__instr_v_, calc_stage_r_2__pipe_comp_v_, calc_stage_r_2__pipe_int_v_, calc_stage_r_2__pipe_mul_v_, calc_stage_r_2__pipe_mem_v_, calc_stage_r_2__pipe_fp_v_, calc_stage_r_2__irf_w_v_, calc_stage_r_2__frf_w_v_, calc_status_o[95:91], calc_stage_r_1__instr_metadata__itag__7_, calc_stage_r_1__instr_metadata__itag__6_, calc_stage_r_1__instr_metadata__itag__5_, calc_stage_r_1__instr_metadata__itag__4_, calc_stage_r_1__instr_metadata__itag__3_, calc_stage_r_1__instr_metadata__itag__2_, calc_stage_r_1__instr_metadata__itag__1_, calc_stage_r_1__instr_metadata__itag__0_, calc_stage_r_1__instr_metadata__pc__63_, calc_stage_r_1__instr_metadata__pc__62_, calc_stage_r_1__instr_metadata__pc__61_, calc_stage_r_1__instr_metadata__pc__60_, calc_stage_r_1__instr_metadata__pc__59_, calc_stage_r_1__instr_metadata__pc__58_, calc_stage_r_1__instr_metadata__pc__57_, calc_stage_r_1__instr_metadata__pc__56_, calc_stage_r_1__instr_metadata__pc__55_, calc_stage_r_1__instr_metadata__pc__54_, calc_stage_r_1__instr_metadata__pc__53_, calc_stage_r_1__instr_metadata__pc__52_, calc_stage_r_1__instr_metadata__pc__51_, calc_stage_r_1__instr_metadata__pc__50_, calc_stage_r_1__instr_metadata__pc__49_, calc_stage_r_1__instr_metadata__pc__48_, calc_stage_r_1__instr_metadata__pc__47_, calc_stage_r_1__instr_metadata__pc__46_, calc_stage_r_1__instr_metadata__pc__45_, calc_stage_r_1__instr_metadata__pc__44_, calc_stage_r_1__instr_metadata__pc__43_, calc_stage_r_1__instr_metadata__pc__42_, calc_stage_r_1__instr_metadata__pc__41_, calc_stage_r_1__instr_metadata__pc__40_, calc_stage_r_1__instr_metadata__pc__39_, calc_stage_r_1__instr_metadata__pc__38_, calc_stage_r_1__instr_metadata__pc__37_, calc_stage_r_1__instr_metadata__pc__36_, calc_stage_r_1__instr_metadata__pc__35_, calc_stage_r_1__instr_metadata__pc__34_, calc_stage_r_1__instr_metadata__pc__33_, calc_stage_r_1__instr_metadata__pc__32_, calc_stage_r_1__instr_metadata__pc__31_, calc_stage_r_1__instr_metadata__pc__30_, calc_stage_r_1__instr_metadata__pc__29_, calc_stage_r_1__instr_metadata__pc__28_, calc_stage_r_1__instr_metadata__pc__27_, calc_stage_r_1__instr_metadata__pc__26_, calc_stage_r_1__instr_metadata__pc__25_, calc_stage_r_1__instr_metadata__pc__24_, calc_stage_r_1__instr_metadata__pc__23_, calc_stage_r_1__instr_metadata__pc__22_, calc_stage_r_1__instr_metadata__pc__21_, calc_stage_r_1__instr_metadata__pc__20_, calc_stage_r_1__instr_metadata__pc__19_, calc_stage_r_1__instr_metadata__pc__18_, calc_stage_r_1__instr_metadata__pc__17_, calc_stage_r_1__instr_metadata__pc__16_, calc_stage_r_1__instr_metadata__pc__15_, calc_stage_r_1__instr_metadata__pc__14_, calc_stage_r_1__instr_metadata__pc__13_, calc_stage_r_1__instr_metadata__pc__12_, calc_stage_r_1__instr_metadata__pc__11_, calc_stage_r_1__instr_metadata__pc__10_, calc_stage_r_1__instr_metadata__pc__9_, calc_stage_r_1__instr_metadata__pc__8_, calc_stage_r_1__instr_metadata__pc__7_, calc_stage_r_1__instr_metadata__pc__6_, calc_stage_r_1__instr_metadata__pc__5_, calc_stage_r_1__instr_metadata__pc__4_, calc_stage_r_1__instr_metadata__pc__3_, calc_stage_r_1__instr_metadata__pc__2_, calc_stage_r_1__instr_metadata__pc__1_, calc_stage_r_1__instr_metadata__pc__0_, calc_stage_r_1__instr_metadata__fe_exception_not_instr_, calc_stage_r_1__instr_metadata__fe_exception_code__1_, calc_stage_r_1__instr_metadata__fe_exception_code__0_, calc_stage_r_1__instr__31_, calc_stage_r_1__instr__30_, calc_stage_r_1__instr__29_, calc_stage_r_1__instr__28_, calc_stage_r_1__instr__27_, calc_stage_r_1__instr__26_, calc_stage_r_1__instr__25_, calc_stage_r_1__instr__24_, calc_stage_r_1__instr__23_, calc_stage_r_1__instr__22_, calc_stage_r_1__instr__21_, calc_stage_r_1__instr__20_, calc_stage_r_1__instr__19_, calc_stage_r_1__instr__18_, calc_stage_r_1__instr__17_, calc_stage_r_1__instr__16_, calc_stage_r_1__instr__15_, calc_stage_r_1__instr__14_, calc_stage_r_1__instr__13_, calc_stage_r_1__instr__12_, calc_stage_r_1__instr__11_, calc_stage_r_1__instr__10_, calc_stage_r_1__instr__9_, calc_stage_r_1__instr__8_, calc_stage_r_1__instr__7_, calc_stage_r_1__instr__6_, calc_stage_r_1__instr__5_, calc_stage_r_1__instr__4_, calc_stage_r_1__instr__3_, calc_stage_r_1__instr__2_, calc_stage_r_1__instr__1_, calc_stage_r_1__instr__0_, calc_stage_r_1__instr_v_, calc_stage_r_1__pipe_comp_v_, calc_stage_r_1__pipe_int_v_, calc_stage_r_1__pipe_mul_v_, calc_stage_r_1__pipe_mem_v_, calc_stage_r_1__pipe_fp_v_, calc_stage_r_1__irf_w_v_, calc_stage_r_1__frf_w_v_, calc_status_o[84:80], calc_stage_r_0__instr_metadata__itag__7_, calc_stage_r_0__instr_metadata__itag__6_, calc_stage_r_0__instr_metadata__itag__5_, calc_stage_r_0__instr_metadata__itag__4_, calc_stage_r_0__instr_metadata__itag__3_, calc_stage_r_0__instr_metadata__itag__2_, calc_stage_r_0__instr_metadata__itag__1_, calc_stage_r_0__instr_metadata__itag__0_, calc_stage_r_0__instr_metadata__pc__63_, calc_stage_r_0__instr_metadata__pc__62_, calc_stage_r_0__instr_metadata__pc__61_, calc_stage_r_0__instr_metadata__pc__60_, calc_stage_r_0__instr_metadata__pc__59_, calc_stage_r_0__instr_metadata__pc__58_, calc_stage_r_0__instr_metadata__pc__57_, calc_stage_r_0__instr_metadata__pc__56_, calc_stage_r_0__instr_metadata__pc__55_, calc_stage_r_0__instr_metadata__pc__54_, calc_stage_r_0__instr_metadata__pc__53_, calc_stage_r_0__instr_metadata__pc__52_, calc_stage_r_0__instr_metadata__pc__51_, calc_stage_r_0__instr_metadata__pc__50_, calc_stage_r_0__instr_metadata__pc__49_, calc_stage_r_0__instr_metadata__pc__48_, calc_stage_r_0__instr_metadata__pc__47_, calc_stage_r_0__instr_metadata__pc__46_, calc_stage_r_0__instr_metadata__pc__45_, calc_stage_r_0__instr_metadata__pc__44_, calc_stage_r_0__instr_metadata__pc__43_, calc_stage_r_0__instr_metadata__pc__42_, calc_stage_r_0__instr_metadata__pc__41_, calc_stage_r_0__instr_metadata__pc__40_, calc_stage_r_0__instr_metadata__pc__39_, calc_stage_r_0__instr_metadata__pc__38_, calc_stage_r_0__instr_metadata__pc__37_, calc_stage_r_0__instr_metadata__pc__36_, calc_stage_r_0__instr_metadata__pc__35_, calc_stage_r_0__instr_metadata__pc__34_, calc_stage_r_0__instr_metadata__pc__33_, calc_stage_r_0__instr_metadata__pc__32_, calc_stage_r_0__instr_metadata__pc__31_, calc_stage_r_0__instr_metadata__pc__30_, calc_stage_r_0__instr_metadata__pc__29_, calc_stage_r_0__instr_metadata__pc__28_, calc_stage_r_0__instr_metadata__pc__27_, calc_stage_r_0__instr_metadata__pc__26_, calc_stage_r_0__instr_metadata__pc__25_, calc_stage_r_0__instr_metadata__pc__24_, calc_stage_r_0__instr_metadata__pc__23_, calc_stage_r_0__instr_metadata__pc__22_, calc_stage_r_0__instr_metadata__pc__21_, calc_stage_r_0__instr_metadata__pc__20_, calc_stage_r_0__instr_metadata__pc__19_, calc_stage_r_0__instr_metadata__pc__18_, calc_stage_r_0__instr_metadata__pc__17_, calc_stage_r_0__instr_metadata__pc__16_, calc_stage_r_0__instr_metadata__pc__15_, calc_stage_r_0__instr_metadata__pc__14_, calc_stage_r_0__instr_metadata__pc__13_, calc_stage_r_0__instr_metadata__pc__12_, calc_stage_r_0__instr_metadata__pc__11_, calc_stage_r_0__instr_metadata__pc__10_, calc_stage_r_0__instr_metadata__pc__9_, calc_stage_r_0__instr_metadata__pc__8_, calc_stage_r_0__instr_metadata__pc__7_, calc_stage_r_0__instr_metadata__pc__6_, calc_stage_r_0__instr_metadata__pc__5_, calc_stage_r_0__instr_metadata__pc__4_, calc_stage_r_0__instr_metadata__pc__3_, calc_stage_r_0__instr_metadata__pc__2_, calc_stage_r_0__instr_metadata__pc__1_, calc_stage_r_0__instr_metadata__pc__0_, calc_stage_r_0__instr_metadata__fe_exception_not_instr_, calc_stage_r_0__instr_metadata__fe_exception_code__1_, calc_stage_r_0__instr_metadata__fe_exception_code__0_, calc_stage_r_0__instr__31_, calc_stage_r_0__instr__30_, calc_stage_r_0__instr__29_, calc_stage_r_0__instr__28_, calc_stage_r_0__instr__27_, calc_stage_r_0__instr__26_, calc_stage_r_0__instr__25_, calc_stage_r_0__instr__24_, calc_stage_r_0__instr__23_, calc_stage_r_0__instr__22_, calc_stage_r_0__instr__21_, calc_stage_r_0__instr__20_, calc_stage_r_0__instr__19_, calc_stage_r_0__instr__18_, calc_stage_r_0__instr__17_, calc_stage_r_0__instr__16_, calc_stage_r_0__instr__15_, calc_stage_r_0__instr__14_, calc_stage_r_0__instr__13_, calc_stage_r_0__instr__12_, calc_stage_r_0__instr__11_, calc_stage_r_0__instr__10_, calc_stage_r_0__instr__9_, calc_stage_r_0__instr__8_, calc_stage_r_0__instr__7_, calc_stage_r_0__instr__6_, calc_stage_r_0__instr__5_, calc_stage_r_0__instr__4_, calc_stage_r_0__instr__3_, calc_stage_r_0__instr__2_, calc_stage_r_0__instr__1_, calc_stage_r_0__instr__0_, calc_stage_r_0__instr_v_, calc_stage_r_0__pipe_comp_v_, calc_stage_r_0__pipe_int_v_, calc_stage_r_0__pipe_mul_v_, calc_stage_r_0__pipe_mem_v_, calc_stage_r_0__pipe_fp_v_, calc_stage_r_0__irf_w_v_, calc_stage_r_0__frf_w_v_, calc_status_o[73:69] })
  );


  bsg_dff_width_p386
  dispatch_pkt_reg
  (
    .clk_i(clk_i),
    .data_i(dispatch_pkt),
    .data_o({ dispatch_pkt_r_instr_metadata__itag__7_, dispatch_pkt_r_instr_metadata__itag__6_, dispatch_pkt_r_instr_metadata__itag__5_, dispatch_pkt_r_instr_metadata__itag__4_, dispatch_pkt_r_instr_metadata__itag__3_, dispatch_pkt_r_instr_metadata__itag__2_, dispatch_pkt_r_instr_metadata__itag__1_, dispatch_pkt_r_instr_metadata__itag__0_, calc_status_o[187:124], dispatch_pkt_r_instr_metadata__fe_exception_not_instr_, dispatch_pkt_r_instr_metadata__fe_exception_code__1_, dispatch_pkt_r_instr_metadata__fe_exception_code__0_, calc_status_o[226:191], dispatch_pkt_r_instr__31_, dispatch_pkt_r_instr__30_, dispatch_pkt_r_instr__29_, dispatch_pkt_r_instr__28_, dispatch_pkt_r_instr__27_, dispatch_pkt_r_instr__26_, dispatch_pkt_r_instr__25_, dispatch_pkt_r_instr__24_, dispatch_pkt_r_instr__23_, dispatch_pkt_r_instr__22_, dispatch_pkt_r_instr__21_, dispatch_pkt_r_instr__20_, dispatch_pkt_r_instr__19_, dispatch_pkt_r_instr__18_, dispatch_pkt_r_instr__17_, dispatch_pkt_r_instr__16_, dispatch_pkt_r_instr__15_, dispatch_pkt_r_instr__14_, dispatch_pkt_r_instr__13_, dispatch_pkt_r_instr__12_, dispatch_pkt_r_instr__11_, dispatch_pkt_r_instr__10_, dispatch_pkt_r_instr__9_, dispatch_pkt_r_instr__8_, dispatch_pkt_r_instr__7_, dispatch_pkt_r_instr__6_, dispatch_pkt_r_instr__5_, dispatch_pkt_r_instr__4_, dispatch_pkt_r_instr__3_, dispatch_pkt_r_instr__2_, dispatch_pkt_r_instr__1_, dispatch_pkt_r_instr__0_, calc_status_o[188:188], dispatch_pkt_r_decode__fe_nop_v_, dispatch_pkt_r_decode__be_nop_v_, dispatch_pkt_r_decode__me_nop_v_, dispatch_pkt_r_decode__pipe_comp_v_, calc_status_o[291:291], dispatch_pkt_r_decode__pipe_mul_v_, dispatch_pkt_r_decode__pipe_mem_v_, dispatch_pkt_r_decode__pipe_fp_v_, dispatch_pkt_r_decode__irf_w_v_, dispatch_pkt_r_decode__frf_w_v_, dispatch_pkt_r_decode__csr_instr_v_, dispatch_pkt_r_decode__mhartid_r_v_, dispatch_pkt_r_decode__mcycle_r_v_, dispatch_pkt_r_decode__mtime_r_v_, dispatch_pkt_r_decode__minstret_r_v_, dispatch_pkt_r_decode__mtvec_rw_v_, dispatch_pkt_r_decode__mtval_rw_v_, dispatch_pkt_r_decode__mepc_rw_v_, dispatch_pkt_r_decode__mscratch_rw_v_, dispatch_pkt_r_decode__dcache_w_v_, dispatch_pkt_r_decode__dcache_r_v_, dispatch_pkt_r_decode__fp_not_int_v_, dispatch_pkt_r_decode__ret_v_, dispatch_pkt_r_decode__amo_v_, dispatch_pkt_r_decode__jmp_v_, dispatch_pkt_r_decode__br_v_, dispatch_pkt_r_decode__opw_v_, dispatch_pkt_r_decode__fu_op__fu_op__3_, dispatch_pkt_r_decode__fu_op__fu_op__2_, dispatch_pkt_r_decode__fu_op__fu_op__1_, dispatch_pkt_r_decode__fu_op__fu_op__0_, dispatch_pkt_r_decode__rs1_addr__4_, dispatch_pkt_r_decode__rs1_addr__3_, dispatch_pkt_r_decode__rs1_addr__2_, dispatch_pkt_r_decode__rs1_addr__1_, dispatch_pkt_r_decode__rs1_addr__0_, dispatch_pkt_r_decode__rs2_addr__4_, dispatch_pkt_r_decode__rs2_addr__3_, dispatch_pkt_r_decode__rs2_addr__2_, dispatch_pkt_r_decode__rs2_addr__1_, dispatch_pkt_r_decode__rs2_addr__0_, dispatch_pkt_r_decode__rd_addr__4_, dispatch_pkt_r_decode__rd_addr__3_, dispatch_pkt_r_decode__rd_addr__2_, dispatch_pkt_r_decode__rd_addr__1_, dispatch_pkt_r_decode__rd_addr__0_, dispatch_pkt_r_decode__src1_sel_, dispatch_pkt_r_decode__src2_sel_, dispatch_pkt_r_decode__baddr_sel_, dispatch_pkt_r_decode__result_sel_, dispatch_pkt_r_rs1__63_, dispatch_pkt_r_rs1__62_, dispatch_pkt_r_rs1__61_, dispatch_pkt_r_rs1__60_, dispatch_pkt_r_rs1__59_, dispatch_pkt_r_rs1__58_, dispatch_pkt_r_rs1__57_, dispatch_pkt_r_rs1__56_, dispatch_pkt_r_rs1__55_, dispatch_pkt_r_rs1__54_, dispatch_pkt_r_rs1__53_, dispatch_pkt_r_rs1__52_, dispatch_pkt_r_rs1__51_, dispatch_pkt_r_rs1__50_, dispatch_pkt_r_rs1__49_, dispatch_pkt_r_rs1__48_, dispatch_pkt_r_rs1__47_, dispatch_pkt_r_rs1__46_, dispatch_pkt_r_rs1__45_, dispatch_pkt_r_rs1__44_, dispatch_pkt_r_rs1__43_, dispatch_pkt_r_rs1__42_, dispatch_pkt_r_rs1__41_, dispatch_pkt_r_rs1__40_, dispatch_pkt_r_rs1__39_, dispatch_pkt_r_rs1__38_, dispatch_pkt_r_rs1__37_, dispatch_pkt_r_rs1__36_, dispatch_pkt_r_rs1__35_, dispatch_pkt_r_rs1__34_, dispatch_pkt_r_rs1__33_, dispatch_pkt_r_rs1__32_, dispatch_pkt_r_rs1__31_, dispatch_pkt_r_rs1__30_, dispatch_pkt_r_rs1__29_, dispatch_pkt_r_rs1__28_, dispatch_pkt_r_rs1__27_, dispatch_pkt_r_rs1__26_, dispatch_pkt_r_rs1__25_, dispatch_pkt_r_rs1__24_, dispatch_pkt_r_rs1__23_, dispatch_pkt_r_rs1__22_, dispatch_pkt_r_rs1__21_, dispatch_pkt_r_rs1__20_, dispatch_pkt_r_rs1__19_, dispatch_pkt_r_rs1__18_, dispatch_pkt_r_rs1__17_, dispatch_pkt_r_rs1__16_, dispatch_pkt_r_rs1__15_, dispatch_pkt_r_rs1__14_, dispatch_pkt_r_rs1__13_, dispatch_pkt_r_rs1__12_, dispatch_pkt_r_rs1__11_, dispatch_pkt_r_rs1__10_, dispatch_pkt_r_rs1__9_, dispatch_pkt_r_rs1__8_, dispatch_pkt_r_rs1__7_, dispatch_pkt_r_rs1__6_, dispatch_pkt_r_rs1__5_, dispatch_pkt_r_rs1__4_, dispatch_pkt_r_rs1__3_, dispatch_pkt_r_rs1__2_, dispatch_pkt_r_rs1__1_, dispatch_pkt_r_rs1__0_, dispatch_pkt_r_rs2__63_, dispatch_pkt_r_rs2__62_, dispatch_pkt_r_rs2__61_, dispatch_pkt_r_rs2__60_, dispatch_pkt_r_rs2__59_, dispatch_pkt_r_rs2__58_, dispatch_pkt_r_rs2__57_, dispatch_pkt_r_rs2__56_, dispatch_pkt_r_rs2__55_, dispatch_pkt_r_rs2__54_, dispatch_pkt_r_rs2__53_, dispatch_pkt_r_rs2__52_, dispatch_pkt_r_rs2__51_, dispatch_pkt_r_rs2__50_, dispatch_pkt_r_rs2__49_, dispatch_pkt_r_rs2__48_, dispatch_pkt_r_rs2__47_, dispatch_pkt_r_rs2__46_, dispatch_pkt_r_rs2__45_, dispatch_pkt_r_rs2__44_, dispatch_pkt_r_rs2__43_, dispatch_pkt_r_rs2__42_, dispatch_pkt_r_rs2__41_, dispatch_pkt_r_rs2__40_, dispatch_pkt_r_rs2__39_, dispatch_pkt_r_rs2__38_, dispatch_pkt_r_rs2__37_, dispatch_pkt_r_rs2__36_, dispatch_pkt_r_rs2__35_, dispatch_pkt_r_rs2__34_, dispatch_pkt_r_rs2__33_, dispatch_pkt_r_rs2__32_, dispatch_pkt_r_rs2__31_, dispatch_pkt_r_rs2__30_, dispatch_pkt_r_rs2__29_, dispatch_pkt_r_rs2__28_, dispatch_pkt_r_rs2__27_, dispatch_pkt_r_rs2__26_, dispatch_pkt_r_rs2__25_, dispatch_pkt_r_rs2__24_, dispatch_pkt_r_rs2__23_, dispatch_pkt_r_rs2__22_, dispatch_pkt_r_rs2__21_, dispatch_pkt_r_rs2__20_, dispatch_pkt_r_rs2__19_, dispatch_pkt_r_rs2__18_, dispatch_pkt_r_rs2__17_, dispatch_pkt_r_rs2__16_, dispatch_pkt_r_rs2__15_, dispatch_pkt_r_rs2__14_, dispatch_pkt_r_rs2__13_, dispatch_pkt_r_rs2__12_, dispatch_pkt_r_rs2__11_, dispatch_pkt_r_rs2__10_, dispatch_pkt_r_rs2__9_, dispatch_pkt_r_rs2__8_, dispatch_pkt_r_rs2__7_, dispatch_pkt_r_rs2__6_, dispatch_pkt_r_rs2__5_, dispatch_pkt_r_rs2__4_, dispatch_pkt_r_rs2__3_, dispatch_pkt_r_rs2__2_, dispatch_pkt_r_rs2__1_, dispatch_pkt_r_rs2__0_, dispatch_pkt_r_imm__63_, dispatch_pkt_r_imm__62_, dispatch_pkt_r_imm__61_, dispatch_pkt_r_imm__60_, dispatch_pkt_r_imm__59_, dispatch_pkt_r_imm__58_, dispatch_pkt_r_imm__57_, dispatch_pkt_r_imm__56_, dispatch_pkt_r_imm__55_, dispatch_pkt_r_imm__54_, dispatch_pkt_r_imm__53_, dispatch_pkt_r_imm__52_, dispatch_pkt_r_imm__51_, dispatch_pkt_r_imm__50_, dispatch_pkt_r_imm__49_, dispatch_pkt_r_imm__48_, dispatch_pkt_r_imm__47_, dispatch_pkt_r_imm__46_, dispatch_pkt_r_imm__45_, dispatch_pkt_r_imm__44_, dispatch_pkt_r_imm__43_, dispatch_pkt_r_imm__42_, dispatch_pkt_r_imm__41_, dispatch_pkt_r_imm__40_, dispatch_pkt_r_imm__39_, dispatch_pkt_r_imm__38_, dispatch_pkt_r_imm__37_, dispatch_pkt_r_imm__36_, dispatch_pkt_r_imm__35_, dispatch_pkt_r_imm__34_, dispatch_pkt_r_imm__33_, dispatch_pkt_r_imm__32_, dispatch_pkt_r_imm__31_, dispatch_pkt_r_imm__30_, dispatch_pkt_r_imm__29_, dispatch_pkt_r_imm__28_, dispatch_pkt_r_imm__27_, dispatch_pkt_r_imm__26_, dispatch_pkt_r_imm__25_, dispatch_pkt_r_imm__24_, dispatch_pkt_r_imm__23_, dispatch_pkt_r_imm__22_, dispatch_pkt_r_imm__21_, dispatch_pkt_r_imm__20_, dispatch_pkt_r_imm__19_, dispatch_pkt_r_imm__18_, dispatch_pkt_r_imm__17_, dispatch_pkt_r_imm__16_, dispatch_pkt_r_imm__15_, dispatch_pkt_r_imm__14_, dispatch_pkt_r_imm__13_, dispatch_pkt_r_imm__12_, dispatch_pkt_r_imm__11_, dispatch_pkt_r_imm__10_, dispatch_pkt_r_imm__9_, dispatch_pkt_r_imm__8_, dispatch_pkt_r_imm__7_, dispatch_pkt_r_imm__6_, dispatch_pkt_r_imm__5_, dispatch_pkt_r_imm__4_, dispatch_pkt_r_imm__3_, dispatch_pkt_r_imm__2_, dispatch_pkt_r_imm__1_, dispatch_pkt_r_imm__0_ })
  );


  bsg_mux_segmented_segments_p5_segment_width_p64
  comp_stage_mux
  (
    .data0_i({ comp_stage_r[255:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .data1_i({ pipe_fp_data_lo, pipe_mem_data_lo, pipe_mul_data_lo, pipe_int_data_lo, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_i({ calc_stage_r_3__pipe_fp_v_, calc_stage_r_2__pipe_mem_v_, calc_stage_r_1__pipe_mul_v_, calc_stage_r_0__pipe_int_v_, 1'b1 }),
    .data_o(comp_stage_n)
  );


  bsg_dff_width_p320
  comp_stage_reg
  (
    .clk_i(clk_i),
    .data_i(comp_stage_n),
    .data_o(comp_stage_r)
  );


  bsg_dff_width_p45
  exc_stage_reg
  (
    .clk_i(clk_i),
    .data_i({ exc_stage_n_4__poison_v_, exc_stage_r_3__roll_v_, exc_stage_r_3__illegal_instr_v_, exc_stage_r_3__ret_instr_v_, exc_stage_r_3__csr_instr_v_, exc_stage_r_3__tlb_miss_v_, exc_stage_r_3__load_fault_v_, exc_stage_r_3__store_fault_v_, exc_stage_r_3__cache_miss_v_, exc_stage_n_3__poison_v_, exc_stage_n_3__roll_v_, exc_stage_r_2__illegal_instr_v_, exc_stage_r_2__ret_instr_v_, exc_stage_r_2__csr_instr_v_, exc_stage_r_2__tlb_miss_v_, exc_stage_r_2__load_fault_v_, exc_stage_r_2__store_fault_v_, exc_stage_n_3__cache_miss_v_, exc_stage_n_2__poison_v_, exc_stage_n_2__roll_v_, exc_stage_r_1__illegal_instr_v_, exc_stage_r_1__ret_instr_v_, exc_stage_r_1__csr_instr_v_, exc_stage_r_1__tlb_miss_v_, exc_stage_r_1__load_fault_v_, exc_stage_r_1__store_fault_v_, exc_stage_r_1__cache_miss_v_, exc_stage_n_1__poison_v_, exc_stage_n_1__roll_v_, exc_stage_r_0__illegal_instr_v_, exc_stage_r_0__ret_instr_v_, exc_stage_r_0__csr_instr_v_, exc_stage_r_0__tlb_miss_v_, exc_stage_r_0__load_fault_v_, exc_stage_r_0__store_fault_v_, exc_stage_r_0__cache_miss_v_, chk_poison_isd_i, chk_roll_i, exc_stage_n_0__illegal_instr_v_, exc_stage_n_0__ret_instr_v_, exc_stage_n_0__csr_instr_v_, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .data_o({ exc_stage_r_4__poison_v_, exc_stage_r_4__roll_v_, exc_stage_r_4__illegal_instr_v_, exc_stage_r_4__ret_instr_v_, exc_stage_r_4__csr_instr_v_, exc_stage_r_4__tlb_miss_v_, exc_stage_r_4__load_fault_v_, exc_stage_r_4__store_fault_v_, exc_stage_r_4__cache_miss_v_, exc_stage_n_4__poison_v_, exc_stage_r_3__roll_v_, exc_stage_r_3__illegal_instr_v_, exc_stage_r_3__ret_instr_v_, exc_stage_r_3__csr_instr_v_, exc_stage_r_3__tlb_miss_v_, exc_stage_r_3__load_fault_v_, exc_stage_r_3__store_fault_v_, exc_stage_r_3__cache_miss_v_, exc_stage_r_2__poison_v_, exc_stage_r_2__roll_v_, exc_stage_r_2__illegal_instr_v_, exc_stage_r_2__ret_instr_v_, exc_stage_r_2__csr_instr_v_, exc_stage_r_2__tlb_miss_v_, exc_stage_r_2__load_fault_v_, exc_stage_r_2__store_fault_v_, exc_stage_r_2__cache_miss_v_, exc_stage_r_1__poison_v_, exc_stage_r_1__roll_v_, exc_stage_r_1__illegal_instr_v_, exc_stage_r_1__ret_instr_v_, exc_stage_r_1__csr_instr_v_, exc_stage_r_1__tlb_miss_v_, exc_stage_r_1__load_fault_v_, exc_stage_r_1__store_fault_v_, exc_stage_r_1__cache_miss_v_, exc_stage_r_0__poison_v_, exc_stage_r_0__roll_v_, exc_stage_r_0__illegal_instr_v_, exc_stage_r_0__ret_instr_v_, exc_stage_r_0__csr_instr_v_, exc_stage_r_0__tlb_miss_v_, exc_stage_r_0__load_fault_v_, exc_stage_r_0__store_fault_v_, exc_stage_r_0__cache_miss_v_ })
  );


  bsg_counter_clear_up_init_val_p0_ptr_width_lp64
  cycle_counter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(1'b0),
    .up_i(1'b1),
    .count_o(cycle_cnt_lo)
  );


  bsg_counter_clear_up_init_val_p0_ptr_width_lp64
  time_counter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(1'b0),
    .up_i(1'b1),
    .count_o(time_cnt_lo)
  );


  bsg_counter_clear_up_init_val_p0_ptr_width_lp64
  instret_counter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(1'b0),
    .up_i(n_63_net_),
    .count_o(instret_cnt_lo)
  );


  bsg_dff_en_width_p64
  mtval_csr_reg
  (
    .clk_i(clk_i),
    .data_i(mtval_mux_lo),
    .en_i(n_64_net_),
    .data_o(mtval_li)
  );


  bsg_mux_width_p64_els_p2
  mtval_mux
  (
    .data_i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, calc_stage_r_2__instr__31_, calc_stage_r_2__instr__30_, calc_stage_r_2__instr__29_, calc_stage_r_2__instr__28_, calc_stage_r_2__instr__27_, calc_stage_r_2__instr__26_, calc_stage_r_2__instr__25_, calc_stage_r_2__instr__24_, calc_stage_r_2__instr__23_, calc_stage_r_2__instr__22_, calc_stage_r_2__instr__21_, calc_stage_r_2__instr__20_, calc_stage_r_2__instr__19_, calc_stage_r_2__instr__18_, calc_stage_r_2__instr__17_, calc_stage_r_2__instr__16_, calc_stage_r_2__instr__15_, calc_stage_r_2__instr__14_, calc_stage_r_2__instr__13_, calc_stage_r_2__instr__12_, calc_stage_r_2__instr__11_, calc_stage_r_2__instr__10_, calc_stage_r_2__instr__9_, calc_stage_r_2__instr__8_, calc_stage_r_2__instr__7_, calc_stage_r_2__instr__6_, calc_stage_r_2__instr__5_, calc_stage_r_2__instr__4_, calc_stage_r_2__instr__3_, calc_stage_r_2__instr__2_, calc_stage_r_2__instr__1_, calc_stage_r_2__instr__0_, mtval_lo }),
    .sel_i(calc_status_o[2]),
    .data_o(mtval_mux_lo)
  );


  bsg_dff_en_width_p64
  mscratch_csr_reg
  (
    .clk_i(clk_i),
    .data_i(mscratch_lo),
    .en_i(mscratch_w_v_lo),
    .data_o(mscratch_li)
  );

  assign dispatch_pkt[0] = issue_pkt_r_imm__0_;
  assign dispatch_pkt[1] = issue_pkt_r_imm__1_;
  assign dispatch_pkt[2] = issue_pkt_r_imm__2_;
  assign dispatch_pkt[3] = issue_pkt_r_imm__3_;
  assign dispatch_pkt[4] = issue_pkt_r_imm__4_;
  assign dispatch_pkt[5] = issue_pkt_r_imm__5_;
  assign dispatch_pkt[6] = issue_pkt_r_imm__6_;
  assign dispatch_pkt[7] = issue_pkt_r_imm__7_;
  assign dispatch_pkt[8] = issue_pkt_r_imm__8_;
  assign dispatch_pkt[9] = issue_pkt_r_imm__9_;
  assign dispatch_pkt[10] = issue_pkt_r_imm__10_;
  assign dispatch_pkt[11] = issue_pkt_r_imm__11_;
  assign dispatch_pkt[12] = issue_pkt_r_imm__12_;
  assign dispatch_pkt[13] = issue_pkt_r_imm__13_;
  assign dispatch_pkt[14] = issue_pkt_r_imm__14_;
  assign dispatch_pkt[15] = issue_pkt_r_imm__15_;
  assign dispatch_pkt[16] = issue_pkt_r_imm__16_;
  assign dispatch_pkt[17] = issue_pkt_r_imm__17_;
  assign dispatch_pkt[18] = issue_pkt_r_imm__18_;
  assign dispatch_pkt[19] = issue_pkt_r_imm__19_;
  assign dispatch_pkt[20] = issue_pkt_r_imm__20_;
  assign dispatch_pkt[21] = issue_pkt_r_imm__21_;
  assign dispatch_pkt[22] = issue_pkt_r_imm__22_;
  assign dispatch_pkt[23] = issue_pkt_r_imm__23_;
  assign dispatch_pkt[24] = issue_pkt_r_imm__24_;
  assign dispatch_pkt[25] = issue_pkt_r_imm__25_;
  assign dispatch_pkt[26] = issue_pkt_r_imm__26_;
  assign dispatch_pkt[27] = issue_pkt_r_imm__27_;
  assign dispatch_pkt[28] = issue_pkt_r_imm__28_;
  assign dispatch_pkt[29] = issue_pkt_r_imm__29_;
  assign dispatch_pkt[30] = issue_pkt_r_imm__30_;
  assign dispatch_pkt[31] = issue_pkt_r_imm__31_;
  assign dispatch_pkt[32] = issue_pkt_r_imm__32_;
  assign dispatch_pkt[33] = issue_pkt_r_imm__33_;
  assign dispatch_pkt[34] = issue_pkt_r_imm__34_;
  assign dispatch_pkt[35] = issue_pkt_r_imm__35_;
  assign dispatch_pkt[36] = issue_pkt_r_imm__36_;
  assign dispatch_pkt[37] = issue_pkt_r_imm__37_;
  assign dispatch_pkt[38] = issue_pkt_r_imm__38_;
  assign dispatch_pkt[39] = issue_pkt_r_imm__39_;
  assign dispatch_pkt[40] = issue_pkt_r_imm__40_;
  assign dispatch_pkt[41] = issue_pkt_r_imm__41_;
  assign dispatch_pkt[42] = issue_pkt_r_imm__42_;
  assign dispatch_pkt[43] = issue_pkt_r_imm__43_;
  assign dispatch_pkt[44] = issue_pkt_r_imm__44_;
  assign dispatch_pkt[45] = issue_pkt_r_imm__45_;
  assign dispatch_pkt[46] = issue_pkt_r_imm__46_;
  assign dispatch_pkt[47] = issue_pkt_r_imm__47_;
  assign dispatch_pkt[48] = issue_pkt_r_imm__48_;
  assign dispatch_pkt[49] = issue_pkt_r_imm__49_;
  assign dispatch_pkt[50] = issue_pkt_r_imm__50_;
  assign dispatch_pkt[51] = issue_pkt_r_imm__51_;
  assign dispatch_pkt[52] = issue_pkt_r_imm__52_;
  assign dispatch_pkt[53] = issue_pkt_r_imm__53_;
  assign dispatch_pkt[54] = issue_pkt_r_imm__54_;
  assign dispatch_pkt[55] = issue_pkt_r_imm__55_;
  assign dispatch_pkt[56] = issue_pkt_r_imm__56_;
  assign dispatch_pkt[57] = issue_pkt_r_imm__57_;
  assign dispatch_pkt[58] = issue_pkt_r_imm__58_;
  assign dispatch_pkt[59] = issue_pkt_r_imm__59_;
  assign dispatch_pkt[60] = issue_pkt_r_imm__60_;
  assign dispatch_pkt[61] = issue_pkt_r_imm__61_;
  assign dispatch_pkt[62] = issue_pkt_r_imm__62_;
  assign dispatch_pkt[63] = issue_pkt_r_imm__63_;
  assign dispatch_pkt[64] = bypass_rs2[0];
  assign dispatch_pkt[65] = bypass_rs2[1];
  assign dispatch_pkt[66] = bypass_rs2[2];
  assign dispatch_pkt[67] = bypass_rs2[3];
  assign dispatch_pkt[68] = bypass_rs2[4];
  assign dispatch_pkt[69] = bypass_rs2[5];
  assign dispatch_pkt[70] = bypass_rs2[6];
  assign dispatch_pkt[71] = bypass_rs2[7];
  assign dispatch_pkt[72] = bypass_rs2[8];
  assign dispatch_pkt[73] = bypass_rs2[9];
  assign dispatch_pkt[74] = bypass_rs2[10];
  assign dispatch_pkt[75] = bypass_rs2[11];
  assign dispatch_pkt[76] = bypass_rs2[12];
  assign dispatch_pkt[77] = bypass_rs2[13];
  assign dispatch_pkt[78] = bypass_rs2[14];
  assign dispatch_pkt[79] = bypass_rs2[15];
  assign dispatch_pkt[80] = bypass_rs2[16];
  assign dispatch_pkt[81] = bypass_rs2[17];
  assign dispatch_pkt[82] = bypass_rs2[18];
  assign dispatch_pkt[83] = bypass_rs2[19];
  assign dispatch_pkt[84] = bypass_rs2[20];
  assign dispatch_pkt[85] = bypass_rs2[21];
  assign dispatch_pkt[86] = bypass_rs2[22];
  assign dispatch_pkt[87] = bypass_rs2[23];
  assign dispatch_pkt[88] = bypass_rs2[24];
  assign dispatch_pkt[89] = bypass_rs2[25];
  assign dispatch_pkt[90] = bypass_rs2[26];
  assign dispatch_pkt[91] = bypass_rs2[27];
  assign dispatch_pkt[92] = bypass_rs2[28];
  assign dispatch_pkt[93] = bypass_rs2[29];
  assign dispatch_pkt[94] = bypass_rs2[30];
  assign dispatch_pkt[95] = bypass_rs2[31];
  assign dispatch_pkt[96] = bypass_rs2[32];
  assign dispatch_pkt[97] = bypass_rs2[33];
  assign dispatch_pkt[98] = bypass_rs2[34];
  assign dispatch_pkt[99] = bypass_rs2[35];
  assign dispatch_pkt[100] = bypass_rs2[36];
  assign dispatch_pkt[101] = bypass_rs2[37];
  assign dispatch_pkt[102] = bypass_rs2[38];
  assign dispatch_pkt[103] = bypass_rs2[39];
  assign dispatch_pkt[104] = bypass_rs2[40];
  assign dispatch_pkt[105] = bypass_rs2[41];
  assign dispatch_pkt[106] = bypass_rs2[42];
  assign dispatch_pkt[107] = bypass_rs2[43];
  assign dispatch_pkt[108] = bypass_rs2[44];
  assign dispatch_pkt[109] = bypass_rs2[45];
  assign dispatch_pkt[110] = bypass_rs2[46];
  assign dispatch_pkt[111] = bypass_rs2[47];
  assign dispatch_pkt[112] = bypass_rs2[48];
  assign dispatch_pkt[113] = bypass_rs2[49];
  assign dispatch_pkt[114] = bypass_rs2[50];
  assign dispatch_pkt[115] = bypass_rs2[51];
  assign dispatch_pkt[116] = bypass_rs2[52];
  assign dispatch_pkt[117] = bypass_rs2[53];
  assign dispatch_pkt[118] = bypass_rs2[54];
  assign dispatch_pkt[119] = bypass_rs2[55];
  assign dispatch_pkt[120] = bypass_rs2[56];
  assign dispatch_pkt[121] = bypass_rs2[57];
  assign dispatch_pkt[122] = bypass_rs2[58];
  assign dispatch_pkt[123] = bypass_rs2[59];
  assign dispatch_pkt[124] = bypass_rs2[60];
  assign dispatch_pkt[125] = bypass_rs2[61];
  assign dispatch_pkt[126] = bypass_rs2[62];
  assign dispatch_pkt[127] = bypass_rs2[63];
  assign dispatch_pkt[128] = bypass_rs1[0];
  assign dispatch_pkt[129] = bypass_rs1[1];
  assign dispatch_pkt[130] = bypass_rs1[2];
  assign dispatch_pkt[131] = bypass_rs1[3];
  assign dispatch_pkt[132] = bypass_rs1[4];
  assign dispatch_pkt[133] = bypass_rs1[5];
  assign dispatch_pkt[134] = bypass_rs1[6];
  assign dispatch_pkt[135] = bypass_rs1[7];
  assign dispatch_pkt[136] = bypass_rs1[8];
  assign dispatch_pkt[137] = bypass_rs1[9];
  assign dispatch_pkt[138] = bypass_rs1[10];
  assign dispatch_pkt[139] = bypass_rs1[11];
  assign dispatch_pkt[140] = bypass_rs1[12];
  assign dispatch_pkt[141] = bypass_rs1[13];
  assign dispatch_pkt[142] = bypass_rs1[14];
  assign dispatch_pkt[143] = bypass_rs1[15];
  assign dispatch_pkt[144] = bypass_rs1[16];
  assign dispatch_pkt[145] = bypass_rs1[17];
  assign dispatch_pkt[146] = bypass_rs1[18];
  assign dispatch_pkt[147] = bypass_rs1[19];
  assign dispatch_pkt[148] = bypass_rs1[20];
  assign dispatch_pkt[149] = bypass_rs1[21];
  assign dispatch_pkt[150] = bypass_rs1[22];
  assign dispatch_pkt[151] = bypass_rs1[23];
  assign dispatch_pkt[152] = bypass_rs1[24];
  assign dispatch_pkt[153] = bypass_rs1[25];
  assign dispatch_pkt[154] = bypass_rs1[26];
  assign dispatch_pkt[155] = bypass_rs1[27];
  assign dispatch_pkt[156] = bypass_rs1[28];
  assign dispatch_pkt[157] = bypass_rs1[29];
  assign dispatch_pkt[158] = bypass_rs1[30];
  assign dispatch_pkt[159] = bypass_rs1[31];
  assign dispatch_pkt[160] = bypass_rs1[32];
  assign dispatch_pkt[161] = bypass_rs1[33];
  assign dispatch_pkt[162] = bypass_rs1[34];
  assign dispatch_pkt[163] = bypass_rs1[35];
  assign dispatch_pkt[164] = bypass_rs1[36];
  assign dispatch_pkt[165] = bypass_rs1[37];
  assign dispatch_pkt[166] = bypass_rs1[38];
  assign dispatch_pkt[167] = bypass_rs1[39];
  assign dispatch_pkt[168] = bypass_rs1[40];
  assign dispatch_pkt[169] = bypass_rs1[41];
  assign dispatch_pkt[170] = bypass_rs1[42];
  assign dispatch_pkt[171] = bypass_rs1[43];
  assign dispatch_pkt[172] = bypass_rs1[44];
  assign dispatch_pkt[173] = bypass_rs1[45];
  assign dispatch_pkt[174] = bypass_rs1[46];
  assign dispatch_pkt[175] = bypass_rs1[47];
  assign dispatch_pkt[176] = bypass_rs1[48];
  assign dispatch_pkt[177] = bypass_rs1[49];
  assign dispatch_pkt[178] = bypass_rs1[50];
  assign dispatch_pkt[179] = bypass_rs1[51];
  assign dispatch_pkt[180] = bypass_rs1[52];
  assign dispatch_pkt[181] = bypass_rs1[53];
  assign dispatch_pkt[182] = bypass_rs1[54];
  assign dispatch_pkt[183] = bypass_rs1[55];
  assign dispatch_pkt[184] = bypass_rs1[56];
  assign dispatch_pkt[185] = bypass_rs1[57];
  assign dispatch_pkt[186] = bypass_rs1[58];
  assign dispatch_pkt[187] = bypass_rs1[59];
  assign dispatch_pkt[188] = bypass_rs1[60];
  assign dispatch_pkt[189] = bypass_rs1[61];
  assign dispatch_pkt[190] = bypass_rs1[62];
  assign dispatch_pkt[191] = bypass_rs1[63];
  assign dispatch_pkt[243] = issue_pkt_r_instr__0_;
  assign dispatch_pkt[244] = issue_pkt_r_instr__1_;
  assign dispatch_pkt[245] = issue_pkt_r_instr__2_;
  assign dispatch_pkt[246] = issue_pkt_r_instr__3_;
  assign dispatch_pkt[247] = issue_pkt_r_instr__4_;
  assign dispatch_pkt[248] = issue_pkt_r_instr__5_;
  assign dispatch_pkt[249] = issue_pkt_r_instr__6_;
  assign dispatch_pkt[250] = issue_pkt_r_instr__7_;
  assign dispatch_pkt[251] = issue_pkt_r_instr__8_;
  assign dispatch_pkt[252] = issue_pkt_r_instr__9_;
  assign dispatch_pkt[253] = issue_pkt_r_instr__10_;
  assign dispatch_pkt[254] = issue_pkt_r_instr__11_;
  assign dispatch_pkt[255] = issue_pkt_r_instr__12_;
  assign dispatch_pkt[256] = issue_pkt_r_instr__13_;
  assign dispatch_pkt[257] = issue_pkt_r_instr__14_;
  assign dispatch_pkt[258] = issue_pkt_r_instr__15_;
  assign dispatch_pkt[259] = issue_pkt_r_instr__16_;
  assign dispatch_pkt[260] = issue_pkt_r_instr__17_;
  assign dispatch_pkt[261] = issue_pkt_r_instr__18_;
  assign dispatch_pkt[262] = issue_pkt_r_instr__19_;
  assign dispatch_pkt[263] = issue_pkt_r_instr__20_;
  assign dispatch_pkt[264] = issue_pkt_r_instr__21_;
  assign dispatch_pkt[265] = issue_pkt_r_instr__22_;
  assign dispatch_pkt[266] = issue_pkt_r_instr__23_;
  assign dispatch_pkt[267] = issue_pkt_r_instr__24_;
  assign dispatch_pkt[268] = issue_pkt_r_instr__25_;
  assign dispatch_pkt[269] = issue_pkt_r_instr__26_;
  assign dispatch_pkt[270] = issue_pkt_r_instr__27_;
  assign dispatch_pkt[271] = issue_pkt_r_instr__28_;
  assign dispatch_pkt[272] = issue_pkt_r_instr__29_;
  assign dispatch_pkt[273] = issue_pkt_r_instr__30_;
  assign dispatch_pkt[274] = issue_pkt_r_instr__31_;
  assign dispatch_pkt[275] = issue_pkt_r_branch_metadata_fwd__0_;
  assign dispatch_pkt[276] = issue_pkt_r_branch_metadata_fwd__1_;
  assign dispatch_pkt[277] = issue_pkt_r_branch_metadata_fwd__2_;
  assign dispatch_pkt[278] = issue_pkt_r_branch_metadata_fwd__3_;
  assign dispatch_pkt[279] = issue_pkt_r_branch_metadata_fwd__4_;
  assign dispatch_pkt[280] = issue_pkt_r_branch_metadata_fwd__5_;
  assign dispatch_pkt[281] = issue_pkt_r_branch_metadata_fwd__6_;
  assign dispatch_pkt[282] = issue_pkt_r_branch_metadata_fwd__7_;
  assign dispatch_pkt[283] = issue_pkt_r_branch_metadata_fwd__8_;
  assign dispatch_pkt[284] = issue_pkt_r_branch_metadata_fwd__9_;
  assign dispatch_pkt[285] = issue_pkt_r_branch_metadata_fwd__10_;
  assign dispatch_pkt[286] = issue_pkt_r_branch_metadata_fwd__11_;
  assign dispatch_pkt[287] = issue_pkt_r_branch_metadata_fwd__12_;
  assign dispatch_pkt[288] = issue_pkt_r_branch_metadata_fwd__13_;
  assign dispatch_pkt[289] = issue_pkt_r_branch_metadata_fwd__14_;
  assign dispatch_pkt[290] = issue_pkt_r_branch_metadata_fwd__15_;
  assign dispatch_pkt[291] = issue_pkt_r_branch_metadata_fwd__16_;
  assign dispatch_pkt[292] = issue_pkt_r_branch_metadata_fwd__17_;
  assign dispatch_pkt[293] = issue_pkt_r_branch_metadata_fwd__18_;
  assign dispatch_pkt[294] = issue_pkt_r_branch_metadata_fwd__19_;
  assign dispatch_pkt[295] = issue_pkt_r_branch_metadata_fwd__20_;
  assign dispatch_pkt[296] = issue_pkt_r_branch_metadata_fwd__21_;
  assign dispatch_pkt[297] = issue_pkt_r_branch_metadata_fwd__22_;
  assign dispatch_pkt[298] = issue_pkt_r_branch_metadata_fwd__23_;
  assign dispatch_pkt[299] = issue_pkt_r_branch_metadata_fwd__24_;
  assign dispatch_pkt[300] = issue_pkt_r_branch_metadata_fwd__25_;
  assign dispatch_pkt[301] = issue_pkt_r_branch_metadata_fwd__26_;
  assign dispatch_pkt[302] = issue_pkt_r_branch_metadata_fwd__27_;
  assign dispatch_pkt[303] = issue_pkt_r_branch_metadata_fwd__28_;
  assign dispatch_pkt[304] = issue_pkt_r_branch_metadata_fwd__29_;
  assign dispatch_pkt[305] = issue_pkt_r_branch_metadata_fwd__30_;
  assign dispatch_pkt[306] = issue_pkt_r_branch_metadata_fwd__31_;
  assign dispatch_pkt[307] = issue_pkt_r_branch_metadata_fwd__32_;
  assign dispatch_pkt[308] = issue_pkt_r_branch_metadata_fwd__33_;
  assign dispatch_pkt[309] = issue_pkt_r_branch_metadata_fwd__34_;
  assign dispatch_pkt[310] = issue_pkt_r_branch_metadata_fwd__35_;
  assign dispatch_pkt[311] = issue_pkt_r_instr_metadata__fe_exception_code__0_;
  assign dispatch_pkt[312] = issue_pkt_r_instr_metadata__fe_exception_code__1_;
  assign dispatch_pkt[313] = issue_pkt_r_instr_metadata__fe_exception_not_instr_;
  assign dispatch_pkt[314] = issue_pkt_r_instr_metadata__pc__0_;
  assign dispatch_pkt[315] = issue_pkt_r_instr_metadata__pc__1_;
  assign dispatch_pkt[316] = issue_pkt_r_instr_metadata__pc__2_;
  assign dispatch_pkt[317] = issue_pkt_r_instr_metadata__pc__3_;
  assign dispatch_pkt[318] = issue_pkt_r_instr_metadata__pc__4_;
  assign dispatch_pkt[319] = issue_pkt_r_instr_metadata__pc__5_;
  assign dispatch_pkt[320] = issue_pkt_r_instr_metadata__pc__6_;
  assign dispatch_pkt[321] = issue_pkt_r_instr_metadata__pc__7_;
  assign dispatch_pkt[322] = issue_pkt_r_instr_metadata__pc__8_;
  assign dispatch_pkt[323] = issue_pkt_r_instr_metadata__pc__9_;
  assign dispatch_pkt[324] = issue_pkt_r_instr_metadata__pc__10_;
  assign dispatch_pkt[325] = issue_pkt_r_instr_metadata__pc__11_;
  assign dispatch_pkt[326] = issue_pkt_r_instr_metadata__pc__12_;
  assign dispatch_pkt[327] = issue_pkt_r_instr_metadata__pc__13_;
  assign dispatch_pkt[328] = issue_pkt_r_instr_metadata__pc__14_;
  assign dispatch_pkt[329] = issue_pkt_r_instr_metadata__pc__15_;
  assign dispatch_pkt[330] = issue_pkt_r_instr_metadata__pc__16_;
  assign dispatch_pkt[331] = issue_pkt_r_instr_metadata__pc__17_;
  assign dispatch_pkt[332] = issue_pkt_r_instr_metadata__pc__18_;
  assign dispatch_pkt[333] = issue_pkt_r_instr_metadata__pc__19_;
  assign dispatch_pkt[334] = issue_pkt_r_instr_metadata__pc__20_;
  assign dispatch_pkt[335] = issue_pkt_r_instr_metadata__pc__21_;
  assign dispatch_pkt[336] = issue_pkt_r_instr_metadata__pc__22_;
  assign dispatch_pkt[337] = issue_pkt_r_instr_metadata__pc__23_;
  assign dispatch_pkt[338] = issue_pkt_r_instr_metadata__pc__24_;
  assign dispatch_pkt[339] = issue_pkt_r_instr_metadata__pc__25_;
  assign dispatch_pkt[340] = issue_pkt_r_instr_metadata__pc__26_;
  assign dispatch_pkt[341] = issue_pkt_r_instr_metadata__pc__27_;
  assign dispatch_pkt[342] = issue_pkt_r_instr_metadata__pc__28_;
  assign dispatch_pkt[343] = issue_pkt_r_instr_metadata__pc__29_;
  assign dispatch_pkt[344] = issue_pkt_r_instr_metadata__pc__30_;
  assign dispatch_pkt[345] = issue_pkt_r_instr_metadata__pc__31_;
  assign dispatch_pkt[346] = issue_pkt_r_instr_metadata__pc__32_;
  assign dispatch_pkt[347] = issue_pkt_r_instr_metadata__pc__33_;
  assign dispatch_pkt[348] = issue_pkt_r_instr_metadata__pc__34_;
  assign dispatch_pkt[349] = issue_pkt_r_instr_metadata__pc__35_;
  assign dispatch_pkt[350] = issue_pkt_r_instr_metadata__pc__36_;
  assign dispatch_pkt[351] = issue_pkt_r_instr_metadata__pc__37_;
  assign dispatch_pkt[352] = issue_pkt_r_instr_metadata__pc__38_;
  assign dispatch_pkt[353] = issue_pkt_r_instr_metadata__pc__39_;
  assign dispatch_pkt[354] = issue_pkt_r_instr_metadata__pc__40_;
  assign dispatch_pkt[355] = issue_pkt_r_instr_metadata__pc__41_;
  assign dispatch_pkt[356] = issue_pkt_r_instr_metadata__pc__42_;
  assign dispatch_pkt[357] = issue_pkt_r_instr_metadata__pc__43_;
  assign dispatch_pkt[358] = issue_pkt_r_instr_metadata__pc__44_;
  assign dispatch_pkt[359] = issue_pkt_r_instr_metadata__pc__45_;
  assign dispatch_pkt[360] = issue_pkt_r_instr_metadata__pc__46_;
  assign dispatch_pkt[361] = issue_pkt_r_instr_metadata__pc__47_;
  assign dispatch_pkt[362] = issue_pkt_r_instr_metadata__pc__48_;
  assign dispatch_pkt[363] = issue_pkt_r_instr_metadata__pc__49_;
  assign dispatch_pkt[364] = issue_pkt_r_instr_metadata__pc__50_;
  assign dispatch_pkt[365] = issue_pkt_r_instr_metadata__pc__51_;
  assign dispatch_pkt[366] = issue_pkt_r_instr_metadata__pc__52_;
  assign dispatch_pkt[367] = issue_pkt_r_instr_metadata__pc__53_;
  assign dispatch_pkt[368] = issue_pkt_r_instr_metadata__pc__54_;
  assign dispatch_pkt[369] = issue_pkt_r_instr_metadata__pc__55_;
  assign dispatch_pkt[370] = issue_pkt_r_instr_metadata__pc__56_;
  assign dispatch_pkt[371] = issue_pkt_r_instr_metadata__pc__57_;
  assign dispatch_pkt[372] = issue_pkt_r_instr_metadata__pc__58_;
  assign dispatch_pkt[373] = issue_pkt_r_instr_metadata__pc__59_;
  assign dispatch_pkt[374] = issue_pkt_r_instr_metadata__pc__60_;
  assign dispatch_pkt[375] = issue_pkt_r_instr_metadata__pc__61_;
  assign dispatch_pkt[376] = issue_pkt_r_instr_metadata__pc__62_;
  assign dispatch_pkt[377] = issue_pkt_r_instr_metadata__pc__63_;
  assign dispatch_pkt[378] = issue_pkt_r_instr_metadata__itag__0_;
  assign dispatch_pkt[379] = issue_pkt_r_instr_metadata__itag__1_;
  assign dispatch_pkt[380] = issue_pkt_r_instr_metadata__itag__2_;
  assign dispatch_pkt[381] = issue_pkt_r_instr_metadata__itag__3_;
  assign dispatch_pkt[382] = issue_pkt_r_instr_metadata__itag__4_;
  assign dispatch_pkt[383] = issue_pkt_r_instr_metadata__itag__5_;
  assign dispatch_pkt[384] = issue_pkt_r_instr_metadata__itag__6_;
  assign dispatch_pkt[385] = issue_pkt_r_instr_metadata__itag__7_;
  assign { N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9 } = (N0)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                                                                                                                                            (N1)? decoded : 1'b0;
  assign N0 = illegal_instr_isd;
  assign N1 = N8;
  assign dispatch_pkt[242:192] = (N2)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                 (N3)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                 (N4)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                 (N7)? { N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9 } : 1'b0;
  assign N2 = fe_nop_v;
  assign N3 = be_nop_v;
  assign N4 = me_nop_v;
  assign issue_pkt_ready_o = chk_dispatch_v_i | N60;
  assign N60 = ~calc_status_o[306];
  assign n_0_net_ = calc_stage_r_3__irf_w_v_ & N61;
  assign N61 = ~exc_stage_n_4__poison_v_;
  assign n_6_net_ = calc_stage_r_4__frf_w_v_ & N62;
  assign N62 = ~exc_stage_r_4__poison_v_;
  assign n_12_net_ = issue_pkt_v_i | chk_dispatch_v_i;
  assign n_28_net_ = N69 | exc_stage_r_0__cache_miss_v_;
  assign N69 = N68 | exc_stage_r_0__store_fault_v_;
  assign N68 = N67 | exc_stage_r_0__load_fault_v_;
  assign N67 = N66 | exc_stage_r_0__tlb_miss_v_;
  assign N66 = N65 | exc_stage_r_0__csr_instr_v_;
  assign N65 = N64 | exc_stage_r_0__ret_instr_v_;
  assign N64 = N63 | exc_stage_r_0__illegal_instr_v_;
  assign N63 = exc_stage_n_1__poison_v_ | exc_stage_n_1__roll_v_;
  assign fe_nop_v = N60 & chk_dispatch_v_i;
  assign be_nop_v = N70 & mmu_cmd_ready_i;
  assign N70 = ~chk_dispatch_v_i;
  assign me_nop_v = N71 & N72;
  assign N71 = ~chk_dispatch_v_i;
  assign N72 = ~mmu_cmd_ready_i;
  assign n_63_net_ = N74 & N75;
  assign N74 = calc_stage_r_2__instr_v_ & N73;
  assign N73 = ~exc_stage_n_3__poison_v_;
  assign N75 = ~exc_stage_n_3__cache_miss_v_;
  assign n_64_net_ = mtval_w_v_lo | calc_status_o[2];
  assign N5 = be_nop_v | fe_nop_v;
  assign N6 = me_nop_v | N5;
  assign N7 = ~N6;
  assign N8 = ~illegal_instr_isd;
  assign calc_status_o[189] = N76 | dispatch_pkt_r_decode__jmp_v_;
  assign N76 = dispatch_pkt_r_decode__br_v_ & pipe_int_data_lo[0];
  assign calc_status_o[190] = dispatch_pkt_r_decode__br_v_ | dispatch_pkt_r_decode__jmp_v_;
  assign calc_status_o[79] = N78 & calc_stage_r_0__irf_w_v_;
  assign N78 = calc_stage_r_0__pipe_int_v_ & N77;
  assign N77 = ~exc_stage_n_1__poison_v_;
  assign calc_status_o[78] = N80 & calc_stage_r_0__irf_w_v_;
  assign N80 = calc_stage_r_0__pipe_mul_v_ & N79;
  assign N79 = ~exc_stage_n_1__poison_v_;
  assign calc_status_o[77] = N82 & calc_stage_r_0__irf_w_v_;
  assign N82 = calc_stage_r_0__pipe_mem_v_ & N81;
  assign N81 = ~exc_stage_n_1__poison_v_;
  assign calc_status_o[76] = N84 & calc_stage_r_0__frf_w_v_;
  assign N84 = calc_stage_r_0__pipe_mem_v_ & N83;
  assign N83 = ~exc_stage_n_1__poison_v_;
  assign calc_status_o[75] = N86 & calc_stage_r_0__frf_w_v_;
  assign N86 = calc_stage_r_0__pipe_fp_v_ & N85;
  assign N85 = ~exc_stage_n_1__poison_v_;
  assign calc_status_o[74] = exc_stage_r_0__csr_instr_v_ | exc_stage_r_0__ret_instr_v_;
  assign calc_status_o[90] = N88 & calc_stage_r_1__irf_w_v_;
  assign N88 = calc_stage_r_1__pipe_int_v_ & N87;
  assign N87 = ~exc_stage_n_2__poison_v_;
  assign calc_status_o[89] = N90 & calc_stage_r_1__irf_w_v_;
  assign N90 = calc_stage_r_1__pipe_mul_v_ & N89;
  assign N89 = ~exc_stage_n_2__poison_v_;
  assign calc_status_o[88] = N92 & calc_stage_r_1__irf_w_v_;
  assign N92 = calc_stage_r_1__pipe_mem_v_ & N91;
  assign N91 = ~exc_stage_n_2__poison_v_;
  assign calc_status_o[87] = N94 & calc_stage_r_1__frf_w_v_;
  assign N94 = calc_stage_r_1__pipe_mem_v_ & N93;
  assign N93 = ~exc_stage_n_2__poison_v_;
  assign calc_status_o[86] = N96 & calc_stage_r_1__frf_w_v_;
  assign N96 = calc_stage_r_1__pipe_fp_v_ & N95;
  assign N95 = ~exc_stage_n_2__poison_v_;
  assign calc_status_o[85] = exc_stage_r_1__csr_instr_v_ | exc_stage_r_1__ret_instr_v_;
  assign calc_status_o[101] = N98 & calc_stage_r_2__irf_w_v_;
  assign N98 = calc_stage_r_2__pipe_int_v_ & N97;
  assign N97 = ~exc_stage_n_3__poison_v_;
  assign calc_status_o[100] = N100 & calc_stage_r_2__irf_w_v_;
  assign N100 = calc_stage_r_2__pipe_mul_v_ & N99;
  assign N99 = ~exc_stage_n_3__poison_v_;
  assign calc_status_o[99] = N102 & calc_stage_r_2__irf_w_v_;
  assign N102 = calc_stage_r_2__pipe_mem_v_ & N101;
  assign N101 = ~exc_stage_n_3__poison_v_;
  assign calc_status_o[98] = N104 & calc_stage_r_2__frf_w_v_;
  assign N104 = calc_stage_r_2__pipe_mem_v_ & N103;
  assign N103 = ~exc_stage_n_3__poison_v_;
  assign calc_status_o[97] = N106 & calc_stage_r_2__frf_w_v_;
  assign N106 = calc_stage_r_2__pipe_fp_v_ & N105;
  assign N105 = ~exc_stage_n_3__poison_v_;
  assign calc_status_o[96] = exc_stage_r_2__csr_instr_v_ | exc_stage_r_2__ret_instr_v_;
  assign calc_status_o[112] = N108 & calc_stage_r_3__irf_w_v_;
  assign N108 = calc_stage_r_3__pipe_int_v_ & N107;
  assign N107 = ~exc_stage_n_4__poison_v_;
  assign calc_status_o[111] = N110 & calc_stage_r_3__irf_w_v_;
  assign N110 = calc_stage_r_3__pipe_mul_v_ & N109;
  assign N109 = ~exc_stage_n_4__poison_v_;
  assign calc_status_o[110] = N112 & calc_stage_r_3__irf_w_v_;
  assign N112 = calc_stage_r_3__pipe_mem_v_ & N111;
  assign N111 = ~exc_stage_n_4__poison_v_;
  assign calc_status_o[109] = N114 & calc_stage_r_3__frf_w_v_;
  assign N114 = calc_stage_r_3__pipe_mem_v_ & N113;
  assign N113 = ~exc_stage_n_4__poison_v_;
  assign calc_status_o[108] = N116 & calc_stage_r_3__frf_w_v_;
  assign N116 = calc_stage_r_3__pipe_fp_v_ & N115;
  assign N115 = ~exc_stage_n_4__poison_v_;
  assign calc_status_o[107] = exc_stage_r_3__csr_instr_v_ | exc_stage_r_3__ret_instr_v_;
  assign calc_status_o[123] = N118 & calc_stage_r_4__irf_w_v_;
  assign N118 = calc_stage_r_4__pipe_int_v_ & N117;
  assign N117 = ~1'b0;
  assign calc_status_o[122] = N120 & calc_stage_r_4__irf_w_v_;
  assign N120 = calc_stage_r_4__pipe_mul_v_ & N119;
  assign N119 = ~1'b0;
  assign calc_status_o[121] = N122 & calc_stage_r_4__irf_w_v_;
  assign N122 = calc_stage_r_4__pipe_mem_v_ & N121;
  assign N121 = ~1'b0;
  assign calc_status_o[120] = N124 & calc_stage_r_4__frf_w_v_;
  assign N124 = calc_stage_r_4__pipe_mem_v_ & N123;
  assign N123 = ~1'b0;
  assign calc_status_o[119] = N126 & calc_stage_r_4__frf_w_v_;
  assign N126 = calc_stage_r_4__pipe_fp_v_ & N125;
  assign N125 = ~1'b0;
  assign calc_status_o[118] = exc_stage_r_4__csr_instr_v_ | exc_stage_r_4__ret_instr_v_;
  assign calc_status_o[68] = calc_stage_r_2__pipe_mem_v_ & N127;
  assign N127 = ~exc_stage_n_3__poison_v_;
  assign calc_status_o[3] = N128 & N129;
  assign N128 = exc_stage_n_3__cache_miss_v_ & calc_stage_r_2__pipe_mem_v_;
  assign N129 = ~exc_stage_r_2__poison_v_;
  assign calc_status_o[2] = exc_stage_r_2__illegal_instr_v_ & N129;
  assign calc_status_o[1] = exc_stage_r_2__ret_instr_v_ & N129;
  assign calc_status_o[0] = calc_stage_r_2__instr_v_ & N130;
  assign N130 = ~exc_stage_r_2__roll_v_;
  assign comp_stage_n_slice_iwb_v[1] = calc_stage_r_0__irf_w_v_ & N131;
  assign N131 = ~exc_stage_n_1__poison_v_;
  assign comp_stage_n_slice_fwb_v[1] = calc_stage_r_0__frf_w_v_ & N132;
  assign N132 = ~exc_stage_n_1__poison_v_;
  assign comp_stage_n_slice_iwb_v[2] = calc_stage_r_1__irf_w_v_ & N133;
  assign N133 = ~exc_stage_n_2__poison_v_;
  assign comp_stage_n_slice_fwb_v[2] = calc_stage_r_1__frf_w_v_ & N134;
  assign N134 = ~exc_stage_n_2__poison_v_;
  assign comp_stage_n_slice_iwb_v[3] = calc_stage_r_2__irf_w_v_ & N135;
  assign N135 = ~exc_stage_n_3__poison_v_;
  assign comp_stage_n_slice_fwb_v[3] = calc_stage_r_2__frf_w_v_ & N136;
  assign N136 = ~exc_stage_n_3__poison_v_;
  assign comp_stage_n_slice_iwb_v[4] = calc_stage_r_3__irf_w_v_ & N137;
  assign N137 = ~exc_stage_n_4__poison_v_;
  assign comp_stage_n_slice_fwb_v[4] = calc_stage_r_3__frf_w_v_ & N138;
  assign N138 = ~exc_stage_n_4__poison_v_;
  assign exc_stage_n_0__illegal_instr_v_ = dispatch_pkt[242] & illegal_instr_isd;
  assign exc_stage_n_1__roll_v_ = exc_stage_r_0__roll_v_ | chk_roll_i;
  assign exc_stage_n_2__roll_v_ = exc_stage_r_1__roll_v_ | chk_roll_i;
  assign exc_stage_n_3__roll_v_ = exc_stage_r_2__roll_v_ | chk_roll_i;
  assign exc_stage_n_1__poison_v_ = exc_stage_r_0__poison_v_ | chk_poison_ex1_i;
  assign exc_stage_n_2__poison_v_ = exc_stage_r_1__poison_v_ | chk_poison_ex2_i;
  assign exc_stage_n_3__poison_v_ = exc_stage_r_2__poison_v_ | chk_poison_ex3_i;

endmodule



module bp_be_dcache_wbuf_queue_width_p97
(
  clk_i,
  data_i,
  el0_en_i,
  el1_en_i,
  mux0_sel_i,
  mux1_sel_i,
  el0_snoop_o,
  el1_snoop_o,
  data_o
);

  input [96:0] data_i;
  output [96:0] el0_snoop_o;
  output [96:0] el1_snoop_o;
  output [96:0] data_o;
  input clk_i;
  input el0_en_i;
  input el1_en_i;
  input mux0_sel_i;
  input mux1_sel_i;
  wire [96:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102;
  reg [96:0] el0_snoop_o,el1_snoop_o;
  assign { N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5 } = (N0)? el0_snoop_o :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                (N1)? data_i : 1'b0;
  assign N0 = mux0_sel_i;
  assign N1 = N4;
  assign data_o = (N2)? el1_snoop_o :
                  (N3)? data_i : 1'b0;
  assign N2 = mux1_sel_i;
  assign N3 = N102;
  assign N4 = ~mux0_sel_i;
  assign N102 = ~mux1_sel_i;

  always @(posedge clk_i) begin
    if(el0_en_i) begin
      { el0_snoop_o[96:0] } <= { data_i[96:0] };
    end
    if(el1_en_i) begin
      { el1_snoop_o[96:0] } <= { N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5 };
    end
  end


endmodule



module bsg_mux_segmented_segments_p8_segment_width_p8
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [63:0] data0_i;
  input [63:0] data1_i;
  input [7:0] sel_i;
  output [63:0] data_o;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15;
  assign data_o[7:0] = (N0)? data1_i[7:0] :
                       (N8)? data0_i[7:0] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[15:8] = (N1)? data1_i[15:8] :
                        (N9)? data0_i[15:8] : 1'b0;
  assign N1 = sel_i[1];
  assign data_o[23:16] = (N2)? data1_i[23:16] :
                         (N10)? data0_i[23:16] : 1'b0;
  assign N2 = sel_i[2];
  assign data_o[31:24] = (N3)? data1_i[31:24] :
                         (N11)? data0_i[31:24] : 1'b0;
  assign N3 = sel_i[3];
  assign data_o[39:32] = (N4)? data1_i[39:32] :
                         (N12)? data0_i[39:32] : 1'b0;
  assign N4 = sel_i[4];
  assign data_o[47:40] = (N5)? data1_i[47:40] :
                         (N13)? data0_i[47:40] : 1'b0;
  assign N5 = sel_i[5];
  assign data_o[55:48] = (N6)? data1_i[55:48] :
                         (N14)? data0_i[55:48] : 1'b0;
  assign N6 = sel_i[6];
  assign data_o[63:56] = (N7)? data1_i[63:56] :
                         (N15)? data0_i[63:56] : 1'b0;
  assign N7 = sel_i[7];
  assign N8 = ~sel_i[0];
  assign N9 = ~sel_i[1];
  assign N10 = ~sel_i[2];
  assign N11 = ~sel_i[3];
  assign N12 = ~sel_i[4];
  assign N13 = ~sel_i[5];
  assign N14 = ~sel_i[6];
  assign N15 = ~sel_i[7];

endmodule



module bp_be_dcache_wbuf_data_width_p64_paddr_width_p22_ways_p8_sets_p64
(
  clk_i,
  reset_i,
  v_i,
  wbuf_entry_i,
  yumi_i,
  v_o,
  wbuf_entry_o,
  empty_o,
  bypass_addr_i,
  bypass_v_i,
  bypass_data_o,
  bypass_mask_o,
  lce_snoop_index_i,
  lce_snoop_way_i,
  lce_snoop_match_o
);

  input [96:0] wbuf_entry_i;
  output [96:0] wbuf_entry_o;
  input [21:0] bypass_addr_i;
  output [63:0] bypass_data_o;
  output [7:0] bypass_mask_o;
  input [5:0] lce_snoop_index_i;
  input [2:0] lce_snoop_way_i;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input bypass_v_i;
  output v_o;
  output empty_o;
  output lce_snoop_match_o;
  wire [96:0] wbuf_entry_o,wbuf_entry_el0,wbuf_entry_el1;
  wire v_o,empty_o,lce_snoop_match_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,
  el0_valid,el1_valid,el0_enable,N14,el1_enable,mux0_sel,mux1_sel,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,tag_hit0_n,tag_hit1_n,tag_hit2_n,n_2_net__7_,
  n_2_net__6_,n_2_net__5_,n_2_net__4_,n_2_net__3_,n_2_net__2_,n_2_net__1_,n_2_net__0_,
  n_4_net__7_,n_4_net__6_,n_4_net__5_,n_4_net__4_,n_4_net__3_,n_4_net__2_,n_4_net__1_,
  n_4_net__0_,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,
  N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,
  N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,
  N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,
  N103,N104,lce_snoop_el2_match,N105,N106,lce_snoop_el0_match,N107,N108,
  lce_snoop_el1_match,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,
  N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,
  N139,N140,N141,N142,N143,N144,N145;
  wire [7:7] tag_hit0x4,tag_hit1x4,tag_hit2x4;
  wire [7:0] bypass_mask_n;
  wire [63:0] el0or1_data,bypass_data_n;
  reg [1:0] num_els_r;
  reg [63:0] bypass_data_o;
  reg [7:0] bypass_mask_o;
  assign N8 = N6 & N7;
  assign N9 = num_els_r[1] | N7;
  assign N11 = N6 | num_els_r[0];
  assign N13 = num_els_r[1] & num_els_r[0];

  bp_be_dcache_wbuf_queue_width_p97
  wbq
  (
    .clk_i(clk_i),
    .data_i(wbuf_entry_i),
    .el0_en_i(el0_enable),
    .el1_en_i(el1_enable),
    .mux0_sel_i(mux0_sel),
    .mux1_sel_i(mux1_sel),
    .el0_snoop_o(wbuf_entry_el0),
    .el1_snoop_o(wbuf_entry_el1),
    .data_o(wbuf_entry_o)
  );

  assign tag_hit0_n = bypass_addr_i[21:3] == wbuf_entry_el0[96:78];
  assign tag_hit1_n = bypass_addr_i[21:3] == wbuf_entry_el1[96:78];
  assign tag_hit2_n = bypass_addr_i[21:3] == wbuf_entry_i[96:78];

  bsg_mux_segmented_segments_p8_segment_width_p8
  mux_segmented_merge0
  (
    .data0_i(wbuf_entry_el1[74:11]),
    .data1_i(wbuf_entry_el0[74:11]),
    .sel_i({ n_2_net__7_, n_2_net__6_, n_2_net__5_, n_2_net__4_, n_2_net__3_, n_2_net__2_, n_2_net__1_, n_2_net__0_ }),
    .data_o(el0or1_data)
  );


  bsg_mux_segmented_segments_p8_segment_width_p8
  mux_segmented_merge1
  (
    .data0_i(el0or1_data),
    .data1_i(wbuf_entry_i[74:11]),
    .sel_i({ n_4_net__7_, n_4_net__6_, n_4_net__5_, n_4_net__4_, n_4_net__3_, n_4_net__2_, n_4_net__1_, n_4_net__0_ }),
    .data_o(bypass_data_n)
  );

  assign N103 = lce_snoop_index_i == wbuf_entry_i[86:81];
  assign N104 = lce_snoop_way_i == wbuf_entry_i[2:0];
  assign N105 = lce_snoop_index_i == wbuf_entry_el0[86:81];
  assign N106 = lce_snoop_way_i == wbuf_entry_el0[2:0];
  assign N107 = lce_snoop_index_i == wbuf_entry_el1[86:81];
  assign N108 = lce_snoop_way_i == wbuf_entry_el1[2:0];
  assign { N21, N20 } = v_i - N19;
  assign { N23, N22 } = num_els_r + { N21, N20 };
  assign v_o = (N0)? v_i :
               (N1)? 1'b1 :
               (N2)? 1'b1 :
               (N3)? 1'b0 : 1'b0;
  assign N0 = N8;
  assign N1 = N10;
  assign N2 = N12;
  assign N3 = N13;
  assign empty_o = (N0)? 1'b1 :
                   (N1)? 1'b0 :
                   (N2)? 1'b0 :
                   (N3)? 1'b0 : 1'b0;
  assign el0_valid = (N0)? 1'b0 :
                     (N1)? 1'b0 :
                     (N2)? 1'b1 :
                     (N3)? 1'b0 : 1'b0;
  assign el1_valid = (N0)? 1'b0 :
                     (N1)? 1'b1 :
                     (N2)? 1'b1 :
                     (N3)? 1'b0 : 1'b0;
  assign el0_enable = (N0)? 1'b0 :
                      (N1)? N15 :
                      (N2)? N17 :
                      (N3)? 1'b0 : 1'b0;
  assign el1_enable = (N0)? N14 :
                      (N1)? N16 :
                      (N2)? yumi_i :
                      (N3)? 1'b0 : 1'b0;
  assign mux0_sel = (N0)? 1'b0 :
                    (N1)? 1'b0 :
                    (N2)? 1'b1 :
                    (N3)? 1'b0 : 1'b0;
  assign mux1_sel = (N0)? 1'b0 :
                    (N1)? 1'b1 :
                    (N2)? 1'b1 :
                    (N3)? 1'b0 : 1'b0;
  assign { N25, N24 } = (N4)? { 1'b0, 1'b0 } :
                        (N5)? { N23, N22 } : 1'b0;
  assign N4 = reset_i;
  assign N5 = N18;
  assign N28 = (N4)? 1'b1 :
               (N102)? 1'b1 :
               (N27)? 1'b0 : 1'b0;
  assign { N36, N35, N34, N33, N32, N31, N30, N29 } = (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                      (N102)? bypass_mask_n : 1'b0;
  assign { N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37 } = (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                                                                                                                                                                                                               (N102)? bypass_data_n : 1'b0;
  assign N6 = ~num_els_r[1];
  assign N7 = ~num_els_r[0];
  assign N10 = ~N9;
  assign N12 = ~N11;
  assign N14 = v_i & N109;
  assign N109 = ~yumi_i;
  assign N15 = v_i & N109;
  assign N16 = v_i & yumi_i;
  assign N17 = v_i & yumi_i;
  assign N18 = ~reset_i;
  assign N19 = v_o & yumi_i;
  assign tag_hit0x4[7] = tag_hit0_n & el0_valid;
  assign tag_hit1x4[7] = tag_hit1_n & el1_valid;
  assign tag_hit2x4[7] = tag_hit2_n & v_i;
  assign bypass_mask_n[7] = N112 | N113;
  assign N112 = N110 | N111;
  assign N110 = tag_hit0x4[7] & wbuf_entry_el0[10];
  assign N111 = tag_hit1x4[7] & wbuf_entry_el1[10];
  assign N113 = tag_hit2x4[7] & wbuf_entry_i[10];
  assign bypass_mask_n[6] = N116 | N117;
  assign N116 = N114 | N115;
  assign N114 = tag_hit0x4[7] & wbuf_entry_el0[9];
  assign N115 = tag_hit1x4[7] & wbuf_entry_el1[9];
  assign N117 = tag_hit2x4[7] & wbuf_entry_i[9];
  assign bypass_mask_n[5] = N120 | N121;
  assign N120 = N118 | N119;
  assign N118 = tag_hit0x4[7] & wbuf_entry_el0[8];
  assign N119 = tag_hit1x4[7] & wbuf_entry_el1[8];
  assign N121 = tag_hit2x4[7] & wbuf_entry_i[8];
  assign bypass_mask_n[4] = N124 | N125;
  assign N124 = N122 | N123;
  assign N122 = tag_hit0x4[7] & wbuf_entry_el0[7];
  assign N123 = tag_hit1x4[7] & wbuf_entry_el1[7];
  assign N125 = tag_hit2x4[7] & wbuf_entry_i[7];
  assign bypass_mask_n[3] = N128 | N129;
  assign N128 = N126 | N127;
  assign N126 = tag_hit0x4[7] & wbuf_entry_el0[6];
  assign N127 = tag_hit1x4[7] & wbuf_entry_el1[6];
  assign N129 = tag_hit2x4[7] & wbuf_entry_i[6];
  assign bypass_mask_n[2] = N132 | N133;
  assign N132 = N130 | N131;
  assign N130 = tag_hit0x4[7] & wbuf_entry_el0[5];
  assign N131 = tag_hit1x4[7] & wbuf_entry_el1[5];
  assign N133 = tag_hit2x4[7] & wbuf_entry_i[5];
  assign bypass_mask_n[1] = N136 | N137;
  assign N136 = N134 | N135;
  assign N134 = tag_hit0x4[7] & wbuf_entry_el0[4];
  assign N135 = tag_hit1x4[7] & wbuf_entry_el1[4];
  assign N137 = tag_hit2x4[7] & wbuf_entry_i[4];
  assign bypass_mask_n[0] = N140 | N141;
  assign N140 = N138 | N139;
  assign N138 = tag_hit0x4[7] & wbuf_entry_el0[3];
  assign N139 = tag_hit1x4[7] & wbuf_entry_el1[3];
  assign N141 = tag_hit2x4[7] & wbuf_entry_i[3];
  assign n_2_net__7_ = tag_hit0x4[7] & wbuf_entry_el0[10];
  assign n_2_net__6_ = tag_hit0x4[7] & wbuf_entry_el0[9];
  assign n_2_net__5_ = tag_hit0x4[7] & wbuf_entry_el0[8];
  assign n_2_net__4_ = tag_hit0x4[7] & wbuf_entry_el0[7];
  assign n_2_net__3_ = tag_hit0x4[7] & wbuf_entry_el0[6];
  assign n_2_net__2_ = tag_hit0x4[7] & wbuf_entry_el0[5];
  assign n_2_net__1_ = tag_hit0x4[7] & wbuf_entry_el0[4];
  assign n_2_net__0_ = tag_hit0x4[7] & wbuf_entry_el0[3];
  assign n_4_net__7_ = tag_hit2x4[7] & wbuf_entry_i[10];
  assign n_4_net__6_ = tag_hit2x4[7] & wbuf_entry_i[9];
  assign n_4_net__5_ = tag_hit2x4[7] & wbuf_entry_i[8];
  assign n_4_net__4_ = tag_hit2x4[7] & wbuf_entry_i[7];
  assign n_4_net__3_ = tag_hit2x4[7] & wbuf_entry_i[6];
  assign n_4_net__2_ = tag_hit2x4[7] & wbuf_entry_i[5];
  assign n_4_net__1_ = tag_hit2x4[7] & wbuf_entry_i[4];
  assign n_4_net__0_ = tag_hit2x4[7] & wbuf_entry_i[3];
  assign N26 = bypass_v_i | reset_i;
  assign N27 = ~N26;
  assign N101 = ~reset_i;
  assign N102 = bypass_v_i & N101;
  assign lce_snoop_el2_match = N142 & N104;
  assign N142 = v_i & N103;
  assign lce_snoop_el0_match = N143 & N106;
  assign N143 = el0_valid & N105;
  assign lce_snoop_el1_match = N144 & N108;
  assign N144 = el1_valid & N107;
  assign lce_snoop_match_o = N145 | lce_snoop_el1_match;
  assign N145 = lce_snoop_el2_match | lce_snoop_el0_match;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { num_els_r[1:0] } <= { N25, N24 };
    end
    if(N28) begin
      { bypass_data_o[63:0] } <= { N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37 };
      { bypass_mask_o[7:0] } <= { N36, N35, N34, N33, N32, N31, N30, N29 };
    end
  end


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p15_els_p64
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [14:0] data_i;
  input [5:0] addr_i;
  input [14:0] w_mask_i;
  output [14:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [14:0] data_o;

  hard_mem_1rw_bit_mask_d64_w15_wrapper
  macro_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bp_be_dcache_lce_req_data_width_p64_paddr_width_p22_num_cce_p1_num_lce_p2_ways_p8
(
  clk_i,
  reset_i,
  lce_id_i,
  load_miss_i,
  store_miss_i,
  miss_addr_i,
  lru_way_i,
  dirty_i,
  uncached_load_req_i,
  uncached_store_req_i,
  store_data_i,
  size_op_i,
  cache_miss_o,
  miss_addr_o,
  tr_data_received_i,
  cce_data_received_i,
  uncached_data_received_i,
  set_tag_received_i,
  set_tag_wakeup_received_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_yumi_i
);

  input [0:0] lce_id_i;
  input [21:0] miss_addr_i;
  input [2:0] lru_way_i;
  input [7:0] dirty_i;
  input [63:0] store_data_i;
  input [1:0] size_op_i;
  output [21:0] miss_addr_o;
  output [96:0] lce_req_o;
  output [25:0] lce_resp_o;
  input clk_i;
  input reset_i;
  input load_miss_i;
  input store_miss_i;
  input uncached_load_req_i;
  input uncached_store_req_i;
  input tr_data_received_i;
  input cce_data_received_i;
  input uncached_data_received_i;
  input set_tag_received_i;
  input set_tag_wakeup_received_i;
  input lce_req_ready_i;
  input lce_resp_yumi_i;
  output cache_miss_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  wire [96:0] lce_req_o;
  wire [25:0] lce_resp_o;
  wire cache_miss_o,lce_req_v_o,lce_resp_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,
  tr_data_received,cce_data_received,set_tag_received,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,dirty_lru_flopped_n,tr_data_received_n,
  cce_data_received_n,set_tag_received_n,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256;
  wire [2:0] state_n;
  reg size_op_r,dirty_lru_flopped_r,tr_data_received_r,cce_data_received_r,
  set_tag_received_r,load_not_store_r,dirty_r;
  reg [2:0] state_r,lru_way_r;
  reg [21:0] miss_addr_o;
  assign lce_resp_o[23] = 1'b1;
  assign lce_resp_o[25] = 1'b0;
  assign lce_req_o[29] = 1'b0;
  assign lce_req_o[32] = 1'b0;
  assign lce_resp_o[21] = miss_addr_o[21];
  assign lce_resp_o[20] = miss_addr_o[20];
  assign lce_resp_o[19] = miss_addr_o[19];
  assign lce_resp_o[18] = miss_addr_o[18];
  assign lce_resp_o[17] = miss_addr_o[17];
  assign lce_resp_o[16] = miss_addr_o[16];
  assign lce_resp_o[15] = miss_addr_o[15];
  assign lce_resp_o[14] = miss_addr_o[14];
  assign lce_resp_o[13] = miss_addr_o[13];
  assign lce_resp_o[12] = miss_addr_o[12];
  assign lce_resp_o[11] = miss_addr_o[11];
  assign lce_resp_o[10] = miss_addr_o[10];
  assign lce_resp_o[9] = miss_addr_o[9];
  assign lce_resp_o[8] = miss_addr_o[8];
  assign lce_resp_o[7] = miss_addr_o[7];
  assign lce_resp_o[6] = miss_addr_o[6];
  assign lce_resp_o[5] = miss_addr_o[5];
  assign lce_resp_o[4] = miss_addr_o[4];
  assign lce_resp_o[3] = miss_addr_o[3];
  assign lce_resp_o[2] = miss_addr_o[2];
  assign lce_resp_o[1] = miss_addr_o[1];
  assign lce_resp_o[0] = miss_addr_o[0];
  assign lce_resp_o[24] = lce_id_i[0];
  assign lce_req_o[31] = lce_id_i[0];
  assign N28 = (N20)? dirty_i[0] :
               (N22)? dirty_i[1] :
               (N24)? dirty_i[2] :
               (N26)? dirty_i[3] :
               (N21)? dirty_i[4] :
               (N23)? dirty_i[5] :
               (N25)? dirty_i[6] :
               (N27)? dirty_i[7] : 1'b0;
  assign N32 = N29 & N30;
  assign N33 = N32 & N31;
  assign N34 = state_r[2] | state_r[1];
  assign N35 = N34 | N31;
  assign N37 = state_r[2] | N30;
  assign N38 = N37 | state_r[0];
  assign N40 = N29 | state_r[1];
  assign N41 = N40 | N31;
  assign N43 = state_r[2] | N30;
  assign N44 = N43 | N31;
  assign N46 = N29 | state_r[1];
  assign N47 = N46 | state_r[0];
  assign N49 = state_r[2] & state_r[1];
  assign lce_req_o[6:4] = (N0)? lru_way_r :
                          (N1)? lru_way_i : 1'b0;
  assign N0 = dirty_lru_flopped_r;
  assign N1 = N12;
  assign lce_req_o[3] = (N0)? dirty_r :
                        (N1)? N28 : 1'b0;
  assign N57 = (N2)? 1'b1 :
               (N167)? 1'b1 :
               (N170)? N54 :
               (N53)? 1'b0 : 1'b0;
  assign N2 = N50;
  assign { N59, N58 } = (N2)? { 1'b0, 1'b1 } :
                        (N167)? { 1'b1, 1'b0 } :
                        (N170)? { 1'b0, 1'b0 } :
                        (N53)? { 1'b0, 1'b0 } : 1'b0;
  assign N60 = (N2)? 1'b0 :
               (N167)? 1'b0 :
               (N170)? 1'b1 :
               (N53)? 1'b0 : 1'b0;
  assign { N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61 } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, miss_addr_o } :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           (N167)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, miss_addr_o } :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           (N170)? { store_data_i, miss_addr_i } :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           (N53)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, miss_addr_o } : 1'b0;
  assign { N158, N157, N156 } = (N3)? { 1'b0, 1'b1, 1'b1 } :
                                (N174)? { 1'b1, 1'b0, 1'b0 } :
                                (N155)? { 1'b1, 1'b0, 1'b1 } : 1'b0;
  assign N3 = tr_data_received;
  assign { N161, N160, N159 } = (N4)? { 1'b0, 1'b0, 1'b0 } :
                                (N172)? { N158, N157, N156 } :
                                (N153)? { 1'b1, 1'b0, 1'b1 } : 1'b0;
  assign N4 = N151;
  assign lce_req_o[1:0] = (N5)? { 1'b0, size_op_r } :
                          (N163)? size_op_i : 1'b0;
  assign N5 = N39;
  assign lce_req_o[2] = (N6)? N60 :
                        (N7)? 1'b0 :
                        (N5)? 1'b1 :
                        (N8)? 1'b0 :
                        (N9)? 1'b0 :
                        (N10)? 1'b0 :
                        (N11)? 1'b0 : 1'b0;
  assign N6 = N33;
  assign N7 = N36;
  assign N8 = N42;
  assign N9 = N45;
  assign N10 = N48;
  assign N11 = N49;
  assign { lce_req_o[96:33], lce_req_o[28:7] } = (N6)? { N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61 } :
                                                 (N165)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, miss_addr_o } : 1'b0;
  assign lce_req_o[30] = (N7)? N147 :
                         (N166)? 1'b0 : 1'b0;
  assign dirty_lru_flopped_n = (N6)? 1'b0 :
                               (N7)? 1'b1 : 1'b0;
  assign tr_data_received_n = (N6)? 1'b0 :
                              (N8)? 1'b1 : 1'b0;
  assign cce_data_received_n = (N6)? 1'b0 :
                               (N8)? 1'b1 : 1'b0;
  assign set_tag_received_n = (N6)? 1'b0 :
                              (N8)? 1'b1 : 1'b0;
  assign cache_miss_o = (N6)? N57 :
                        (N7)? 1'b1 :
                        (N5)? 1'b1 :
                        (N8)? 1'b1 :
                        (N9)? 1'b1 :
                        (N10)? 1'b1 :
                        (N11)? 1'b0 : 1'b0;
  assign state_n = (N6)? { 1'b0, N59, N58 } :
                   (N7)? { lce_req_ready_i, 1'b0, 1'b1 } :
                   (N5)? { lce_req_ready_i, N54, lce_req_ready_i } :
                   (N8)? { N161, N160, N159 } :
                   (N9)? { 1'b0, N162, N162 } :
                   (N10)? { N162, 1'b0, 1'b0 } :
                   (N11)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_req_v_o = (N6)? N60 :
                       (N7)? 1'b1 :
                       (N5)? 1'b1 :
                       (N8)? 1'b0 :
                       (N9)? 1'b0 :
                       (N10)? 1'b0 :
                       (N11)? 1'b0 : 1'b0;
  assign lce_resp_v_o = (N6)? 1'b0 :
                        (N7)? 1'b0 :
                        (N5)? 1'b0 :
                        (N8)? 1'b0 :
                        (N9)? 1'b1 :
                        (N10)? 1'b1 :
                        (N11)? 1'b0 : 1'b0;
  assign lce_resp_o[22] = (N6)? 1'b0 :
                          (N7)? 1'b0 :
                          (N5)? 1'b0 :
                          (N8)? 1'b0 :
                          (N9)? 1'b0 :
                          (N10)? 1'b1 :
                          (N11)? 1'b0 : 1'b0;
  assign tr_data_received = tr_data_received_r | tr_data_received_i;
  assign cce_data_received = cce_data_received_r | cce_data_received_i;
  assign set_tag_received = set_tag_received_r | set_tag_received_i;
  assign N12 = ~dirty_lru_flopped_r;
  assign N13 = ~lru_way_i[0];
  assign N14 = ~lru_way_i[1];
  assign N15 = N13 & N14;
  assign N16 = N13 & lru_way_i[1];
  assign N17 = lru_way_i[0] & N14;
  assign N18 = lru_way_i[0] & lru_way_i[1];
  assign N19 = ~lru_way_i[2];
  assign N20 = N15 & N19;
  assign N21 = N15 & lru_way_i[2];
  assign N22 = N17 & N19;
  assign N23 = N17 & lru_way_i[2];
  assign N24 = N16 & N19;
  assign N25 = N16 & lru_way_i[2];
  assign N26 = N18 & N19;
  assign N27 = N18 & lru_way_i[2];
  assign N29 = ~state_r[2];
  assign N30 = ~state_r[1];
  assign N31 = ~state_r[0];
  assign N36 = ~N35;
  assign N39 = ~N38;
  assign N42 = ~N41;
  assign N45 = ~N44;
  assign N48 = ~N47;
  assign N50 = load_miss_i | store_miss_i;
  assign N51 = uncached_load_req_i | N50;
  assign N52 = uncached_store_req_i | N51;
  assign N53 = ~N52;
  assign N54 = ~lce_req_ready_i;
  assign N55 = ~N51;
  assign N56 = ~N50;
  assign N147 = ~load_not_store_r;
  assign N148 = ~tr_data_received_i;
  assign N149 = ~cce_data_received_i;
  assign N150 = ~set_tag_received_i;
  assign N151 = set_tag_wakeup_received_i | uncached_data_received_i;
  assign N152 = set_tag_received | N151;
  assign N153 = ~N152;
  assign N154 = cce_data_received | tr_data_received;
  assign N155 = ~N154;
  assign N162 = ~lce_resp_yumi_i;
  assign N163 = N38;
  assign N164 = ~N33;
  assign N165 = N164;
  assign N166 = N35;
  assign N167 = uncached_load_req_i & N56;
  assign N168 = ~uncached_load_req_i;
  assign N169 = N56 & N168;
  assign N170 = uncached_store_req_i & N169;
  assign N171 = ~N151;
  assign N172 = set_tag_received & N171;
  assign N173 = ~tr_data_received;
  assign N174 = cce_data_received & N173;
  assign N175 = ~reset_i;
  assign N176 = N33 & N175;
  assign N177 = N50 & N176;
  assign N178 = N55 & N176;
  assign N179 = N177 | N178;
  assign N180 = N36 & N175;
  assign N181 = N179 | N180;
  assign N182 = N39 & N175;
  assign N183 = N181 | N182;
  assign N184 = N42 & N175;
  assign N185 = N183 | N184;
  assign N186 = N45 & N175;
  assign N187 = N185 | N186;
  assign N188 = N48 & N175;
  assign N189 = N187 | N188;
  assign N190 = N49 & N175;
  assign N191 = N189 | N190;
  assign N192 = ~N191;
  assign N193 = N175 & N192;
  assign N194 = N56 & N33;
  assign N195 = N194 | N39;
  assign N196 = N195 | N42;
  assign N197 = N196 | N45;
  assign N198 = N197 | N48;
  assign N199 = N198 | N49;
  assign N200 = ~N199;
  assign N201 = N55 & N33;
  assign N202 = N201 | N36;
  assign N203 = N202 | N39;
  assign N204 = N148 & N42;
  assign N205 = N203 | N204;
  assign N206 = N205 | N45;
  assign N207 = N206 | N48;
  assign N208 = N207 | N49;
  assign N209 = ~N208;
  assign N210 = N149 & N42;
  assign N211 = N203 | N210;
  assign N212 = N211 | N45;
  assign N213 = N212 | N48;
  assign N214 = N213 | N49;
  assign N215 = ~N214;
  assign N216 = N150 & N42;
  assign N217 = N203 | N216;
  assign N218 = N217 | N45;
  assign N219 = N218 | N48;
  assign N220 = N219 | N49;
  assign N221 = ~N220;
  assign N222 = N56 & N176;
  assign N223 = N222 | N180;
  assign N224 = N223 | N182;
  assign N225 = N224 | N184;
  assign N226 = N225 | N186;
  assign N227 = N226 | N188;
  assign N228 = N227 | N190;
  assign N229 = ~N228;
  assign N230 = N175 & N229;
  assign N231 = dirty_lru_flopped_r & N180;
  assign N232 = N176 | N231;
  assign N233 = N232 | N182;
  assign N234 = N233 | N184;
  assign N235 = N234 | N186;
  assign N236 = N235 | N188;
  assign N237 = N236 | N190;
  assign N238 = ~N237;
  assign N239 = N175 & N238;
  assign N240 = dirty_lru_flopped_r & N180;
  assign N241 = N176 | N240;
  assign N242 = N241 | N182;
  assign N243 = N242 | N184;
  assign N244 = N243 | N186;
  assign N245 = N244 | N188;
  assign N246 = N245 | N190;
  assign N247 = ~N246;
  assign N248 = N175 & N247;
  assign N249 = N178 | N180;
  assign N250 = N249 | N182;
  assign N251 = N250 | N184;
  assign N252 = N251 | N186;
  assign N253 = N252 | N188;
  assign N254 = N253 | N190;
  assign N255 = ~N254;
  assign N256 = N175 & N255;

  always @(posedge clk_i) begin
    if(N193) begin
      size_op_r <= size_op_i[0];
    end
    if(reset_i) begin
      { state_r[2:0] } <= { 1'b0, 1'b0, 1'b0 };
    end else if(1'b1) begin
      { state_r[2:0] } <= { state_n[2:0] };
    end
    if(reset_i) begin
      dirty_lru_flopped_r <= 1'b0;
    end else if(N200) begin
      dirty_lru_flopped_r <= dirty_lru_flopped_n;
    end
    if(reset_i) begin
      tr_data_received_r <= 1'b0;
    end else if(N209) begin
      tr_data_received_r <= tr_data_received_n;
    end
    if(reset_i) begin
      cce_data_received_r <= 1'b0;
    end else if(N215) begin
      cce_data_received_r <= cce_data_received_n;
    end
    if(reset_i) begin
      set_tag_received_r <= 1'b0;
    end else if(N221) begin
      set_tag_received_r <= set_tag_received_n;
    end
    if(N230) begin
      load_not_store_r <= load_miss_i;
    end
    if(N239) begin
      { lru_way_r[2:0] } <= { lru_way_i[2:0] };
    end
    if(N248) begin
      dirty_r <= N28;
    end
    if(N256) begin
      { miss_addr_o[21:0] } <= { miss_addr_i[21:0] };
    end
  end


endmodule



module bp_be_dcache_lce_cmd_num_cce_p1_num_lce_p2_paddr_width_p22_lce_data_width_p512_sets_p64_ways_p8_data_width_p64
(
  clk_i,
  reset_i,
  lce_id_i,
  lce_sync_done_o,
  set_tag_received_o,
  set_tag_wakeup_received_o,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_yumi_o,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_yumi_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i,
  data_mem_pkt_v_o,
  data_mem_pkt_o,
  data_mem_data_i,
  data_mem_pkt_yumi_i,
  tag_mem_pkt_v_o,
  tag_mem_pkt_o,
  tag_mem_pkt_yumi_i,
  stat_mem_pkt_v_o,
  stat_mem_pkt_o,
  dirty_i,
  stat_mem_pkt_yumi_i
);

  input [0:0] lce_id_i;
  input [35:0] lce_cmd_i;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  output [517:0] lce_data_cmd_o;
  output [522:0] data_mem_pkt_o;
  input [511:0] data_mem_data_i;
  output [22:0] tag_mem_pkt_o;
  output [10:0] stat_mem_pkt_o;
  input [7:0] dirty_i;
  input clk_i;
  input reset_i;
  input lce_cmd_v_i;
  input lce_resp_yumi_i;
  input lce_data_resp_ready_i;
  input lce_data_cmd_ready_i;
  input data_mem_pkt_yumi_i;
  input tag_mem_pkt_yumi_i;
  input stat_mem_pkt_yumi_i;
  output lce_sync_done_o;
  output set_tag_received_o;
  output set_tag_wakeup_received_o;
  output lce_cmd_yumi_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_data_cmd_v_o;
  output data_mem_pkt_v_o;
  output tag_mem_pkt_v_o;
  output stat_mem_pkt_v_o;
  wire [25:0] lce_resp_o;
  wire [536:0] lce_data_resp_o;
  wire [517:0] lce_data_cmd_o;
  wire [522:0] data_mem_pkt_o;
  wire [22:0] tag_mem_pkt_o;
  wire [10:0] stat_mem_pkt_o;
  wire lce_sync_done_o,set_tag_received_o,set_tag_wakeup_received_o,lce_cmd_yumi_o,
  lce_resp_v_o,lce_data_resp_v_o,lce_data_cmd_v_o,data_mem_pkt_v_o,tag_mem_pkt_v_o,
  stat_mem_pkt_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,lce_tr_done,lce_data_resp_done,N28,N29,N30,
  N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,
  N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,
  N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,
  N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,
  N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,
  N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,
  N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,
  N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,
  N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,
  N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,
  N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,
  N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,
  N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,
  N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,
  N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,
  N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,
  N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,
  N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,
  N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
  N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,
  N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,
  N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,
  N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,
  N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,
  N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,
  N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,
  N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,
  N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,
  N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,
  N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,
  N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,
  N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,
  N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,
  N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,
  N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,
  N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,
  N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,
  N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,
  N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,
  N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,
  N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,
  N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,
  N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,
  N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,
  N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,
  N765,N766,N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,
  N781,N782,N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,
  N797,N798,N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,
  N813,N814,N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,
  N829,N830,N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
  N845,N846,N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,
  N861,N862,N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,
  N877,N878,N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,
  N893,N894,N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,
  N909,N910,N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,
  N925,N926,N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,
  N941,N942,N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,
  N957,N958,N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,
  N973,N974,N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,
  N989,N990,N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,
  N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,
  N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,
  N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,
  N1044,N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,
  N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,
  N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,
  N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,
  N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,
  N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,
  N1124,N1125,N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,
  N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,
  N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,
  N1164,N1165,N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,
  N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,
  N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,
  N1204,N1205,N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,
  N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,
  N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,
  N1244,N1245,N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,
  N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,
  N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,
  N1284,N1285,N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,
  N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,
  N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,
  N1324,N1325,N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,
  N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,
  N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,
  N1364,N1365,N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,
  N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,
  N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,
  N1404,N1405,N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,
  N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,
  N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,
  N1444,N1445,N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,
  N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,
  N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,
  N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,
  N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,
  N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,
  N1524,N1525,N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,
  N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,
  N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,
  N1564,N1565,N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,
  N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,
  N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,
  N1604,N1605,N1607,N1608;
  wire [2:0] state_n;
  reg [511:0] data_buf_r;
  reg [2:0] state_r;
  reg [0:0] sync_ack_count_r;
  reg tr_data_buffered_r,wb_data_buffered_r,wb_data_read_r,wb_dirty_cleared_r,
  invalidated_tag_r;
  assign data_mem_pkt_o[1] = 1'b0;
  assign data_mem_pkt_o[2] = 1'b0;
  assign data_mem_pkt_o[3] = 1'b0;
  assign data_mem_pkt_o[4] = 1'b0;
  assign data_mem_pkt_o[5] = 1'b0;
  assign data_mem_pkt_o[6] = 1'b0;
  assign data_mem_pkt_o[7] = 1'b0;
  assign data_mem_pkt_o[8] = 1'b0;
  assign data_mem_pkt_o[9] = 1'b0;
  assign data_mem_pkt_o[10] = 1'b0;
  assign data_mem_pkt_o[11] = 1'b0;
  assign data_mem_pkt_o[12] = 1'b0;
  assign data_mem_pkt_o[13] = 1'b0;
  assign data_mem_pkt_o[14] = 1'b0;
  assign data_mem_pkt_o[15] = 1'b0;
  assign data_mem_pkt_o[16] = 1'b0;
  assign data_mem_pkt_o[17] = 1'b0;
  assign data_mem_pkt_o[18] = 1'b0;
  assign data_mem_pkt_o[19] = 1'b0;
  assign data_mem_pkt_o[20] = 1'b0;
  assign data_mem_pkt_o[21] = 1'b0;
  assign data_mem_pkt_o[22] = 1'b0;
  assign data_mem_pkt_o[23] = 1'b0;
  assign data_mem_pkt_o[24] = 1'b0;
  assign data_mem_pkt_o[25] = 1'b0;
  assign data_mem_pkt_o[26] = 1'b0;
  assign data_mem_pkt_o[27] = 1'b0;
  assign data_mem_pkt_o[28] = 1'b0;
  assign data_mem_pkt_o[29] = 1'b0;
  assign data_mem_pkt_o[30] = 1'b0;
  assign data_mem_pkt_o[31] = 1'b0;
  assign data_mem_pkt_o[32] = 1'b0;
  assign data_mem_pkt_o[33] = 1'b0;
  assign data_mem_pkt_o[34] = 1'b0;
  assign data_mem_pkt_o[35] = 1'b0;
  assign data_mem_pkt_o[36] = 1'b0;
  assign data_mem_pkt_o[37] = 1'b0;
  assign data_mem_pkt_o[38] = 1'b0;
  assign data_mem_pkt_o[39] = 1'b0;
  assign data_mem_pkt_o[40] = 1'b0;
  assign data_mem_pkt_o[41] = 1'b0;
  assign data_mem_pkt_o[42] = 1'b0;
  assign data_mem_pkt_o[43] = 1'b0;
  assign data_mem_pkt_o[44] = 1'b0;
  assign data_mem_pkt_o[45] = 1'b0;
  assign data_mem_pkt_o[46] = 1'b0;
  assign data_mem_pkt_o[47] = 1'b0;
  assign data_mem_pkt_o[48] = 1'b0;
  assign data_mem_pkt_o[49] = 1'b0;
  assign data_mem_pkt_o[50] = 1'b0;
  assign data_mem_pkt_o[51] = 1'b0;
  assign data_mem_pkt_o[52] = 1'b0;
  assign data_mem_pkt_o[53] = 1'b0;
  assign data_mem_pkt_o[54] = 1'b0;
  assign data_mem_pkt_o[55] = 1'b0;
  assign data_mem_pkt_o[56] = 1'b0;
  assign data_mem_pkt_o[57] = 1'b0;
  assign data_mem_pkt_o[58] = 1'b0;
  assign data_mem_pkt_o[59] = 1'b0;
  assign data_mem_pkt_o[60] = 1'b0;
  assign data_mem_pkt_o[61] = 1'b0;
  assign data_mem_pkt_o[62] = 1'b0;
  assign data_mem_pkt_o[63] = 1'b0;
  assign data_mem_pkt_o[64] = 1'b0;
  assign data_mem_pkt_o[65] = 1'b0;
  assign data_mem_pkt_o[66] = 1'b0;
  assign data_mem_pkt_o[67] = 1'b0;
  assign data_mem_pkt_o[68] = 1'b0;
  assign data_mem_pkt_o[69] = 1'b0;
  assign data_mem_pkt_o[70] = 1'b0;
  assign data_mem_pkt_o[71] = 1'b0;
  assign data_mem_pkt_o[72] = 1'b0;
  assign data_mem_pkt_o[73] = 1'b0;
  assign data_mem_pkt_o[74] = 1'b0;
  assign data_mem_pkt_o[75] = 1'b0;
  assign data_mem_pkt_o[76] = 1'b0;
  assign data_mem_pkt_o[77] = 1'b0;
  assign data_mem_pkt_o[78] = 1'b0;
  assign data_mem_pkt_o[79] = 1'b0;
  assign data_mem_pkt_o[80] = 1'b0;
  assign data_mem_pkt_o[81] = 1'b0;
  assign data_mem_pkt_o[82] = 1'b0;
  assign data_mem_pkt_o[83] = 1'b0;
  assign data_mem_pkt_o[84] = 1'b0;
  assign data_mem_pkt_o[85] = 1'b0;
  assign data_mem_pkt_o[86] = 1'b0;
  assign data_mem_pkt_o[87] = 1'b0;
  assign data_mem_pkt_o[88] = 1'b0;
  assign data_mem_pkt_o[89] = 1'b0;
  assign data_mem_pkt_o[90] = 1'b0;
  assign data_mem_pkt_o[91] = 1'b0;
  assign data_mem_pkt_o[92] = 1'b0;
  assign data_mem_pkt_o[93] = 1'b0;
  assign data_mem_pkt_o[94] = 1'b0;
  assign data_mem_pkt_o[95] = 1'b0;
  assign data_mem_pkt_o[96] = 1'b0;
  assign data_mem_pkt_o[97] = 1'b0;
  assign data_mem_pkt_o[98] = 1'b0;
  assign data_mem_pkt_o[99] = 1'b0;
  assign data_mem_pkt_o[100] = 1'b0;
  assign data_mem_pkt_o[101] = 1'b0;
  assign data_mem_pkt_o[102] = 1'b0;
  assign data_mem_pkt_o[103] = 1'b0;
  assign data_mem_pkt_o[104] = 1'b0;
  assign data_mem_pkt_o[105] = 1'b0;
  assign data_mem_pkt_o[106] = 1'b0;
  assign data_mem_pkt_o[107] = 1'b0;
  assign data_mem_pkt_o[108] = 1'b0;
  assign data_mem_pkt_o[109] = 1'b0;
  assign data_mem_pkt_o[110] = 1'b0;
  assign data_mem_pkt_o[111] = 1'b0;
  assign data_mem_pkt_o[112] = 1'b0;
  assign data_mem_pkt_o[113] = 1'b0;
  assign data_mem_pkt_o[114] = 1'b0;
  assign data_mem_pkt_o[115] = 1'b0;
  assign data_mem_pkt_o[116] = 1'b0;
  assign data_mem_pkt_o[117] = 1'b0;
  assign data_mem_pkt_o[118] = 1'b0;
  assign data_mem_pkt_o[119] = 1'b0;
  assign data_mem_pkt_o[120] = 1'b0;
  assign data_mem_pkt_o[121] = 1'b0;
  assign data_mem_pkt_o[122] = 1'b0;
  assign data_mem_pkt_o[123] = 1'b0;
  assign data_mem_pkt_o[124] = 1'b0;
  assign data_mem_pkt_o[125] = 1'b0;
  assign data_mem_pkt_o[126] = 1'b0;
  assign data_mem_pkt_o[127] = 1'b0;
  assign data_mem_pkt_o[128] = 1'b0;
  assign data_mem_pkt_o[129] = 1'b0;
  assign data_mem_pkt_o[130] = 1'b0;
  assign data_mem_pkt_o[131] = 1'b0;
  assign data_mem_pkt_o[132] = 1'b0;
  assign data_mem_pkt_o[133] = 1'b0;
  assign data_mem_pkt_o[134] = 1'b0;
  assign data_mem_pkt_o[135] = 1'b0;
  assign data_mem_pkt_o[136] = 1'b0;
  assign data_mem_pkt_o[137] = 1'b0;
  assign data_mem_pkt_o[138] = 1'b0;
  assign data_mem_pkt_o[139] = 1'b0;
  assign data_mem_pkt_o[140] = 1'b0;
  assign data_mem_pkt_o[141] = 1'b0;
  assign data_mem_pkt_o[142] = 1'b0;
  assign data_mem_pkt_o[143] = 1'b0;
  assign data_mem_pkt_o[144] = 1'b0;
  assign data_mem_pkt_o[145] = 1'b0;
  assign data_mem_pkt_o[146] = 1'b0;
  assign data_mem_pkt_o[147] = 1'b0;
  assign data_mem_pkt_o[148] = 1'b0;
  assign data_mem_pkt_o[149] = 1'b0;
  assign data_mem_pkt_o[150] = 1'b0;
  assign data_mem_pkt_o[151] = 1'b0;
  assign data_mem_pkt_o[152] = 1'b0;
  assign data_mem_pkt_o[153] = 1'b0;
  assign data_mem_pkt_o[154] = 1'b0;
  assign data_mem_pkt_o[155] = 1'b0;
  assign data_mem_pkt_o[156] = 1'b0;
  assign data_mem_pkt_o[157] = 1'b0;
  assign data_mem_pkt_o[158] = 1'b0;
  assign data_mem_pkt_o[159] = 1'b0;
  assign data_mem_pkt_o[160] = 1'b0;
  assign data_mem_pkt_o[161] = 1'b0;
  assign data_mem_pkt_o[162] = 1'b0;
  assign data_mem_pkt_o[163] = 1'b0;
  assign data_mem_pkt_o[164] = 1'b0;
  assign data_mem_pkt_o[165] = 1'b0;
  assign data_mem_pkt_o[166] = 1'b0;
  assign data_mem_pkt_o[167] = 1'b0;
  assign data_mem_pkt_o[168] = 1'b0;
  assign data_mem_pkt_o[169] = 1'b0;
  assign data_mem_pkt_o[170] = 1'b0;
  assign data_mem_pkt_o[171] = 1'b0;
  assign data_mem_pkt_o[172] = 1'b0;
  assign data_mem_pkt_o[173] = 1'b0;
  assign data_mem_pkt_o[174] = 1'b0;
  assign data_mem_pkt_o[175] = 1'b0;
  assign data_mem_pkt_o[176] = 1'b0;
  assign data_mem_pkt_o[177] = 1'b0;
  assign data_mem_pkt_o[178] = 1'b0;
  assign data_mem_pkt_o[179] = 1'b0;
  assign data_mem_pkt_o[180] = 1'b0;
  assign data_mem_pkt_o[181] = 1'b0;
  assign data_mem_pkt_o[182] = 1'b0;
  assign data_mem_pkt_o[183] = 1'b0;
  assign data_mem_pkt_o[184] = 1'b0;
  assign data_mem_pkt_o[185] = 1'b0;
  assign data_mem_pkt_o[186] = 1'b0;
  assign data_mem_pkt_o[187] = 1'b0;
  assign data_mem_pkt_o[188] = 1'b0;
  assign data_mem_pkt_o[189] = 1'b0;
  assign data_mem_pkt_o[190] = 1'b0;
  assign data_mem_pkt_o[191] = 1'b0;
  assign data_mem_pkt_o[192] = 1'b0;
  assign data_mem_pkt_o[193] = 1'b0;
  assign data_mem_pkt_o[194] = 1'b0;
  assign data_mem_pkt_o[195] = 1'b0;
  assign data_mem_pkt_o[196] = 1'b0;
  assign data_mem_pkt_o[197] = 1'b0;
  assign data_mem_pkt_o[198] = 1'b0;
  assign data_mem_pkt_o[199] = 1'b0;
  assign data_mem_pkt_o[200] = 1'b0;
  assign data_mem_pkt_o[201] = 1'b0;
  assign data_mem_pkt_o[202] = 1'b0;
  assign data_mem_pkt_o[203] = 1'b0;
  assign data_mem_pkt_o[204] = 1'b0;
  assign data_mem_pkt_o[205] = 1'b0;
  assign data_mem_pkt_o[206] = 1'b0;
  assign data_mem_pkt_o[207] = 1'b0;
  assign data_mem_pkt_o[208] = 1'b0;
  assign data_mem_pkt_o[209] = 1'b0;
  assign data_mem_pkt_o[210] = 1'b0;
  assign data_mem_pkt_o[211] = 1'b0;
  assign data_mem_pkt_o[212] = 1'b0;
  assign data_mem_pkt_o[213] = 1'b0;
  assign data_mem_pkt_o[214] = 1'b0;
  assign data_mem_pkt_o[215] = 1'b0;
  assign data_mem_pkt_o[216] = 1'b0;
  assign data_mem_pkt_o[217] = 1'b0;
  assign data_mem_pkt_o[218] = 1'b0;
  assign data_mem_pkt_o[219] = 1'b0;
  assign data_mem_pkt_o[220] = 1'b0;
  assign data_mem_pkt_o[221] = 1'b0;
  assign data_mem_pkt_o[222] = 1'b0;
  assign data_mem_pkt_o[223] = 1'b0;
  assign data_mem_pkt_o[224] = 1'b0;
  assign data_mem_pkt_o[225] = 1'b0;
  assign data_mem_pkt_o[226] = 1'b0;
  assign data_mem_pkt_o[227] = 1'b0;
  assign data_mem_pkt_o[228] = 1'b0;
  assign data_mem_pkt_o[229] = 1'b0;
  assign data_mem_pkt_o[230] = 1'b0;
  assign data_mem_pkt_o[231] = 1'b0;
  assign data_mem_pkt_o[232] = 1'b0;
  assign data_mem_pkt_o[233] = 1'b0;
  assign data_mem_pkt_o[234] = 1'b0;
  assign data_mem_pkt_o[235] = 1'b0;
  assign data_mem_pkt_o[236] = 1'b0;
  assign data_mem_pkt_o[237] = 1'b0;
  assign data_mem_pkt_o[238] = 1'b0;
  assign data_mem_pkt_o[239] = 1'b0;
  assign data_mem_pkt_o[240] = 1'b0;
  assign data_mem_pkt_o[241] = 1'b0;
  assign data_mem_pkt_o[242] = 1'b0;
  assign data_mem_pkt_o[243] = 1'b0;
  assign data_mem_pkt_o[244] = 1'b0;
  assign data_mem_pkt_o[245] = 1'b0;
  assign data_mem_pkt_o[246] = 1'b0;
  assign data_mem_pkt_o[247] = 1'b0;
  assign data_mem_pkt_o[248] = 1'b0;
  assign data_mem_pkt_o[249] = 1'b0;
  assign data_mem_pkt_o[250] = 1'b0;
  assign data_mem_pkt_o[251] = 1'b0;
  assign data_mem_pkt_o[252] = 1'b0;
  assign data_mem_pkt_o[253] = 1'b0;
  assign data_mem_pkt_o[254] = 1'b0;
  assign data_mem_pkt_o[255] = 1'b0;
  assign data_mem_pkt_o[256] = 1'b0;
  assign data_mem_pkt_o[257] = 1'b0;
  assign data_mem_pkt_o[258] = 1'b0;
  assign data_mem_pkt_o[259] = 1'b0;
  assign data_mem_pkt_o[260] = 1'b0;
  assign data_mem_pkt_o[261] = 1'b0;
  assign data_mem_pkt_o[262] = 1'b0;
  assign data_mem_pkt_o[263] = 1'b0;
  assign data_mem_pkt_o[264] = 1'b0;
  assign data_mem_pkt_o[265] = 1'b0;
  assign data_mem_pkt_o[266] = 1'b0;
  assign data_mem_pkt_o[267] = 1'b0;
  assign data_mem_pkt_o[268] = 1'b0;
  assign data_mem_pkt_o[269] = 1'b0;
  assign data_mem_pkt_o[270] = 1'b0;
  assign data_mem_pkt_o[271] = 1'b0;
  assign data_mem_pkt_o[272] = 1'b0;
  assign data_mem_pkt_o[273] = 1'b0;
  assign data_mem_pkt_o[274] = 1'b0;
  assign data_mem_pkt_o[275] = 1'b0;
  assign data_mem_pkt_o[276] = 1'b0;
  assign data_mem_pkt_o[277] = 1'b0;
  assign data_mem_pkt_o[278] = 1'b0;
  assign data_mem_pkt_o[279] = 1'b0;
  assign data_mem_pkt_o[280] = 1'b0;
  assign data_mem_pkt_o[281] = 1'b0;
  assign data_mem_pkt_o[282] = 1'b0;
  assign data_mem_pkt_o[283] = 1'b0;
  assign data_mem_pkt_o[284] = 1'b0;
  assign data_mem_pkt_o[285] = 1'b0;
  assign data_mem_pkt_o[286] = 1'b0;
  assign data_mem_pkt_o[287] = 1'b0;
  assign data_mem_pkt_o[288] = 1'b0;
  assign data_mem_pkt_o[289] = 1'b0;
  assign data_mem_pkt_o[290] = 1'b0;
  assign data_mem_pkt_o[291] = 1'b0;
  assign data_mem_pkt_o[292] = 1'b0;
  assign data_mem_pkt_o[293] = 1'b0;
  assign data_mem_pkt_o[294] = 1'b0;
  assign data_mem_pkt_o[295] = 1'b0;
  assign data_mem_pkt_o[296] = 1'b0;
  assign data_mem_pkt_o[297] = 1'b0;
  assign data_mem_pkt_o[298] = 1'b0;
  assign data_mem_pkt_o[299] = 1'b0;
  assign data_mem_pkt_o[300] = 1'b0;
  assign data_mem_pkt_o[301] = 1'b0;
  assign data_mem_pkt_o[302] = 1'b0;
  assign data_mem_pkt_o[303] = 1'b0;
  assign data_mem_pkt_o[304] = 1'b0;
  assign data_mem_pkt_o[305] = 1'b0;
  assign data_mem_pkt_o[306] = 1'b0;
  assign data_mem_pkt_o[307] = 1'b0;
  assign data_mem_pkt_o[308] = 1'b0;
  assign data_mem_pkt_o[309] = 1'b0;
  assign data_mem_pkt_o[310] = 1'b0;
  assign data_mem_pkt_o[311] = 1'b0;
  assign data_mem_pkt_o[312] = 1'b0;
  assign data_mem_pkt_o[313] = 1'b0;
  assign data_mem_pkt_o[314] = 1'b0;
  assign data_mem_pkt_o[315] = 1'b0;
  assign data_mem_pkt_o[316] = 1'b0;
  assign data_mem_pkt_o[317] = 1'b0;
  assign data_mem_pkt_o[318] = 1'b0;
  assign data_mem_pkt_o[319] = 1'b0;
  assign data_mem_pkt_o[320] = 1'b0;
  assign data_mem_pkt_o[321] = 1'b0;
  assign data_mem_pkt_o[322] = 1'b0;
  assign data_mem_pkt_o[323] = 1'b0;
  assign data_mem_pkt_o[324] = 1'b0;
  assign data_mem_pkt_o[325] = 1'b0;
  assign data_mem_pkt_o[326] = 1'b0;
  assign data_mem_pkt_o[327] = 1'b0;
  assign data_mem_pkt_o[328] = 1'b0;
  assign data_mem_pkt_o[329] = 1'b0;
  assign data_mem_pkt_o[330] = 1'b0;
  assign data_mem_pkt_o[331] = 1'b0;
  assign data_mem_pkt_o[332] = 1'b0;
  assign data_mem_pkt_o[333] = 1'b0;
  assign data_mem_pkt_o[334] = 1'b0;
  assign data_mem_pkt_o[335] = 1'b0;
  assign data_mem_pkt_o[336] = 1'b0;
  assign data_mem_pkt_o[337] = 1'b0;
  assign data_mem_pkt_o[338] = 1'b0;
  assign data_mem_pkt_o[339] = 1'b0;
  assign data_mem_pkt_o[340] = 1'b0;
  assign data_mem_pkt_o[341] = 1'b0;
  assign data_mem_pkt_o[342] = 1'b0;
  assign data_mem_pkt_o[343] = 1'b0;
  assign data_mem_pkt_o[344] = 1'b0;
  assign data_mem_pkt_o[345] = 1'b0;
  assign data_mem_pkt_o[346] = 1'b0;
  assign data_mem_pkt_o[347] = 1'b0;
  assign data_mem_pkt_o[348] = 1'b0;
  assign data_mem_pkt_o[349] = 1'b0;
  assign data_mem_pkt_o[350] = 1'b0;
  assign data_mem_pkt_o[351] = 1'b0;
  assign data_mem_pkt_o[352] = 1'b0;
  assign data_mem_pkt_o[353] = 1'b0;
  assign data_mem_pkt_o[354] = 1'b0;
  assign data_mem_pkt_o[355] = 1'b0;
  assign data_mem_pkt_o[356] = 1'b0;
  assign data_mem_pkt_o[357] = 1'b0;
  assign data_mem_pkt_o[358] = 1'b0;
  assign data_mem_pkt_o[359] = 1'b0;
  assign data_mem_pkt_o[360] = 1'b0;
  assign data_mem_pkt_o[361] = 1'b0;
  assign data_mem_pkt_o[362] = 1'b0;
  assign data_mem_pkt_o[363] = 1'b0;
  assign data_mem_pkt_o[364] = 1'b0;
  assign data_mem_pkt_o[365] = 1'b0;
  assign data_mem_pkt_o[366] = 1'b0;
  assign data_mem_pkt_o[367] = 1'b0;
  assign data_mem_pkt_o[368] = 1'b0;
  assign data_mem_pkt_o[369] = 1'b0;
  assign data_mem_pkt_o[370] = 1'b0;
  assign data_mem_pkt_o[371] = 1'b0;
  assign data_mem_pkt_o[372] = 1'b0;
  assign data_mem_pkt_o[373] = 1'b0;
  assign data_mem_pkt_o[374] = 1'b0;
  assign data_mem_pkt_o[375] = 1'b0;
  assign data_mem_pkt_o[376] = 1'b0;
  assign data_mem_pkt_o[377] = 1'b0;
  assign data_mem_pkt_o[378] = 1'b0;
  assign data_mem_pkt_o[379] = 1'b0;
  assign data_mem_pkt_o[380] = 1'b0;
  assign data_mem_pkt_o[381] = 1'b0;
  assign data_mem_pkt_o[382] = 1'b0;
  assign data_mem_pkt_o[383] = 1'b0;
  assign data_mem_pkt_o[384] = 1'b0;
  assign data_mem_pkt_o[385] = 1'b0;
  assign data_mem_pkt_o[386] = 1'b0;
  assign data_mem_pkt_o[387] = 1'b0;
  assign data_mem_pkt_o[388] = 1'b0;
  assign data_mem_pkt_o[389] = 1'b0;
  assign data_mem_pkt_o[390] = 1'b0;
  assign data_mem_pkt_o[391] = 1'b0;
  assign data_mem_pkt_o[392] = 1'b0;
  assign data_mem_pkt_o[393] = 1'b0;
  assign data_mem_pkt_o[394] = 1'b0;
  assign data_mem_pkt_o[395] = 1'b0;
  assign data_mem_pkt_o[396] = 1'b0;
  assign data_mem_pkt_o[397] = 1'b0;
  assign data_mem_pkt_o[398] = 1'b0;
  assign data_mem_pkt_o[399] = 1'b0;
  assign data_mem_pkt_o[400] = 1'b0;
  assign data_mem_pkt_o[401] = 1'b0;
  assign data_mem_pkt_o[402] = 1'b0;
  assign data_mem_pkt_o[403] = 1'b0;
  assign data_mem_pkt_o[404] = 1'b0;
  assign data_mem_pkt_o[405] = 1'b0;
  assign data_mem_pkt_o[406] = 1'b0;
  assign data_mem_pkt_o[407] = 1'b0;
  assign data_mem_pkt_o[408] = 1'b0;
  assign data_mem_pkt_o[409] = 1'b0;
  assign data_mem_pkt_o[410] = 1'b0;
  assign data_mem_pkt_o[411] = 1'b0;
  assign data_mem_pkt_o[412] = 1'b0;
  assign data_mem_pkt_o[413] = 1'b0;
  assign data_mem_pkt_o[414] = 1'b0;
  assign data_mem_pkt_o[415] = 1'b0;
  assign data_mem_pkt_o[416] = 1'b0;
  assign data_mem_pkt_o[417] = 1'b0;
  assign data_mem_pkt_o[418] = 1'b0;
  assign data_mem_pkt_o[419] = 1'b0;
  assign data_mem_pkt_o[420] = 1'b0;
  assign data_mem_pkt_o[421] = 1'b0;
  assign data_mem_pkt_o[422] = 1'b0;
  assign data_mem_pkt_o[423] = 1'b0;
  assign data_mem_pkt_o[424] = 1'b0;
  assign data_mem_pkt_o[425] = 1'b0;
  assign data_mem_pkt_o[426] = 1'b0;
  assign data_mem_pkt_o[427] = 1'b0;
  assign data_mem_pkt_o[428] = 1'b0;
  assign data_mem_pkt_o[429] = 1'b0;
  assign data_mem_pkt_o[430] = 1'b0;
  assign data_mem_pkt_o[431] = 1'b0;
  assign data_mem_pkt_o[432] = 1'b0;
  assign data_mem_pkt_o[433] = 1'b0;
  assign data_mem_pkt_o[434] = 1'b0;
  assign data_mem_pkt_o[435] = 1'b0;
  assign data_mem_pkt_o[436] = 1'b0;
  assign data_mem_pkt_o[437] = 1'b0;
  assign data_mem_pkt_o[438] = 1'b0;
  assign data_mem_pkt_o[439] = 1'b0;
  assign data_mem_pkt_o[440] = 1'b0;
  assign data_mem_pkt_o[441] = 1'b0;
  assign data_mem_pkt_o[442] = 1'b0;
  assign data_mem_pkt_o[443] = 1'b0;
  assign data_mem_pkt_o[444] = 1'b0;
  assign data_mem_pkt_o[445] = 1'b0;
  assign data_mem_pkt_o[446] = 1'b0;
  assign data_mem_pkt_o[447] = 1'b0;
  assign data_mem_pkt_o[448] = 1'b0;
  assign data_mem_pkt_o[449] = 1'b0;
  assign data_mem_pkt_o[450] = 1'b0;
  assign data_mem_pkt_o[451] = 1'b0;
  assign data_mem_pkt_o[452] = 1'b0;
  assign data_mem_pkt_o[453] = 1'b0;
  assign data_mem_pkt_o[454] = 1'b0;
  assign data_mem_pkt_o[455] = 1'b0;
  assign data_mem_pkt_o[456] = 1'b0;
  assign data_mem_pkt_o[457] = 1'b0;
  assign data_mem_pkt_o[458] = 1'b0;
  assign data_mem_pkt_o[459] = 1'b0;
  assign data_mem_pkt_o[460] = 1'b0;
  assign data_mem_pkt_o[461] = 1'b0;
  assign data_mem_pkt_o[462] = 1'b0;
  assign data_mem_pkt_o[463] = 1'b0;
  assign data_mem_pkt_o[464] = 1'b0;
  assign data_mem_pkt_o[465] = 1'b0;
  assign data_mem_pkt_o[466] = 1'b0;
  assign data_mem_pkt_o[467] = 1'b0;
  assign data_mem_pkt_o[468] = 1'b0;
  assign data_mem_pkt_o[469] = 1'b0;
  assign data_mem_pkt_o[470] = 1'b0;
  assign data_mem_pkt_o[471] = 1'b0;
  assign data_mem_pkt_o[472] = 1'b0;
  assign data_mem_pkt_o[473] = 1'b0;
  assign data_mem_pkt_o[474] = 1'b0;
  assign data_mem_pkt_o[475] = 1'b0;
  assign data_mem_pkt_o[476] = 1'b0;
  assign data_mem_pkt_o[477] = 1'b0;
  assign data_mem_pkt_o[478] = 1'b0;
  assign data_mem_pkt_o[479] = 1'b0;
  assign data_mem_pkt_o[480] = 1'b0;
  assign data_mem_pkt_o[481] = 1'b0;
  assign data_mem_pkt_o[482] = 1'b0;
  assign data_mem_pkt_o[483] = 1'b0;
  assign data_mem_pkt_o[484] = 1'b0;
  assign data_mem_pkt_o[485] = 1'b0;
  assign data_mem_pkt_o[486] = 1'b0;
  assign data_mem_pkt_o[487] = 1'b0;
  assign data_mem_pkt_o[488] = 1'b0;
  assign data_mem_pkt_o[489] = 1'b0;
  assign data_mem_pkt_o[490] = 1'b0;
  assign data_mem_pkt_o[491] = 1'b0;
  assign data_mem_pkt_o[492] = 1'b0;
  assign data_mem_pkt_o[493] = 1'b0;
  assign data_mem_pkt_o[494] = 1'b0;
  assign data_mem_pkt_o[495] = 1'b0;
  assign data_mem_pkt_o[496] = 1'b0;
  assign data_mem_pkt_o[497] = 1'b0;
  assign data_mem_pkt_o[498] = 1'b0;
  assign data_mem_pkt_o[499] = 1'b0;
  assign data_mem_pkt_o[500] = 1'b0;
  assign data_mem_pkt_o[501] = 1'b0;
  assign data_mem_pkt_o[502] = 1'b0;
  assign data_mem_pkt_o[503] = 1'b0;
  assign data_mem_pkt_o[504] = 1'b0;
  assign data_mem_pkt_o[505] = 1'b0;
  assign data_mem_pkt_o[506] = 1'b0;
  assign data_mem_pkt_o[507] = 1'b0;
  assign data_mem_pkt_o[508] = 1'b0;
  assign data_mem_pkt_o[509] = 1'b0;
  assign data_mem_pkt_o[510] = 1'b0;
  assign data_mem_pkt_o[511] = 1'b0;
  assign data_mem_pkt_o[512] = 1'b0;
  assign data_mem_pkt_o[513] = 1'b0;
  assign lce_data_cmd_o[3] = 1'b0;
  assign lce_data_cmd_o[4] = 1'b0;
  assign lce_resp_o[23] = 1'b0;
  assign lce_data_resp_o[23] = lce_id_i[0];
  assign lce_resp_o[24] = lce_id_i[0];
  assign N31 = N28 & N29;
  assign N32 = N31 & N30;
  assign N33 = state_r[2] | state_r[1];
  assign N34 = N33 | N30;
  assign N36 = state_r[2] | N29;
  assign N37 = N36 | state_r[0];
  assign N39 = state_r[2] | N29;
  assign N40 = N39 | N30;
  assign N42 = N28 | state_r[1];
  assign N43 = N42 | state_r[0];
  assign N45 = N28 | state_r[1];
  assign N46 = N45 | N30;
  assign N48 = state_r[2] & state_r[1];
  assign N49 = N86 & N75;
  assign N50 = lce_cmd_i[33] | lce_cmd_i[32];
  assign N51 = N50 | N75;
  assign N68 = N70 | lce_cmd_i[31];
  assign N70 = lce_cmd_i[33] | N80;
  assign N71 = N70 | N75;
  assign N73 = N76 | lce_cmd_i[31];
  assign N76 = N79 | lce_cmd_i[32];
  assign N77 = N76 | N75;
  assign N81 = N79 | N80;
  assign N82 = N81 | lce_cmd_i[31];
  assign N84 = lce_cmd_i[33] & lce_cmd_i[32];
  assign N85 = N84 & lce_cmd_i[31];
  assign N86 = N79 & N80;
  assign N699 = (N691)? dirty_i[0] :
                (N693)? dirty_i[1] :
                (N695)? dirty_i[2] :
                (N697)? dirty_i[3] :
                (N692)? dirty_i[4] :
                (N694)? dirty_i[5] :
                (N696)? dirty_i[6] :
                (N698)? dirty_i[7] : 1'b0;
  assign N1605 = state_r[1] | state_r[2];
  assign lce_sync_done_o = state_r[0] | N1605;
  assign N1607 = ~sync_ack_count_r[0];
  assign N55 = sync_ack_count_r[0] ^ 1'b1;
  assign N58 = (N0)? lce_cmd_i[34] :
               (N1)? 1'b0 :
               (N2)? 1'b0 : 1'b0;
  assign N0 = N49;
  assign N1 = N52;
  assign N2 = N53;
  assign N59 = (N0)? lce_cmd_v_i :
               (N1)? 1'b0 :
               (N2)? 1'b0 : 1'b0;
  assign N60 = (N0)? lce_resp_yumi_i :
               (N1)? N57 :
               (N2)? 1'b0 : 1'b0;
  assign { N66, N65, N64, N63, N62, N61 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                            (N1)? lce_cmd_i[20:15] :
                                            (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N67 = (N0)? 1'b0 :
               (N1)? lce_cmd_v_i :
               (N2)? 1'b0 : 1'b0;
  assign N90 = (N3)? 1'b0 :
               (N4)? lce_cmd_v_i : 1'b0;
  assign N3 = invalidated_tag_r;
  assign N4 = N89;
  assign N93 = (N5)? 1'b0 :
               (N1238)? 1'b1 :
               (N92)? tag_mem_pkt_yumi_i : 1'b0;
  assign N5 = lce_resp_yumi_i;
  assign { N104, N103, N102, N101, N100, N99, N98, N97, N96, N95 } = (N6)? { lce_cmd_i[20:15], lce_cmd_i[8:6], 1'b1 } :
                                                                     (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                     (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                     (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                     (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                     (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N6 = N69;
  assign N7 = N72;
  assign N8 = N74;
  assign N9 = N78;
  assign N10 = N83;
  assign N11 = N87;
  assign N105 = (N6)? lce_cmd_v_i :
                (N7)? 1'b0 :
                (N8)? 1'b0 :
                (N9)? 1'b0 :
                (N10)? 1'b0 :
                (N11)? 1'b0 : 1'b0;
  assign { N107, N106 } = (N6)? { data_mem_pkt_yumi_i, N88 } :
                          (N7)? { stat_mem_pkt_yumi_i, 1'b1 } : 1'b0;
  assign { N117, N116, N115, N114, N113, N112, N111, N110, N109, N108 } = (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                          (N7)? { lce_cmd_i[20:15], lce_cmd_i[8:6], 1'b1 } :
                                                                          (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                          (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                          (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                          (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N118 = (N6)? 1'b0 :
                (N7)? lce_cmd_v_i :
                (N8)? 1'b0 :
                (N9)? 1'b0 :
                (N10)? 1'b0 :
                (N11)? 1'b0 : 1'b0;
  assign { N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119 } = (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                  (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                  (N8)? { lce_cmd_i[20:15], lce_cmd_i[8:4], lce_cmd_i[30:21], 1'b1 } :
                                                                                                                                                  (N9)? { lce_cmd_i[20:15], lce_cmd_i[8:4], lce_cmd_i[30:21], 1'b1 } :
                                                                                                                                                  (N10)? { lce_cmd_i[20:15], lce_cmd_i[8:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                  (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N141 = (N6)? 1'b0 :
                (N7)? 1'b0 :
                (N8)? lce_cmd_v_i :
                (N9)? lce_cmd_v_i :
                (N10)? N90 :
                (N11)? 1'b0 : 1'b0;
  assign N142 = (N6)? 1'b0 :
                (N7)? 1'b0 :
                (N8)? tag_mem_pkt_yumi_i :
                (N9)? tag_mem_pkt_yumi_i :
                (N10)? lce_resp_yumi_i :
                (N11)? 1'b0 : 1'b0;
  assign N143 = (N6)? 1'b0 :
                (N7)? 1'b0 :
                (N8)? tag_mem_pkt_yumi_i :
                (N9)? 1'b0 :
                (N10)? 1'b0 :
                (N11)? 1'b0 : 1'b0;
  assign N144 = (N6)? 1'b0 :
                (N7)? 1'b0 :
                (N8)? 1'b0 :
                (N9)? tag_mem_pkt_yumi_i :
                (N10)? 1'b0 :
                (N11)? 1'b0 : 1'b0;
  assign { N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145 } = (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                              (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                              (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                              (N10)? { lce_cmd_i[34:34], 1'b1, lce_cmd_i[30:9] } :
                                                                                                                                                              (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N169 = (N6)? 1'b0 :
                (N7)? 1'b0 :
                (N8)? 1'b0 :
                (N9)? 1'b0 :
                (N10)? N94 :
                (N11)? 1'b0 : 1'b0;
  assign { N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172 } = (N12)? data_buf_r :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N13)? data_mem_data_i : 1'b0;
  assign N12 = tr_data_buffered_r;
  assign N13 = N171;
  assign N700 = ~N699;
  assign N711 = (N14)? 1'b0 :
                (N1242)? 1'b1 :
                (N710)? wb_data_read_r : 1'b0;
  assign N14 = lce_data_resp_done;
  assign N714 = (N14)? 1'b0 :
                (N1243)? 1'b1 :
                (N713)? data_mem_pkt_yumi_i : 1'b0;
  assign N717 = (N15)? 1'b0 :
                (N16)? N716 : 1'b0;
  assign N15 = wb_dirty_cleared_r;
  assign N16 = N715;
  assign N720 = (N14)? 1'b0 :
                (N1244)? 1'b1 :
                (N719)? stat_mem_pkt_yumi_i : 1'b0;
  assign { N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722 } = (N17)? data_buf_r :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N18)? data_mem_data_i : 1'b0;
  assign N17 = wb_data_buffered_r;
  assign N18 = N721;
  assign stat_mem_pkt_o[0] = (N19)? N108 :
                             (N1236)? 1'b0 : 1'b0;
  assign N19 = N35;
  assign stat_mem_pkt_o[10:2] = (N20)? { N66, N65, N64, N63, N62, N61, 1'b0, 1'b0, 1'b0 } :
                                (N19)? { N117, N116, N115, N114, N113, N112, N111, N110, N109 } :
                                (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                (N23)? { lce_cmd_i[20:15], lce_cmd_i[8:6] } :
                                (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N20 = N32;
  assign N21 = N38;
  assign N22 = N41;
  assign N23 = stat_mem_pkt_o[1];
  assign N24 = N47;
  assign N25 = N48;
  assign stat_mem_pkt_v_o = (N20)? N67 :
                            (N19)? N118 :
                            (N21)? 1'b0 :
                            (N22)? 1'b0 :
                            (N23)? N717 :
                            (N24)? 1'b0 :
                            (N25)? 1'b0 : 1'b0;
  assign { lce_resp_o[25:25], lce_resp_o[22:0] } = (N20)? { N58, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                   (N19)? { N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145 } :
                                                   (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                   (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                   (N23)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                   (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                   (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_resp_v_o = (N20)? N59 :
                        (N19)? N169 :
                        (N21)? 1'b0 :
                        (N22)? 1'b0 :
                        (N23)? 1'b0 :
                        (N24)? 1'b0 :
                        (N25)? 1'b0 : 1'b0;
  assign lce_cmd_yumi_o = (N20)? N60 :
                          (N19)? N142 :
                          (N21)? lce_tr_done :
                          (N22)? 1'b0 :
                          (N23)? lce_data_resp_done :
                          (N24)? lce_data_resp_done :
                          (N25)? 1'b0 : 1'b0;
  assign state_n = (N20)? { 1'b0, 1'b0, N56 } :
                   (N19)? { 1'b0, N107, N106 } :
                   (N21)? { 1'b0, N170, lce_tr_done } :
                   (N22)? { 1'b1, 1'b0, N700 } :
                   (N23)? { N1235, 1'b0, lce_data_resp_done } :
                   (N24)? { N1235, 1'b0, 1'b1 } :
                   (N25)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_mem_pkt_o = (N20)? { N66, N65, N64, N63, N62, N61, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                         (N19)? { N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N83 } :
                         (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                         (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                         (N23)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                         (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                         (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_mem_pkt_v_o = (N20)? N67 :
                           (N19)? N141 :
                           (N21)? 1'b0 :
                           (N22)? 1'b0 :
                           (N23)? 1'b0 :
                           (N24)? 1'b0 :
                           (N25)? 1'b0 : 1'b0;
  assign { data_mem_pkt_o[522:514], data_mem_pkt_o[0:0] } = (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                            (N19)? { N104, N103, N102, N101, N100, N99, N98, N97, N96, N95 } :
                                                            (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                            (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                            (N23)? { lce_cmd_i[20:15], lce_cmd_i[8:6], 1'b1 } :
                                                            (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                            (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign data_mem_pkt_v_o = (N20)? 1'b0 :
                            (N19)? N105 :
                            (N21)? 1'b0 :
                            (N22)? 1'b0 :
                            (N23)? N701 :
                            (N24)? 1'b0 :
                            (N25)? 1'b0 : 1'b0;
  assign set_tag_received_o = (N20)? 1'b0 :
                              (N19)? N143 :
                              (N21)? 1'b0 :
                              (N22)? 1'b0 :
                              (N23)? 1'b0 :
                              (N24)? 1'b0 :
                              (N25)? 1'b0 : 1'b0;
  assign set_tag_wakeup_received_o = (N20)? 1'b0 :
                                     (N19)? N144 :
                                     (N21)? 1'b0 :
                                     (N22)? 1'b0 :
                                     (N23)? 1'b0 :
                                     (N24)? 1'b0 :
                                     (N25)? 1'b0 : 1'b0;
  assign { lce_data_cmd_o[517:5], lce_data_cmd_o[2:0] } = (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                          (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                          (N21)? { N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, lce_cmd_i[3:0] } :
                                                          (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                          (N23)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                          (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                          (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_data_cmd_v_o = (N20)? 1'b0 :
                            (N19)? 1'b0 :
                            (N21)? 1'b1 :
                            (N22)? 1'b0 :
                            (N23)? 1'b0 :
                            (N24)? 1'b0 :
                            (N25)? 1'b0 : 1'b0;
  assign { lce_data_resp_o[536:24], lce_data_resp_o[22:0] } = (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                              (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                              (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                              (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                              (N23)? { N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, lce_cmd_i[34:34], 1'b0, lce_cmd_i[30:9] } :
                                                              (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_cmd_i[34:34], 1'b1, lce_cmd_i[30:9] } :
                                                              (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign lce_data_resp_v_o = (N20)? 1'b0 :
                             (N19)? 1'b0 :
                             (N21)? 1'b0 :
                             (N22)? 1'b0 :
                             (N23)? N1234 :
                             (N24)? 1'b1 :
                             (N25)? 1'b0 : 1'b0;
  assign { N1248, N1247, N1246 } = (N26)? { 1'b0, 1'b0, 1'b0 } :
                                   (N27)? state_n : 1'b0;
  assign N26 = reset_i;
  assign N27 = N1245;
  assign N1249 = (N26)? 1'b0 :
                 (N27)? N55 : 1'b0;
  assign N1250 = (N26)? 1'b0 :
                 (N27)? N170 : 1'b0;
  assign N1251 = (N26)? 1'b0 :
                 (N27)? N711 : 1'b0;
  assign N1252 = (N26)? 1'b0 :
                 (N27)? N714 : 1'b0;
  assign N1253 = (N26)? 1'b0 :
                 (N27)? N720 : 1'b0;
  assign N1254 = (N26)? 1'b0 :
                 (N27)? N93 : 1'b0;
  assign lce_tr_done = lce_data_cmd_v_o & lce_data_cmd_ready_i;
  assign lce_data_resp_done = lce_data_resp_ready_i & lce_data_resp_v_o;
  assign N28 = ~state_r[2];
  assign N29 = ~state_r[1];
  assign N30 = ~state_r[0];
  assign N35 = ~N34;
  assign N38 = ~N37;
  assign N41 = ~N40;
  assign N44 = ~N43;
  assign N47 = ~N46;
  assign stat_mem_pkt_o[1] = N44;
  assign N52 = ~N51;
  assign N53 = lce_cmd_i[33] | lce_cmd_i[32];
  assign N54 = ~lce_resp_yumi_i;
  assign N56 = N1607 & lce_resp_yumi_i;
  assign N57 = tag_mem_pkt_yumi_i & stat_mem_pkt_yumi_i;
  assign N69 = ~N68;
  assign N72 = ~N71;
  assign N74 = ~N73;
  assign N75 = ~lce_cmd_i[31];
  assign N78 = ~N77;
  assign N79 = ~lce_cmd_i[33];
  assign N80 = ~lce_cmd_i[32];
  assign N83 = ~N82;
  assign N87 = N85 | N86;
  assign N88 = ~data_mem_pkt_yumi_i;
  assign N89 = ~invalidated_tag_r;
  assign N91 = invalidated_tag_r | lce_resp_yumi_i;
  assign N92 = ~N91;
  assign N94 = invalidated_tag_r | tag_mem_pkt_yumi_i;
  assign N170 = ~lce_tr_done;
  assign N171 = ~tr_data_buffered_r;
  assign N684 = ~lce_cmd_i[6];
  assign N685 = ~lce_cmd_i[7];
  assign N686 = N684 & N685;
  assign N687 = N684 & lce_cmd_i[7];
  assign N688 = lce_cmd_i[6] & N685;
  assign N689 = lce_cmd_i[6] & lce_cmd_i[7];
  assign N690 = ~lce_cmd_i[8];
  assign N691 = N686 & N690;
  assign N692 = N686 & lce_cmd_i[8];
  assign N693 = N688 & N690;
  assign N694 = N688 & lce_cmd_i[8];
  assign N695 = N687 & N690;
  assign N696 = N687 & lce_cmd_i[8];
  assign N697 = N689 & N690;
  assign N698 = N689 & lce_cmd_i[8];
  assign N701 = ~wb_data_read_r;
  assign N702 = ~N1240;
  assign N703 = N702;
  assign N704 = N702;
  assign N705 = N702;
  assign N706 = N702;
  assign N707 = N702;
  assign N708 = N702;
  assign N709 = wb_data_buffered_r | lce_data_resp_done;
  assign N710 = ~N709;
  assign N712 = wb_data_read_r | lce_data_resp_done;
  assign N713 = ~N712;
  assign N715 = ~wb_dirty_cleared_r;
  assign N716 = wb_data_read_r | data_mem_pkt_yumi_i;
  assign N718 = wb_dirty_cleared_r | lce_data_resp_done;
  assign N719 = ~N718;
  assign N721 = ~wb_data_buffered_r;
  assign N1234 = wb_data_read_r & N1608;
  assign N1608 = wb_dirty_cleared_r | stat_mem_pkt_yumi_i;
  assign N1235 = ~lce_data_resp_done;
  assign N1236 = N34;
  assign N1237 = ~lce_resp_yumi_i;
  assign N1238 = invalidated_tag_r & N1237;
  assign N1239 = ~wb_data_buffered_r;
  assign N1240 = wb_data_read_r & N1239;
  assign N1241 = ~lce_data_resp_done;
  assign N1242 = wb_data_buffered_r & N1241;
  assign N1243 = wb_data_read_r & N1241;
  assign N1244 = wb_dirty_cleared_r & N1241;
  assign N1245 = ~reset_i;
  assign N1255 = N32 & N1245;
  assign N1256 = N35 & N1245;
  assign N1257 = N1255 | N1256;
  assign N1258 = N38 & N1245;
  assign N1259 = tr_data_buffered_r & N1258;
  assign N1260 = N1257 | N1259;
  assign N1261 = N41 & N1245;
  assign N1262 = N1260 | N1261;
  assign N1263 = stat_mem_pkt_o[1] & N1245;
  assign N1264 = N703 & N1263;
  assign N1265 = N1262 | N1264;
  assign N1266 = N47 & N1245;
  assign N1267 = N1265 | N1266;
  assign N1268 = N48 & N1245;
  assign N1269 = N1267 | N1268;
  assign N1270 = ~N1269;
  assign N1271 = N1245 & N1270;
  assign N1272 = N32 & N1245;
  assign N1273 = N35 & N1245;
  assign N1274 = N1272 | N1273;
  assign N1275 = N38 & N1245;
  assign N1276 = tr_data_buffered_r & N1275;
  assign N1277 = N1274 | N1276;
  assign N1278 = N41 & N1245;
  assign N1279 = N1277 | N1278;
  assign N1280 = stat_mem_pkt_o[1] & N1245;
  assign N1281 = N703 & N1280;
  assign N1282 = N1279 | N1281;
  assign N1283 = N47 & N1245;
  assign N1284 = N1282 | N1283;
  assign N1285 = N48 & N1245;
  assign N1286 = N1284 | N1285;
  assign N1287 = ~N1286;
  assign N1288 = N1245 & N1287;
  assign N1289 = N32 & N1245;
  assign N1290 = N35 & N1245;
  assign N1291 = N1289 | N1290;
  assign N1292 = N38 & N1245;
  assign N1293 = tr_data_buffered_r & N1292;
  assign N1294 = N1291 | N1293;
  assign N1295 = N41 & N1245;
  assign N1296 = N1294 | N1295;
  assign N1297 = stat_mem_pkt_o[1] & N1245;
  assign N1298 = N703 & N1297;
  assign N1299 = N1296 | N1298;
  assign N1300 = N47 & N1245;
  assign N1301 = N1299 | N1300;
  assign N1302 = N48 & N1245;
  assign N1303 = N1301 | N1302;
  assign N1304 = ~N1303;
  assign N1305 = N1245 & N1304;
  assign N1306 = N32 & N1245;
  assign N1307 = N35 & N1245;
  assign N1308 = N1306 | N1307;
  assign N1309 = N38 & N1245;
  assign N1310 = tr_data_buffered_r & N1309;
  assign N1311 = N1308 | N1310;
  assign N1312 = N41 & N1245;
  assign N1313 = N1311 | N1312;
  assign N1314 = stat_mem_pkt_o[1] & N1245;
  assign N1315 = N703 & N1314;
  assign N1316 = N1313 | N1315;
  assign N1317 = N47 & N1245;
  assign N1318 = N1316 | N1317;
  assign N1319 = N48 & N1245;
  assign N1320 = N1318 | N1319;
  assign N1321 = ~N1320;
  assign N1322 = N1245 & N1321;
  assign N1323 = N32 & N1245;
  assign N1324 = N35 & N1245;
  assign N1325 = N1323 | N1324;
  assign N1326 = N38 & N1245;
  assign N1327 = tr_data_buffered_r & N1326;
  assign N1328 = N1325 | N1327;
  assign N1329 = N41 & N1245;
  assign N1330 = N1328 | N1329;
  assign N1331 = stat_mem_pkt_o[1] & N1245;
  assign N1332 = N703 & N1331;
  assign N1333 = N1330 | N1332;
  assign N1334 = N47 & N1245;
  assign N1335 = N1333 | N1334;
  assign N1336 = N48 & N1245;
  assign N1337 = N1335 | N1336;
  assign N1338 = ~N1337;
  assign N1339 = N1245 & N1338;
  assign N1340 = N32 & N1245;
  assign N1341 = N35 & N1245;
  assign N1342 = N1340 | N1341;
  assign N1343 = N38 & N1245;
  assign N1344 = tr_data_buffered_r & N1343;
  assign N1345 = N1342 | N1344;
  assign N1346 = N41 & N1245;
  assign N1347 = N1345 | N1346;
  assign N1348 = stat_mem_pkt_o[1] & N1245;
  assign N1349 = N703 & N1348;
  assign N1350 = N1347 | N1349;
  assign N1351 = N47 & N1245;
  assign N1352 = N1350 | N1351;
  assign N1353 = N48 & N1245;
  assign N1354 = N1352 | N1353;
  assign N1355 = ~N1354;
  assign N1356 = N1245 & N1355;
  assign N1357 = N1347 | N1332;
  assign N1358 = N1357 | N1351;
  assign N1359 = N1358 | N1353;
  assign N1360 = ~N1359;
  assign N1361 = N1245 & N1360;
  assign N1362 = N1342 | N1327;
  assign N1363 = N1362 | N1346;
  assign N1364 = N1363 | N1332;
  assign N1365 = N1364 | N1351;
  assign N1366 = N1365 | N1353;
  assign N1367 = ~N1366;
  assign N1368 = N1245 & N1367;
  assign N1369 = N1362 | N1329;
  assign N1370 = N1369 | N1332;
  assign N1371 = N1370 | N1334;
  assign N1372 = N1371 | N1336;
  assign N1373 = ~N1372;
  assign N1374 = N1245 & N1373;
  assign N1375 = N1323 | N1341;
  assign N1376 = N1375 | N1327;
  assign N1377 = N1376 | N1329;
  assign N1378 = N1377 | N1332;
  assign N1379 = N1378 | N1334;
  assign N1380 = N1379 | N1336;
  assign N1381 = ~N1380;
  assign N1382 = N1245 & N1381;
  assign N1383 = N704 & N1331;
  assign N1384 = N1330 | N1383;
  assign N1385 = N1384 | N1334;
  assign N1386 = N1385 | N1336;
  assign N1387 = ~N1386;
  assign N1388 = N1245 & N1387;
  assign N1389 = N704 & N1314;
  assign N1390 = N1330 | N1389;
  assign N1391 = N1390 | N1334;
  assign N1392 = N1391 | N1336;
  assign N1393 = ~N1392;
  assign N1394 = N1245 & N1393;
  assign N1395 = N1325 | N1310;
  assign N1396 = N1395 | N1329;
  assign N1397 = N1396 | N1389;
  assign N1398 = N1397 | N1334;
  assign N1399 = N1398 | N1336;
  assign N1400 = ~N1399;
  assign N1401 = N1245 & N1400;
  assign N1402 = N1395 | N1312;
  assign N1403 = N1402 | N1389;
  assign N1404 = N1403 | N1317;
  assign N1405 = N1404 | N1319;
  assign N1406 = ~N1405;
  assign N1407 = N1245 & N1406;
  assign N1408 = N1306 | N1324;
  assign N1409 = N1408 | N1310;
  assign N1410 = N1409 | N1312;
  assign N1411 = N1410 | N1389;
  assign N1412 = N1411 | N1317;
  assign N1413 = N1412 | N1319;
  assign N1414 = ~N1413;
  assign N1415 = N1245 & N1414;
  assign N1416 = N1313 | N1389;
  assign N1417 = N1416 | N1317;
  assign N1418 = N1417 | N1319;
  assign N1419 = ~N1418;
  assign N1420 = N1245 & N1419;
  assign N1421 = N705 & N1314;
  assign N1422 = N1313 | N1421;
  assign N1423 = N1422 | N1317;
  assign N1424 = N1423 | N1319;
  assign N1425 = ~N1424;
  assign N1426 = N1245 & N1425;
  assign N1427 = N705 & N1297;
  assign N1428 = N1313 | N1427;
  assign N1429 = N1428 | N1317;
  assign N1430 = N1429 | N1319;
  assign N1431 = ~N1430;
  assign N1432 = N1245 & N1431;
  assign N1433 = N1308 | N1293;
  assign N1434 = N1433 | N1312;
  assign N1435 = N1434 | N1427;
  assign N1436 = N1435 | N1317;
  assign N1437 = N1436 | N1319;
  assign N1438 = ~N1437;
  assign N1439 = N1245 & N1438;
  assign N1440 = N1433 | N1295;
  assign N1441 = N1440 | N1427;
  assign N1442 = N1441 | N1300;
  assign N1443 = N1442 | N1302;
  assign N1444 = ~N1443;
  assign N1445 = N1245 & N1444;
  assign N1446 = N1289 | N1307;
  assign N1447 = N1446 | N1293;
  assign N1448 = N1447 | N1295;
  assign N1449 = N1448 | N1427;
  assign N1450 = N1449 | N1300;
  assign N1451 = N1450 | N1302;
  assign N1452 = ~N1451;
  assign N1453 = N1245 & N1452;
  assign N1454 = N1296 | N1427;
  assign N1455 = N1454 | N1300;
  assign N1456 = N1455 | N1302;
  assign N1457 = ~N1456;
  assign N1458 = N1245 & N1457;
  assign N1459 = N706 & N1297;
  assign N1460 = N1296 | N1459;
  assign N1461 = N1460 | N1300;
  assign N1462 = N1461 | N1302;
  assign N1463 = ~N1462;
  assign N1464 = N1245 & N1463;
  assign N1465 = N706 & N1280;
  assign N1466 = N1296 | N1465;
  assign N1467 = N1466 | N1300;
  assign N1468 = N1467 | N1302;
  assign N1469 = ~N1468;
  assign N1470 = N1245 & N1469;
  assign N1471 = N1291 | N1276;
  assign N1472 = N1471 | N1295;
  assign N1473 = N1472 | N1465;
  assign N1474 = N1473 | N1300;
  assign N1475 = N1474 | N1302;
  assign N1476 = ~N1475;
  assign N1477 = N1245 & N1476;
  assign N1478 = N1471 | N1278;
  assign N1479 = N1478 | N1465;
  assign N1480 = N1479 | N1283;
  assign N1481 = N1480 | N1285;
  assign N1482 = ~N1481;
  assign N1483 = N1245 & N1482;
  assign N1484 = N1272 | N1290;
  assign N1485 = N1484 | N1276;
  assign N1486 = N1485 | N1278;
  assign N1487 = N1486 | N1465;
  assign N1488 = N1487 | N1283;
  assign N1489 = N1488 | N1285;
  assign N1490 = ~N1489;
  assign N1491 = N1245 & N1490;
  assign N1492 = N1279 | N1465;
  assign N1493 = N1492 | N1283;
  assign N1494 = N1493 | N1285;
  assign N1495 = ~N1494;
  assign N1496 = N1245 & N1495;
  assign N1497 = N707 & N1280;
  assign N1498 = N1279 | N1497;
  assign N1499 = N1498 | N1283;
  assign N1500 = N1499 | N1285;
  assign N1501 = ~N1500;
  assign N1502 = N1245 & N1501;
  assign N1503 = N707 & N1263;
  assign N1504 = N1279 | N1503;
  assign N1505 = N1504 | N1283;
  assign N1506 = N1505 | N1285;
  assign N1507 = ~N1506;
  assign N1508 = N1245 & N1507;
  assign N1509 = N1274 | N1259;
  assign N1510 = N1509 | N1278;
  assign N1511 = N1510 | N1503;
  assign N1512 = N1511 | N1283;
  assign N1513 = N1512 | N1285;
  assign N1514 = ~N1513;
  assign N1515 = N1245 & N1514;
  assign N1516 = N1509 | N1261;
  assign N1517 = N1516 | N1503;
  assign N1518 = N1517 | N1266;
  assign N1519 = N1518 | N1268;
  assign N1520 = ~N1519;
  assign N1521 = N1245 & N1520;
  assign N1522 = N1255 | N1273;
  assign N1523 = N1522 | N1259;
  assign N1524 = N1523 | N1261;
  assign N1525 = N1524 | N1503;
  assign N1526 = N1525 | N1266;
  assign N1527 = N1526 | N1268;
  assign N1528 = ~N1527;
  assign N1529 = N1245 & N1528;
  assign N1530 = N1262 | N1503;
  assign N1531 = N1530 | N1266;
  assign N1532 = N1531 | N1268;
  assign N1533 = ~N1532;
  assign N1534 = N1245 & N1533;
  assign N1535 = N708 & N1263;
  assign N1536 = N1262 | N1535;
  assign N1537 = N1536 | N1266;
  assign N1538 = N1537 | N1268;
  assign N1539 = ~N1538;
  assign N1540 = N1245 & N1539;
  assign N1541 = N706 & N1263;
  assign N1542 = N1262 | N1541;
  assign N1543 = N1542 | N1266;
  assign N1544 = N1543 | N1268;
  assign N1545 = ~N1544;
  assign N1546 = N1245 & N1545;
  assign N1547 = N705 & N1263;
  assign N1548 = N1262 | N1547;
  assign N1549 = N1548 | N1266;
  assign N1550 = N1549 | N1268;
  assign N1551 = ~N1550;
  assign N1552 = N1245 & N1551;
  assign N1553 = N704 & N1263;
  assign N1554 = N1262 | N1553;
  assign N1555 = N1554 | N1266;
  assign N1556 = N1555 | N1268;
  assign N1557 = ~N1556;
  assign N1558 = N1245 & N1557;
  assign N1559 = N52 & N1255;
  assign N1560 = N53 & N1255;
  assign N1561 = N1559 | N1560;
  assign N1562 = N74 & N1256;
  assign N1563 = N1561 | N1562;
  assign N1564 = N78 & N1256;
  assign N1565 = N1563 | N1564;
  assign N1566 = N83 & N1256;
  assign N1567 = N1565 | N1566;
  assign N1568 = N87 & N1256;
  assign N1569 = N1567 | N1568;
  assign N1570 = ~N1569;
  assign N1571 = N49 & N1255;
  assign N1572 = N54 & N1571;
  assign N1573 = N1572 | N1559;
  assign N1574 = N1573 | N1560;
  assign N1575 = N1574 | N1256;
  assign N1576 = N1575 | N1258;
  assign N1577 = N1576 | N1261;
  assign N1578 = N1577 | N1263;
  assign N1579 = N1578 | N1266;
  assign N1580 = N1579 | N1268;
  assign N1581 = ~N1580;
  assign N1582 = N1257 | N1261;
  assign N1583 = N1582 | N1263;
  assign N1584 = N1583 | N1266;
  assign N1585 = N1584 | N1268;
  assign N1586 = ~N1585;
  assign N1587 = N1257 | N1258;
  assign N1588 = N1587 | N1261;
  assign N1589 = N1588 | N1266;
  assign N1590 = N1589 | N1268;
  assign N1591 = ~N1590;
  assign N1592 = N69 & N1256;
  assign N1593 = N1255 | N1592;
  assign N1594 = N72 & N1256;
  assign N1595 = N1593 | N1594;
  assign N1596 = N1595 | N1562;
  assign N1597 = N1596 | N1564;
  assign N1598 = N1597 | N1568;
  assign N1599 = N1598 | N1258;
  assign N1600 = N1599 | N1261;
  assign N1601 = N1600 | N1263;
  assign N1602 = N1601 | N1266;
  assign N1603 = N1602 | N1268;
  assign N1604 = ~N1603;

  always @(posedge clk_i) begin
    if(N1271) begin
      { data_buf_r[511:511], data_buf_r[0:0] } <= { data_mem_data_i[511:511], data_mem_data_i[0:0] };
    end
    if(N1288) begin
      { data_buf_r[510:510] } <= { data_mem_data_i[510:510] };
    end
    if(N1305) begin
      { data_buf_r[509:509] } <= { data_mem_data_i[509:509] };
    end
    if(N1322) begin
      { data_buf_r[508:508] } <= { data_mem_data_i[508:508] };
    end
    if(N1339) begin
      { data_buf_r[507:507], data_buf_r[472:413] } <= { data_mem_data_i[507:507], data_mem_data_i[472:413] };
    end
    if(N1356) begin
      { data_buf_r[506:492] } <= { data_mem_data_i[506:492] };
    end
    if(N1361) begin
      { data_buf_r[491:490] } <= { data_mem_data_i[491:490] };
    end
    if(N1368) begin
      { data_buf_r[489:489] } <= { data_mem_data_i[489:489] };
    end
    if(N1374) begin
      { data_buf_r[488:481] } <= { data_mem_data_i[488:481] };
    end
    if(N1382) begin
      { data_buf_r[480:473] } <= { data_mem_data_i[480:473] };
    end
    if(N1388) begin
      { data_buf_r[412:393] } <= { data_mem_data_i[412:393] };
    end
    if(N1394) begin
      { data_buf_r[392:391] } <= { data_mem_data_i[392:391] };
    end
    if(N1401) begin
      { data_buf_r[390:390] } <= { data_mem_data_i[390:390] };
    end
    if(N1407) begin
      { data_buf_r[389:382] } <= { data_mem_data_i[389:382] };
    end
    if(N1415) begin
      { data_buf_r[381:374] } <= { data_mem_data_i[381:374] };
    end
    if(N1420) begin
      { data_buf_r[373:314] } <= { data_mem_data_i[373:314] };
    end
    if(N1426) begin
      { data_buf_r[313:294] } <= { data_mem_data_i[313:294] };
    end
    if(N1432) begin
      { data_buf_r[293:292] } <= { data_mem_data_i[293:292] };
    end
    if(N1439) begin
      { data_buf_r[291:291] } <= { data_mem_data_i[291:291] };
    end
    if(N1445) begin
      { data_buf_r[290:283] } <= { data_mem_data_i[290:283] };
    end
    if(N1453) begin
      { data_buf_r[282:275] } <= { data_mem_data_i[282:275] };
    end
    if(N1458) begin
      { data_buf_r[274:215] } <= { data_mem_data_i[274:215] };
    end
    if(N1464) begin
      { data_buf_r[214:195] } <= { data_mem_data_i[214:195] };
    end
    if(N1470) begin
      { data_buf_r[194:193] } <= { data_mem_data_i[194:193] };
    end
    if(N1477) begin
      { data_buf_r[192:192] } <= { data_mem_data_i[192:192] };
    end
    if(N1483) begin
      { data_buf_r[191:184] } <= { data_mem_data_i[191:184] };
    end
    if(N1491) begin
      { data_buf_r[183:176] } <= { data_mem_data_i[183:176] };
    end
    if(N1496) begin
      { data_buf_r[175:116] } <= { data_mem_data_i[175:116] };
    end
    if(N1502) begin
      { data_buf_r[115:96] } <= { data_mem_data_i[115:96] };
    end
    if(N1508) begin
      { data_buf_r[95:94] } <= { data_mem_data_i[95:94] };
    end
    if(N1515) begin
      { data_buf_r[93:93] } <= { data_mem_data_i[93:93] };
    end
    if(N1521) begin
      { data_buf_r[92:85] } <= { data_mem_data_i[92:85] };
    end
    if(N1529) begin
      { data_buf_r[84:77] } <= { data_mem_data_i[84:77] };
    end
    if(N1534) begin
      { data_buf_r[76:17], data_buf_r[4:4] } <= { data_mem_data_i[76:17], data_mem_data_i[4:4] };
    end
    if(N1540) begin
      { data_buf_r[16:5] } <= { data_mem_data_i[16:5] };
    end
    if(N1546) begin
      { data_buf_r[3:3] } <= { data_mem_data_i[3:3] };
    end
    if(N1552) begin
      { data_buf_r[2:2] } <= { data_mem_data_i[2:2] };
    end
    if(N1558) begin
      { data_buf_r[1:1] } <= { data_mem_data_i[1:1] };
    end
    if(N1570) begin
      { state_r[2:0] } <= { N1248, N1247, N1246 };
    end
    if(N1581) begin
      { sync_ack_count_r[0:0] } <= { N1249 };
    end
    if(N1586) begin
      tr_data_buffered_r <= N1250;
    end
    if(N1591) begin
      wb_data_buffered_r <= N1251;
      wb_data_read_r <= N1252;
      wb_dirty_cleared_r <= N1253;
    end
    if(N1604) begin
      invalidated_tag_r <= N1254;
    end
  end


endmodule



module bp_be_dcache_lce_data_cmd_num_cce_p1_num_lce_p2_data_width_p64_paddr_width_p22_lce_data_width_p512_ways_p8_sets_p64
(
  cce_data_received_o,
  tr_data_received_o,
  uncached_data_received_o,
  miss_addr_i,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_yumi_o,
  data_mem_pkt_v_o,
  data_mem_pkt_o,
  data_mem_pkt_yumi_i
);

  input [21:0] miss_addr_i;
  input [517:0] lce_data_cmd_i;
  output [522:0] data_mem_pkt_o;
  input lce_data_cmd_v_i;
  input data_mem_pkt_yumi_i;
  output cce_data_received_o;
  output tr_data_received_o;
  output uncached_data_received_o;
  output lce_data_cmd_yumi_o;
  output data_mem_pkt_v_o;
  wire [522:0] data_mem_pkt_o;
  wire cce_data_received_o,tr_data_received_o,uncached_data_received_o,
  lce_data_cmd_yumi_o,data_mem_pkt_v_o,data_mem_pkt_yumi_i,lce_data_cmd_v_i,N0,N1,N2,N3,N4,N5,N6,
  N7;
  assign data_mem_pkt_o[0] = 1'b0;
  assign data_mem_pkt_o[516] = lce_data_cmd_i[2];
  assign data_mem_pkt_o[515] = lce_data_cmd_i[1];
  assign data_mem_pkt_o[514] = lce_data_cmd_i[0];
  assign data_mem_pkt_o[513] = lce_data_cmd_i[517];
  assign data_mem_pkt_o[512] = lce_data_cmd_i[516];
  assign data_mem_pkt_o[511] = lce_data_cmd_i[515];
  assign data_mem_pkt_o[510] = lce_data_cmd_i[514];
  assign data_mem_pkt_o[509] = lce_data_cmd_i[513];
  assign data_mem_pkt_o[508] = lce_data_cmd_i[512];
  assign data_mem_pkt_o[507] = lce_data_cmd_i[511];
  assign data_mem_pkt_o[506] = lce_data_cmd_i[510];
  assign data_mem_pkt_o[505] = lce_data_cmd_i[509];
  assign data_mem_pkt_o[504] = lce_data_cmd_i[508];
  assign data_mem_pkt_o[503] = lce_data_cmd_i[507];
  assign data_mem_pkt_o[502] = lce_data_cmd_i[506];
  assign data_mem_pkt_o[501] = lce_data_cmd_i[505];
  assign data_mem_pkt_o[500] = lce_data_cmd_i[504];
  assign data_mem_pkt_o[499] = lce_data_cmd_i[503];
  assign data_mem_pkt_o[498] = lce_data_cmd_i[502];
  assign data_mem_pkt_o[497] = lce_data_cmd_i[501];
  assign data_mem_pkt_o[496] = lce_data_cmd_i[500];
  assign data_mem_pkt_o[495] = lce_data_cmd_i[499];
  assign data_mem_pkt_o[494] = lce_data_cmd_i[498];
  assign data_mem_pkt_o[493] = lce_data_cmd_i[497];
  assign data_mem_pkt_o[492] = lce_data_cmd_i[496];
  assign data_mem_pkt_o[491] = lce_data_cmd_i[495];
  assign data_mem_pkt_o[490] = lce_data_cmd_i[494];
  assign data_mem_pkt_o[489] = lce_data_cmd_i[493];
  assign data_mem_pkt_o[488] = lce_data_cmd_i[492];
  assign data_mem_pkt_o[487] = lce_data_cmd_i[491];
  assign data_mem_pkt_o[486] = lce_data_cmd_i[490];
  assign data_mem_pkt_o[485] = lce_data_cmd_i[489];
  assign data_mem_pkt_o[484] = lce_data_cmd_i[488];
  assign data_mem_pkt_o[483] = lce_data_cmd_i[487];
  assign data_mem_pkt_o[482] = lce_data_cmd_i[486];
  assign data_mem_pkt_o[481] = lce_data_cmd_i[485];
  assign data_mem_pkt_o[480] = lce_data_cmd_i[484];
  assign data_mem_pkt_o[479] = lce_data_cmd_i[483];
  assign data_mem_pkt_o[478] = lce_data_cmd_i[482];
  assign data_mem_pkt_o[477] = lce_data_cmd_i[481];
  assign data_mem_pkt_o[476] = lce_data_cmd_i[480];
  assign data_mem_pkt_o[475] = lce_data_cmd_i[479];
  assign data_mem_pkt_o[474] = lce_data_cmd_i[478];
  assign data_mem_pkt_o[473] = lce_data_cmd_i[477];
  assign data_mem_pkt_o[472] = lce_data_cmd_i[476];
  assign data_mem_pkt_o[471] = lce_data_cmd_i[475];
  assign data_mem_pkt_o[470] = lce_data_cmd_i[474];
  assign data_mem_pkt_o[469] = lce_data_cmd_i[473];
  assign data_mem_pkt_o[468] = lce_data_cmd_i[472];
  assign data_mem_pkt_o[467] = lce_data_cmd_i[471];
  assign data_mem_pkt_o[466] = lce_data_cmd_i[470];
  assign data_mem_pkt_o[465] = lce_data_cmd_i[469];
  assign data_mem_pkt_o[464] = lce_data_cmd_i[468];
  assign data_mem_pkt_o[463] = lce_data_cmd_i[467];
  assign data_mem_pkt_o[462] = lce_data_cmd_i[466];
  assign data_mem_pkt_o[461] = lce_data_cmd_i[465];
  assign data_mem_pkt_o[460] = lce_data_cmd_i[464];
  assign data_mem_pkt_o[459] = lce_data_cmd_i[463];
  assign data_mem_pkt_o[458] = lce_data_cmd_i[462];
  assign data_mem_pkt_o[457] = lce_data_cmd_i[461];
  assign data_mem_pkt_o[456] = lce_data_cmd_i[460];
  assign data_mem_pkt_o[455] = lce_data_cmd_i[459];
  assign data_mem_pkt_o[454] = lce_data_cmd_i[458];
  assign data_mem_pkt_o[453] = lce_data_cmd_i[457];
  assign data_mem_pkt_o[452] = lce_data_cmd_i[456];
  assign data_mem_pkt_o[451] = lce_data_cmd_i[455];
  assign data_mem_pkt_o[450] = lce_data_cmd_i[454];
  assign data_mem_pkt_o[449] = lce_data_cmd_i[453];
  assign data_mem_pkt_o[448] = lce_data_cmd_i[452];
  assign data_mem_pkt_o[447] = lce_data_cmd_i[451];
  assign data_mem_pkt_o[446] = lce_data_cmd_i[450];
  assign data_mem_pkt_o[445] = lce_data_cmd_i[449];
  assign data_mem_pkt_o[444] = lce_data_cmd_i[448];
  assign data_mem_pkt_o[443] = lce_data_cmd_i[447];
  assign data_mem_pkt_o[442] = lce_data_cmd_i[446];
  assign data_mem_pkt_o[441] = lce_data_cmd_i[445];
  assign data_mem_pkt_o[440] = lce_data_cmd_i[444];
  assign data_mem_pkt_o[439] = lce_data_cmd_i[443];
  assign data_mem_pkt_o[438] = lce_data_cmd_i[442];
  assign data_mem_pkt_o[437] = lce_data_cmd_i[441];
  assign data_mem_pkt_o[436] = lce_data_cmd_i[440];
  assign data_mem_pkt_o[435] = lce_data_cmd_i[439];
  assign data_mem_pkt_o[434] = lce_data_cmd_i[438];
  assign data_mem_pkt_o[433] = lce_data_cmd_i[437];
  assign data_mem_pkt_o[432] = lce_data_cmd_i[436];
  assign data_mem_pkt_o[431] = lce_data_cmd_i[435];
  assign data_mem_pkt_o[430] = lce_data_cmd_i[434];
  assign data_mem_pkt_o[429] = lce_data_cmd_i[433];
  assign data_mem_pkt_o[428] = lce_data_cmd_i[432];
  assign data_mem_pkt_o[427] = lce_data_cmd_i[431];
  assign data_mem_pkt_o[426] = lce_data_cmd_i[430];
  assign data_mem_pkt_o[425] = lce_data_cmd_i[429];
  assign data_mem_pkt_o[424] = lce_data_cmd_i[428];
  assign data_mem_pkt_o[423] = lce_data_cmd_i[427];
  assign data_mem_pkt_o[422] = lce_data_cmd_i[426];
  assign data_mem_pkt_o[421] = lce_data_cmd_i[425];
  assign data_mem_pkt_o[420] = lce_data_cmd_i[424];
  assign data_mem_pkt_o[419] = lce_data_cmd_i[423];
  assign data_mem_pkt_o[418] = lce_data_cmd_i[422];
  assign data_mem_pkt_o[417] = lce_data_cmd_i[421];
  assign data_mem_pkt_o[416] = lce_data_cmd_i[420];
  assign data_mem_pkt_o[415] = lce_data_cmd_i[419];
  assign data_mem_pkt_o[414] = lce_data_cmd_i[418];
  assign data_mem_pkt_o[413] = lce_data_cmd_i[417];
  assign data_mem_pkt_o[412] = lce_data_cmd_i[416];
  assign data_mem_pkt_o[411] = lce_data_cmd_i[415];
  assign data_mem_pkt_o[410] = lce_data_cmd_i[414];
  assign data_mem_pkt_o[409] = lce_data_cmd_i[413];
  assign data_mem_pkt_o[408] = lce_data_cmd_i[412];
  assign data_mem_pkt_o[407] = lce_data_cmd_i[411];
  assign data_mem_pkt_o[406] = lce_data_cmd_i[410];
  assign data_mem_pkt_o[405] = lce_data_cmd_i[409];
  assign data_mem_pkt_o[404] = lce_data_cmd_i[408];
  assign data_mem_pkt_o[403] = lce_data_cmd_i[407];
  assign data_mem_pkt_o[402] = lce_data_cmd_i[406];
  assign data_mem_pkt_o[401] = lce_data_cmd_i[405];
  assign data_mem_pkt_o[400] = lce_data_cmd_i[404];
  assign data_mem_pkt_o[399] = lce_data_cmd_i[403];
  assign data_mem_pkt_o[398] = lce_data_cmd_i[402];
  assign data_mem_pkt_o[397] = lce_data_cmd_i[401];
  assign data_mem_pkt_o[396] = lce_data_cmd_i[400];
  assign data_mem_pkt_o[395] = lce_data_cmd_i[399];
  assign data_mem_pkt_o[394] = lce_data_cmd_i[398];
  assign data_mem_pkt_o[393] = lce_data_cmd_i[397];
  assign data_mem_pkt_o[392] = lce_data_cmd_i[396];
  assign data_mem_pkt_o[391] = lce_data_cmd_i[395];
  assign data_mem_pkt_o[390] = lce_data_cmd_i[394];
  assign data_mem_pkt_o[389] = lce_data_cmd_i[393];
  assign data_mem_pkt_o[388] = lce_data_cmd_i[392];
  assign data_mem_pkt_o[387] = lce_data_cmd_i[391];
  assign data_mem_pkt_o[386] = lce_data_cmd_i[390];
  assign data_mem_pkt_o[385] = lce_data_cmd_i[389];
  assign data_mem_pkt_o[384] = lce_data_cmd_i[388];
  assign data_mem_pkt_o[383] = lce_data_cmd_i[387];
  assign data_mem_pkt_o[382] = lce_data_cmd_i[386];
  assign data_mem_pkt_o[381] = lce_data_cmd_i[385];
  assign data_mem_pkt_o[380] = lce_data_cmd_i[384];
  assign data_mem_pkt_o[379] = lce_data_cmd_i[383];
  assign data_mem_pkt_o[378] = lce_data_cmd_i[382];
  assign data_mem_pkt_o[377] = lce_data_cmd_i[381];
  assign data_mem_pkt_o[376] = lce_data_cmd_i[380];
  assign data_mem_pkt_o[375] = lce_data_cmd_i[379];
  assign data_mem_pkt_o[374] = lce_data_cmd_i[378];
  assign data_mem_pkt_o[373] = lce_data_cmd_i[377];
  assign data_mem_pkt_o[372] = lce_data_cmd_i[376];
  assign data_mem_pkt_o[371] = lce_data_cmd_i[375];
  assign data_mem_pkt_o[370] = lce_data_cmd_i[374];
  assign data_mem_pkt_o[369] = lce_data_cmd_i[373];
  assign data_mem_pkt_o[368] = lce_data_cmd_i[372];
  assign data_mem_pkt_o[367] = lce_data_cmd_i[371];
  assign data_mem_pkt_o[366] = lce_data_cmd_i[370];
  assign data_mem_pkt_o[365] = lce_data_cmd_i[369];
  assign data_mem_pkt_o[364] = lce_data_cmd_i[368];
  assign data_mem_pkt_o[363] = lce_data_cmd_i[367];
  assign data_mem_pkt_o[362] = lce_data_cmd_i[366];
  assign data_mem_pkt_o[361] = lce_data_cmd_i[365];
  assign data_mem_pkt_o[360] = lce_data_cmd_i[364];
  assign data_mem_pkt_o[359] = lce_data_cmd_i[363];
  assign data_mem_pkt_o[358] = lce_data_cmd_i[362];
  assign data_mem_pkt_o[357] = lce_data_cmd_i[361];
  assign data_mem_pkt_o[356] = lce_data_cmd_i[360];
  assign data_mem_pkt_o[355] = lce_data_cmd_i[359];
  assign data_mem_pkt_o[354] = lce_data_cmd_i[358];
  assign data_mem_pkt_o[353] = lce_data_cmd_i[357];
  assign data_mem_pkt_o[352] = lce_data_cmd_i[356];
  assign data_mem_pkt_o[351] = lce_data_cmd_i[355];
  assign data_mem_pkt_o[350] = lce_data_cmd_i[354];
  assign data_mem_pkt_o[349] = lce_data_cmd_i[353];
  assign data_mem_pkt_o[348] = lce_data_cmd_i[352];
  assign data_mem_pkt_o[347] = lce_data_cmd_i[351];
  assign data_mem_pkt_o[346] = lce_data_cmd_i[350];
  assign data_mem_pkt_o[345] = lce_data_cmd_i[349];
  assign data_mem_pkt_o[344] = lce_data_cmd_i[348];
  assign data_mem_pkt_o[343] = lce_data_cmd_i[347];
  assign data_mem_pkt_o[342] = lce_data_cmd_i[346];
  assign data_mem_pkt_o[341] = lce_data_cmd_i[345];
  assign data_mem_pkt_o[340] = lce_data_cmd_i[344];
  assign data_mem_pkt_o[339] = lce_data_cmd_i[343];
  assign data_mem_pkt_o[338] = lce_data_cmd_i[342];
  assign data_mem_pkt_o[337] = lce_data_cmd_i[341];
  assign data_mem_pkt_o[336] = lce_data_cmd_i[340];
  assign data_mem_pkt_o[335] = lce_data_cmd_i[339];
  assign data_mem_pkt_o[334] = lce_data_cmd_i[338];
  assign data_mem_pkt_o[333] = lce_data_cmd_i[337];
  assign data_mem_pkt_o[332] = lce_data_cmd_i[336];
  assign data_mem_pkt_o[331] = lce_data_cmd_i[335];
  assign data_mem_pkt_o[330] = lce_data_cmd_i[334];
  assign data_mem_pkt_o[329] = lce_data_cmd_i[333];
  assign data_mem_pkt_o[328] = lce_data_cmd_i[332];
  assign data_mem_pkt_o[327] = lce_data_cmd_i[331];
  assign data_mem_pkt_o[326] = lce_data_cmd_i[330];
  assign data_mem_pkt_o[325] = lce_data_cmd_i[329];
  assign data_mem_pkt_o[324] = lce_data_cmd_i[328];
  assign data_mem_pkt_o[323] = lce_data_cmd_i[327];
  assign data_mem_pkt_o[322] = lce_data_cmd_i[326];
  assign data_mem_pkt_o[321] = lce_data_cmd_i[325];
  assign data_mem_pkt_o[320] = lce_data_cmd_i[324];
  assign data_mem_pkt_o[319] = lce_data_cmd_i[323];
  assign data_mem_pkt_o[318] = lce_data_cmd_i[322];
  assign data_mem_pkt_o[317] = lce_data_cmd_i[321];
  assign data_mem_pkt_o[316] = lce_data_cmd_i[320];
  assign data_mem_pkt_o[315] = lce_data_cmd_i[319];
  assign data_mem_pkt_o[314] = lce_data_cmd_i[318];
  assign data_mem_pkt_o[313] = lce_data_cmd_i[317];
  assign data_mem_pkt_o[312] = lce_data_cmd_i[316];
  assign data_mem_pkt_o[311] = lce_data_cmd_i[315];
  assign data_mem_pkt_o[310] = lce_data_cmd_i[314];
  assign data_mem_pkt_o[309] = lce_data_cmd_i[313];
  assign data_mem_pkt_o[308] = lce_data_cmd_i[312];
  assign data_mem_pkt_o[307] = lce_data_cmd_i[311];
  assign data_mem_pkt_o[306] = lce_data_cmd_i[310];
  assign data_mem_pkt_o[305] = lce_data_cmd_i[309];
  assign data_mem_pkt_o[304] = lce_data_cmd_i[308];
  assign data_mem_pkt_o[303] = lce_data_cmd_i[307];
  assign data_mem_pkt_o[302] = lce_data_cmd_i[306];
  assign data_mem_pkt_o[301] = lce_data_cmd_i[305];
  assign data_mem_pkt_o[300] = lce_data_cmd_i[304];
  assign data_mem_pkt_o[299] = lce_data_cmd_i[303];
  assign data_mem_pkt_o[298] = lce_data_cmd_i[302];
  assign data_mem_pkt_o[297] = lce_data_cmd_i[301];
  assign data_mem_pkt_o[296] = lce_data_cmd_i[300];
  assign data_mem_pkt_o[295] = lce_data_cmd_i[299];
  assign data_mem_pkt_o[294] = lce_data_cmd_i[298];
  assign data_mem_pkt_o[293] = lce_data_cmd_i[297];
  assign data_mem_pkt_o[292] = lce_data_cmd_i[296];
  assign data_mem_pkt_o[291] = lce_data_cmd_i[295];
  assign data_mem_pkt_o[290] = lce_data_cmd_i[294];
  assign data_mem_pkt_o[289] = lce_data_cmd_i[293];
  assign data_mem_pkt_o[288] = lce_data_cmd_i[292];
  assign data_mem_pkt_o[287] = lce_data_cmd_i[291];
  assign data_mem_pkt_o[286] = lce_data_cmd_i[290];
  assign data_mem_pkt_o[285] = lce_data_cmd_i[289];
  assign data_mem_pkt_o[284] = lce_data_cmd_i[288];
  assign data_mem_pkt_o[283] = lce_data_cmd_i[287];
  assign data_mem_pkt_o[282] = lce_data_cmd_i[286];
  assign data_mem_pkt_o[281] = lce_data_cmd_i[285];
  assign data_mem_pkt_o[280] = lce_data_cmd_i[284];
  assign data_mem_pkt_o[279] = lce_data_cmd_i[283];
  assign data_mem_pkt_o[278] = lce_data_cmd_i[282];
  assign data_mem_pkt_o[277] = lce_data_cmd_i[281];
  assign data_mem_pkt_o[276] = lce_data_cmd_i[280];
  assign data_mem_pkt_o[275] = lce_data_cmd_i[279];
  assign data_mem_pkt_o[274] = lce_data_cmd_i[278];
  assign data_mem_pkt_o[273] = lce_data_cmd_i[277];
  assign data_mem_pkt_o[272] = lce_data_cmd_i[276];
  assign data_mem_pkt_o[271] = lce_data_cmd_i[275];
  assign data_mem_pkt_o[270] = lce_data_cmd_i[274];
  assign data_mem_pkt_o[269] = lce_data_cmd_i[273];
  assign data_mem_pkt_o[268] = lce_data_cmd_i[272];
  assign data_mem_pkt_o[267] = lce_data_cmd_i[271];
  assign data_mem_pkt_o[266] = lce_data_cmd_i[270];
  assign data_mem_pkt_o[265] = lce_data_cmd_i[269];
  assign data_mem_pkt_o[264] = lce_data_cmd_i[268];
  assign data_mem_pkt_o[263] = lce_data_cmd_i[267];
  assign data_mem_pkt_o[262] = lce_data_cmd_i[266];
  assign data_mem_pkt_o[261] = lce_data_cmd_i[265];
  assign data_mem_pkt_o[260] = lce_data_cmd_i[264];
  assign data_mem_pkt_o[259] = lce_data_cmd_i[263];
  assign data_mem_pkt_o[258] = lce_data_cmd_i[262];
  assign data_mem_pkt_o[257] = lce_data_cmd_i[261];
  assign data_mem_pkt_o[256] = lce_data_cmd_i[260];
  assign data_mem_pkt_o[255] = lce_data_cmd_i[259];
  assign data_mem_pkt_o[254] = lce_data_cmd_i[258];
  assign data_mem_pkt_o[253] = lce_data_cmd_i[257];
  assign data_mem_pkt_o[252] = lce_data_cmd_i[256];
  assign data_mem_pkt_o[251] = lce_data_cmd_i[255];
  assign data_mem_pkt_o[250] = lce_data_cmd_i[254];
  assign data_mem_pkt_o[249] = lce_data_cmd_i[253];
  assign data_mem_pkt_o[248] = lce_data_cmd_i[252];
  assign data_mem_pkt_o[247] = lce_data_cmd_i[251];
  assign data_mem_pkt_o[246] = lce_data_cmd_i[250];
  assign data_mem_pkt_o[245] = lce_data_cmd_i[249];
  assign data_mem_pkt_o[244] = lce_data_cmd_i[248];
  assign data_mem_pkt_o[243] = lce_data_cmd_i[247];
  assign data_mem_pkt_o[242] = lce_data_cmd_i[246];
  assign data_mem_pkt_o[241] = lce_data_cmd_i[245];
  assign data_mem_pkt_o[240] = lce_data_cmd_i[244];
  assign data_mem_pkt_o[239] = lce_data_cmd_i[243];
  assign data_mem_pkt_o[238] = lce_data_cmd_i[242];
  assign data_mem_pkt_o[237] = lce_data_cmd_i[241];
  assign data_mem_pkt_o[236] = lce_data_cmd_i[240];
  assign data_mem_pkt_o[235] = lce_data_cmd_i[239];
  assign data_mem_pkt_o[234] = lce_data_cmd_i[238];
  assign data_mem_pkt_o[233] = lce_data_cmd_i[237];
  assign data_mem_pkt_o[232] = lce_data_cmd_i[236];
  assign data_mem_pkt_o[231] = lce_data_cmd_i[235];
  assign data_mem_pkt_o[230] = lce_data_cmd_i[234];
  assign data_mem_pkt_o[229] = lce_data_cmd_i[233];
  assign data_mem_pkt_o[228] = lce_data_cmd_i[232];
  assign data_mem_pkt_o[227] = lce_data_cmd_i[231];
  assign data_mem_pkt_o[226] = lce_data_cmd_i[230];
  assign data_mem_pkt_o[225] = lce_data_cmd_i[229];
  assign data_mem_pkt_o[224] = lce_data_cmd_i[228];
  assign data_mem_pkt_o[223] = lce_data_cmd_i[227];
  assign data_mem_pkt_o[222] = lce_data_cmd_i[226];
  assign data_mem_pkt_o[221] = lce_data_cmd_i[225];
  assign data_mem_pkt_o[220] = lce_data_cmd_i[224];
  assign data_mem_pkt_o[219] = lce_data_cmd_i[223];
  assign data_mem_pkt_o[218] = lce_data_cmd_i[222];
  assign data_mem_pkt_o[217] = lce_data_cmd_i[221];
  assign data_mem_pkt_o[216] = lce_data_cmd_i[220];
  assign data_mem_pkt_o[215] = lce_data_cmd_i[219];
  assign data_mem_pkt_o[214] = lce_data_cmd_i[218];
  assign data_mem_pkt_o[213] = lce_data_cmd_i[217];
  assign data_mem_pkt_o[212] = lce_data_cmd_i[216];
  assign data_mem_pkt_o[211] = lce_data_cmd_i[215];
  assign data_mem_pkt_o[210] = lce_data_cmd_i[214];
  assign data_mem_pkt_o[209] = lce_data_cmd_i[213];
  assign data_mem_pkt_o[208] = lce_data_cmd_i[212];
  assign data_mem_pkt_o[207] = lce_data_cmd_i[211];
  assign data_mem_pkt_o[206] = lce_data_cmd_i[210];
  assign data_mem_pkt_o[205] = lce_data_cmd_i[209];
  assign data_mem_pkt_o[204] = lce_data_cmd_i[208];
  assign data_mem_pkt_o[203] = lce_data_cmd_i[207];
  assign data_mem_pkt_o[202] = lce_data_cmd_i[206];
  assign data_mem_pkt_o[201] = lce_data_cmd_i[205];
  assign data_mem_pkt_o[200] = lce_data_cmd_i[204];
  assign data_mem_pkt_o[199] = lce_data_cmd_i[203];
  assign data_mem_pkt_o[198] = lce_data_cmd_i[202];
  assign data_mem_pkt_o[197] = lce_data_cmd_i[201];
  assign data_mem_pkt_o[196] = lce_data_cmd_i[200];
  assign data_mem_pkt_o[195] = lce_data_cmd_i[199];
  assign data_mem_pkt_o[194] = lce_data_cmd_i[198];
  assign data_mem_pkt_o[193] = lce_data_cmd_i[197];
  assign data_mem_pkt_o[192] = lce_data_cmd_i[196];
  assign data_mem_pkt_o[191] = lce_data_cmd_i[195];
  assign data_mem_pkt_o[190] = lce_data_cmd_i[194];
  assign data_mem_pkt_o[189] = lce_data_cmd_i[193];
  assign data_mem_pkt_o[188] = lce_data_cmd_i[192];
  assign data_mem_pkt_o[187] = lce_data_cmd_i[191];
  assign data_mem_pkt_o[186] = lce_data_cmd_i[190];
  assign data_mem_pkt_o[185] = lce_data_cmd_i[189];
  assign data_mem_pkt_o[184] = lce_data_cmd_i[188];
  assign data_mem_pkt_o[183] = lce_data_cmd_i[187];
  assign data_mem_pkt_o[182] = lce_data_cmd_i[186];
  assign data_mem_pkt_o[181] = lce_data_cmd_i[185];
  assign data_mem_pkt_o[180] = lce_data_cmd_i[184];
  assign data_mem_pkt_o[179] = lce_data_cmd_i[183];
  assign data_mem_pkt_o[178] = lce_data_cmd_i[182];
  assign data_mem_pkt_o[177] = lce_data_cmd_i[181];
  assign data_mem_pkt_o[176] = lce_data_cmd_i[180];
  assign data_mem_pkt_o[175] = lce_data_cmd_i[179];
  assign data_mem_pkt_o[174] = lce_data_cmd_i[178];
  assign data_mem_pkt_o[173] = lce_data_cmd_i[177];
  assign data_mem_pkt_o[172] = lce_data_cmd_i[176];
  assign data_mem_pkt_o[171] = lce_data_cmd_i[175];
  assign data_mem_pkt_o[170] = lce_data_cmd_i[174];
  assign data_mem_pkt_o[169] = lce_data_cmd_i[173];
  assign data_mem_pkt_o[168] = lce_data_cmd_i[172];
  assign data_mem_pkt_o[167] = lce_data_cmd_i[171];
  assign data_mem_pkt_o[166] = lce_data_cmd_i[170];
  assign data_mem_pkt_o[165] = lce_data_cmd_i[169];
  assign data_mem_pkt_o[164] = lce_data_cmd_i[168];
  assign data_mem_pkt_o[163] = lce_data_cmd_i[167];
  assign data_mem_pkt_o[162] = lce_data_cmd_i[166];
  assign data_mem_pkt_o[161] = lce_data_cmd_i[165];
  assign data_mem_pkt_o[160] = lce_data_cmd_i[164];
  assign data_mem_pkt_o[159] = lce_data_cmd_i[163];
  assign data_mem_pkt_o[158] = lce_data_cmd_i[162];
  assign data_mem_pkt_o[157] = lce_data_cmd_i[161];
  assign data_mem_pkt_o[156] = lce_data_cmd_i[160];
  assign data_mem_pkt_o[155] = lce_data_cmd_i[159];
  assign data_mem_pkt_o[154] = lce_data_cmd_i[158];
  assign data_mem_pkt_o[153] = lce_data_cmd_i[157];
  assign data_mem_pkt_o[152] = lce_data_cmd_i[156];
  assign data_mem_pkt_o[151] = lce_data_cmd_i[155];
  assign data_mem_pkt_o[150] = lce_data_cmd_i[154];
  assign data_mem_pkt_o[149] = lce_data_cmd_i[153];
  assign data_mem_pkt_o[148] = lce_data_cmd_i[152];
  assign data_mem_pkt_o[147] = lce_data_cmd_i[151];
  assign data_mem_pkt_o[146] = lce_data_cmd_i[150];
  assign data_mem_pkt_o[145] = lce_data_cmd_i[149];
  assign data_mem_pkt_o[144] = lce_data_cmd_i[148];
  assign data_mem_pkt_o[143] = lce_data_cmd_i[147];
  assign data_mem_pkt_o[142] = lce_data_cmd_i[146];
  assign data_mem_pkt_o[141] = lce_data_cmd_i[145];
  assign data_mem_pkt_o[140] = lce_data_cmd_i[144];
  assign data_mem_pkt_o[139] = lce_data_cmd_i[143];
  assign data_mem_pkt_o[138] = lce_data_cmd_i[142];
  assign data_mem_pkt_o[137] = lce_data_cmd_i[141];
  assign data_mem_pkt_o[136] = lce_data_cmd_i[140];
  assign data_mem_pkt_o[135] = lce_data_cmd_i[139];
  assign data_mem_pkt_o[134] = lce_data_cmd_i[138];
  assign data_mem_pkt_o[133] = lce_data_cmd_i[137];
  assign data_mem_pkt_o[132] = lce_data_cmd_i[136];
  assign data_mem_pkt_o[131] = lce_data_cmd_i[135];
  assign data_mem_pkt_o[130] = lce_data_cmd_i[134];
  assign data_mem_pkt_o[129] = lce_data_cmd_i[133];
  assign data_mem_pkt_o[128] = lce_data_cmd_i[132];
  assign data_mem_pkt_o[127] = lce_data_cmd_i[131];
  assign data_mem_pkt_o[126] = lce_data_cmd_i[130];
  assign data_mem_pkt_o[125] = lce_data_cmd_i[129];
  assign data_mem_pkt_o[124] = lce_data_cmd_i[128];
  assign data_mem_pkt_o[123] = lce_data_cmd_i[127];
  assign data_mem_pkt_o[122] = lce_data_cmd_i[126];
  assign data_mem_pkt_o[121] = lce_data_cmd_i[125];
  assign data_mem_pkt_o[120] = lce_data_cmd_i[124];
  assign data_mem_pkt_o[119] = lce_data_cmd_i[123];
  assign data_mem_pkt_o[118] = lce_data_cmd_i[122];
  assign data_mem_pkt_o[117] = lce_data_cmd_i[121];
  assign data_mem_pkt_o[116] = lce_data_cmd_i[120];
  assign data_mem_pkt_o[115] = lce_data_cmd_i[119];
  assign data_mem_pkt_o[114] = lce_data_cmd_i[118];
  assign data_mem_pkt_o[113] = lce_data_cmd_i[117];
  assign data_mem_pkt_o[112] = lce_data_cmd_i[116];
  assign data_mem_pkt_o[111] = lce_data_cmd_i[115];
  assign data_mem_pkt_o[110] = lce_data_cmd_i[114];
  assign data_mem_pkt_o[109] = lce_data_cmd_i[113];
  assign data_mem_pkt_o[108] = lce_data_cmd_i[112];
  assign data_mem_pkt_o[107] = lce_data_cmd_i[111];
  assign data_mem_pkt_o[106] = lce_data_cmd_i[110];
  assign data_mem_pkt_o[105] = lce_data_cmd_i[109];
  assign data_mem_pkt_o[104] = lce_data_cmd_i[108];
  assign data_mem_pkt_o[103] = lce_data_cmd_i[107];
  assign data_mem_pkt_o[102] = lce_data_cmd_i[106];
  assign data_mem_pkt_o[101] = lce_data_cmd_i[105];
  assign data_mem_pkt_o[100] = lce_data_cmd_i[104];
  assign data_mem_pkt_o[99] = lce_data_cmd_i[103];
  assign data_mem_pkt_o[98] = lce_data_cmd_i[102];
  assign data_mem_pkt_o[97] = lce_data_cmd_i[101];
  assign data_mem_pkt_o[96] = lce_data_cmd_i[100];
  assign data_mem_pkt_o[95] = lce_data_cmd_i[99];
  assign data_mem_pkt_o[94] = lce_data_cmd_i[98];
  assign data_mem_pkt_o[93] = lce_data_cmd_i[97];
  assign data_mem_pkt_o[92] = lce_data_cmd_i[96];
  assign data_mem_pkt_o[91] = lce_data_cmd_i[95];
  assign data_mem_pkt_o[90] = lce_data_cmd_i[94];
  assign data_mem_pkt_o[89] = lce_data_cmd_i[93];
  assign data_mem_pkt_o[88] = lce_data_cmd_i[92];
  assign data_mem_pkt_o[87] = lce_data_cmd_i[91];
  assign data_mem_pkt_o[86] = lce_data_cmd_i[90];
  assign data_mem_pkt_o[85] = lce_data_cmd_i[89];
  assign data_mem_pkt_o[84] = lce_data_cmd_i[88];
  assign data_mem_pkt_o[83] = lce_data_cmd_i[87];
  assign data_mem_pkt_o[82] = lce_data_cmd_i[86];
  assign data_mem_pkt_o[81] = lce_data_cmd_i[85];
  assign data_mem_pkt_o[80] = lce_data_cmd_i[84];
  assign data_mem_pkt_o[79] = lce_data_cmd_i[83];
  assign data_mem_pkt_o[78] = lce_data_cmd_i[82];
  assign data_mem_pkt_o[77] = lce_data_cmd_i[81];
  assign data_mem_pkt_o[76] = lce_data_cmd_i[80];
  assign data_mem_pkt_o[75] = lce_data_cmd_i[79];
  assign data_mem_pkt_o[74] = lce_data_cmd_i[78];
  assign data_mem_pkt_o[73] = lce_data_cmd_i[77];
  assign data_mem_pkt_o[72] = lce_data_cmd_i[76];
  assign data_mem_pkt_o[71] = lce_data_cmd_i[75];
  assign data_mem_pkt_o[70] = lce_data_cmd_i[74];
  assign data_mem_pkt_o[69] = lce_data_cmd_i[73];
  assign data_mem_pkt_o[68] = lce_data_cmd_i[72];
  assign data_mem_pkt_o[67] = lce_data_cmd_i[71];
  assign data_mem_pkt_o[66] = lce_data_cmd_i[70];
  assign data_mem_pkt_o[65] = lce_data_cmd_i[69];
  assign data_mem_pkt_o[64] = lce_data_cmd_i[68];
  assign data_mem_pkt_o[63] = lce_data_cmd_i[67];
  assign data_mem_pkt_o[62] = lce_data_cmd_i[66];
  assign data_mem_pkt_o[61] = lce_data_cmd_i[65];
  assign data_mem_pkt_o[60] = lce_data_cmd_i[64];
  assign data_mem_pkt_o[59] = lce_data_cmd_i[63];
  assign data_mem_pkt_o[58] = lce_data_cmd_i[62];
  assign data_mem_pkt_o[57] = lce_data_cmd_i[61];
  assign data_mem_pkt_o[56] = lce_data_cmd_i[60];
  assign data_mem_pkt_o[55] = lce_data_cmd_i[59];
  assign data_mem_pkt_o[54] = lce_data_cmd_i[58];
  assign data_mem_pkt_o[53] = lce_data_cmd_i[57];
  assign data_mem_pkt_o[52] = lce_data_cmd_i[56];
  assign data_mem_pkt_o[51] = lce_data_cmd_i[55];
  assign data_mem_pkt_o[50] = lce_data_cmd_i[54];
  assign data_mem_pkt_o[49] = lce_data_cmd_i[53];
  assign data_mem_pkt_o[48] = lce_data_cmd_i[52];
  assign data_mem_pkt_o[47] = lce_data_cmd_i[51];
  assign data_mem_pkt_o[46] = lce_data_cmd_i[50];
  assign data_mem_pkt_o[45] = lce_data_cmd_i[49];
  assign data_mem_pkt_o[44] = lce_data_cmd_i[48];
  assign data_mem_pkt_o[43] = lce_data_cmd_i[47];
  assign data_mem_pkt_o[42] = lce_data_cmd_i[46];
  assign data_mem_pkt_o[41] = lce_data_cmd_i[45];
  assign data_mem_pkt_o[40] = lce_data_cmd_i[44];
  assign data_mem_pkt_o[39] = lce_data_cmd_i[43];
  assign data_mem_pkt_o[38] = lce_data_cmd_i[42];
  assign data_mem_pkt_o[37] = lce_data_cmd_i[41];
  assign data_mem_pkt_o[36] = lce_data_cmd_i[40];
  assign data_mem_pkt_o[35] = lce_data_cmd_i[39];
  assign data_mem_pkt_o[34] = lce_data_cmd_i[38];
  assign data_mem_pkt_o[33] = lce_data_cmd_i[37];
  assign data_mem_pkt_o[32] = lce_data_cmd_i[36];
  assign data_mem_pkt_o[31] = lce_data_cmd_i[35];
  assign data_mem_pkt_o[30] = lce_data_cmd_i[34];
  assign data_mem_pkt_o[29] = lce_data_cmd_i[33];
  assign data_mem_pkt_o[28] = lce_data_cmd_i[32];
  assign data_mem_pkt_o[27] = lce_data_cmd_i[31];
  assign data_mem_pkt_o[26] = lce_data_cmd_i[30];
  assign data_mem_pkt_o[25] = lce_data_cmd_i[29];
  assign data_mem_pkt_o[24] = lce_data_cmd_i[28];
  assign data_mem_pkt_o[23] = lce_data_cmd_i[27];
  assign data_mem_pkt_o[22] = lce_data_cmd_i[26];
  assign data_mem_pkt_o[21] = lce_data_cmd_i[25];
  assign data_mem_pkt_o[20] = lce_data_cmd_i[24];
  assign data_mem_pkt_o[19] = lce_data_cmd_i[23];
  assign data_mem_pkt_o[18] = lce_data_cmd_i[22];
  assign data_mem_pkt_o[17] = lce_data_cmd_i[21];
  assign data_mem_pkt_o[16] = lce_data_cmd_i[20];
  assign data_mem_pkt_o[15] = lce_data_cmd_i[19];
  assign data_mem_pkt_o[14] = lce_data_cmd_i[18];
  assign data_mem_pkt_o[13] = lce_data_cmd_i[17];
  assign data_mem_pkt_o[12] = lce_data_cmd_i[16];
  assign data_mem_pkt_o[11] = lce_data_cmd_i[15];
  assign data_mem_pkt_o[10] = lce_data_cmd_i[14];
  assign data_mem_pkt_o[9] = lce_data_cmd_i[13];
  assign data_mem_pkt_o[8] = lce_data_cmd_i[12];
  assign data_mem_pkt_o[7] = lce_data_cmd_i[11];
  assign data_mem_pkt_o[6] = lce_data_cmd_i[10];
  assign data_mem_pkt_o[5] = lce_data_cmd_i[9];
  assign data_mem_pkt_o[4] = lce_data_cmd_i[8];
  assign data_mem_pkt_o[3] = lce_data_cmd_i[7];
  assign data_mem_pkt_o[2] = lce_data_cmd_i[6];
  assign lce_data_cmd_yumi_o = data_mem_pkt_yumi_i;
  assign data_mem_pkt_v_o = lce_data_cmd_v_i;
  assign data_mem_pkt_o[522] = miss_addr_i[11];
  assign data_mem_pkt_o[521] = miss_addr_i[10];
  assign data_mem_pkt_o[520] = miss_addr_i[9];
  assign data_mem_pkt_o[519] = miss_addr_i[8];
  assign data_mem_pkt_o[518] = miss_addr_i[7];
  assign data_mem_pkt_o[517] = miss_addr_i[6];
  assign N0 = ~lce_data_cmd_i[3];
  assign N1 = N0 | lce_data_cmd_i[4];
  assign N2 = ~N1;
  assign N3 = lce_data_cmd_i[3] | lce_data_cmd_i[4];
  assign N4 = ~N3;
  assign N5 = ~lce_data_cmd_i[4];
  assign N6 = lce_data_cmd_i[3] | N5;
  assign N7 = ~N6;
  assign data_mem_pkt_o[1] = N7;
  assign cce_data_received_o = data_mem_pkt_yumi_i & N2;
  assign tr_data_received_o = data_mem_pkt_yumi_i & N4;
  assign uncached_data_received_o = data_mem_pkt_yumi_i & N7;

endmodule



module bp_be_dcache_lce_data_width_p64_paddr_width_p22_lce_data_width_p512_sets_p64_ways_p8_num_cce_p1_num_lce_p2
(
  clk_i,
  reset_i,
  lce_id_i,
  ready_o,
  cache_miss_o,
  load_miss_i,
  store_miss_i,
  uncached_load_req_i,
  uncached_store_req_i,
  miss_addr_i,
  store_data_i,
  size_op_i,
  data_mem_pkt_v_o,
  data_mem_pkt_o,
  data_mem_data_i,
  data_mem_pkt_yumi_i,
  tag_mem_pkt_v_o,
  tag_mem_pkt_o,
  tag_mem_pkt_yumi_i,
  stat_mem_pkt_v_o,
  stat_mem_pkt_o,
  lru_way_i,
  dirty_i,
  stat_mem_pkt_yumi_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i
);

  input [0:0] lce_id_i;
  input [21:0] miss_addr_i;
  input [63:0] store_data_i;
  input [1:0] size_op_i;
  output [522:0] data_mem_pkt_o;
  input [511:0] data_mem_data_i;
  output [22:0] tag_mem_pkt_o;
  output [10:0] stat_mem_pkt_o;
  input [2:0] lru_way_i;
  input [7:0] dirty_i;
  output [96:0] lce_req_o;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  input [35:0] lce_cmd_i;
  input [517:0] lce_data_cmd_i;
  output [517:0] lce_data_cmd_o;
  input clk_i;
  input reset_i;
  input load_miss_i;
  input store_miss_i;
  input uncached_load_req_i;
  input uncached_store_req_i;
  input data_mem_pkt_yumi_i;
  input tag_mem_pkt_yumi_i;
  input stat_mem_pkt_yumi_i;
  input lce_req_ready_i;
  input lce_resp_ready_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_v_i;
  input lce_data_cmd_ready_i;
  output ready_o;
  output cache_miss_o;
  output data_mem_pkt_v_o;
  output tag_mem_pkt_v_o;
  output stat_mem_pkt_v_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_ready_o;
  output lce_data_cmd_ready_o;
  output lce_data_cmd_v_o;
  wire [522:0] data_mem_pkt_o,lce_cmd_data_mem_pkt_lo,lce_data_cmd_data_mem_pkt_lo;
  wire [22:0] tag_mem_pkt_o;
  wire [10:0] stat_mem_pkt_o;
  wire [96:0] lce_req_o;
  wire [25:0] lce_resp_o,lce_req_to_lce_resp_lo,lce_cmd_to_lce_resp_lo;
  wire [536:0] lce_data_resp_o;
  wire [517:0] lce_data_cmd_o;
  wire ready_o,cache_miss_o,data_mem_pkt_v_o,tag_mem_pkt_v_o,stat_mem_pkt_v_o,
  lce_req_v_o,lce_resp_v_o,lce_data_resp_v_o,lce_cmd_ready_o,lce_data_cmd_ready_o,
  lce_data_cmd_v_o,N0,N1,N2,N3,N4,N5,N6,tr_data_received,cce_data_received,
  uncached_data_received,set_tag_received,set_tag_wakeup_received,lce_req_to_lce_resp_v_lo,
  lce_req_to_lce_resp_yumi_li,lce_sync_done_lo,lce_cmd_to_lce_resp_v_lo,
  lce_cmd_to_lce_resp_yumi_li,lce_cmd_data_mem_pkt_v_lo,lce_cmd_data_mem_pkt_yumi_li,
  lce_data_cmd_data_mem_pkt_v_lo,lce_data_cmd_data_mem_pkt_yumi_li,N7,N8,N9,N10,timeout,N11,N12,
  N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,
  N33,N34,N35,N36,N37;
  wire [21:0] miss_addr_lo;
  wire [2:0] timeout_count_n;
  reg [2:0] timeout_count_r;

  bp_be_dcache_lce_req_data_width_p64_paddr_width_p22_num_cce_p1_num_lce_p2_ways_p8
  lce_req_inst
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .lce_id_i(lce_id_i[0]),
    .load_miss_i(load_miss_i),
    .store_miss_i(store_miss_i),
    .miss_addr_i(miss_addr_i),
    .lru_way_i(lru_way_i),
    .dirty_i(dirty_i),
    .uncached_load_req_i(uncached_load_req_i),
    .uncached_store_req_i(uncached_store_req_i),
    .store_data_i(store_data_i),
    .size_op_i(size_op_i),
    .cache_miss_o(cache_miss_o),
    .miss_addr_o(miss_addr_lo),
    .tr_data_received_i(tr_data_received),
    .cce_data_received_i(cce_data_received),
    .uncached_data_received_i(uncached_data_received),
    .set_tag_received_i(set_tag_received),
    .set_tag_wakeup_received_i(set_tag_wakeup_received),
    .lce_req_o(lce_req_o),
    .lce_req_v_o(lce_req_v_o),
    .lce_req_ready_i(lce_req_ready_i),
    .lce_resp_o(lce_req_to_lce_resp_lo),
    .lce_resp_v_o(lce_req_to_lce_resp_v_lo),
    .lce_resp_yumi_i(lce_req_to_lce_resp_yumi_li)
  );


  bp_be_dcache_lce_cmd_num_cce_p1_num_lce_p2_paddr_width_p22_lce_data_width_p512_sets_p64_ways_p8_data_width_p64
  lce_cmd_inst
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .lce_id_i(lce_id_i[0]),
    .lce_sync_done_o(lce_sync_done_lo),
    .set_tag_received_o(set_tag_received),
    .set_tag_wakeup_received_o(set_tag_wakeup_received),
    .lce_cmd_i(lce_cmd_i),
    .lce_cmd_v_i(lce_cmd_v_i),
    .lce_cmd_yumi_o(lce_cmd_ready_o),
    .lce_resp_o(lce_cmd_to_lce_resp_lo),
    .lce_resp_v_o(lce_cmd_to_lce_resp_v_lo),
    .lce_resp_yumi_i(lce_cmd_to_lce_resp_yumi_li),
    .lce_data_resp_o(lce_data_resp_o),
    .lce_data_resp_v_o(lce_data_resp_v_o),
    .lce_data_resp_ready_i(lce_data_resp_ready_i),
    .lce_data_cmd_o(lce_data_cmd_o),
    .lce_data_cmd_v_o(lce_data_cmd_v_o),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_i),
    .data_mem_pkt_v_o(lce_cmd_data_mem_pkt_v_lo),
    .data_mem_pkt_o(lce_cmd_data_mem_pkt_lo),
    .data_mem_data_i(data_mem_data_i),
    .data_mem_pkt_yumi_i(lce_cmd_data_mem_pkt_yumi_li),
    .tag_mem_pkt_v_o(tag_mem_pkt_v_o),
    .tag_mem_pkt_o(tag_mem_pkt_o),
    .tag_mem_pkt_yumi_i(tag_mem_pkt_yumi_i),
    .stat_mem_pkt_v_o(stat_mem_pkt_v_o),
    .stat_mem_pkt_o(stat_mem_pkt_o),
    .dirty_i(dirty_i),
    .stat_mem_pkt_yumi_i(stat_mem_pkt_yumi_i)
  );


  bp_be_dcache_lce_data_cmd_num_cce_p1_num_lce_p2_data_width_p64_paddr_width_p22_lce_data_width_p512_ways_p8_sets_p64
  lce_data_cmd_inst
  (
    .cce_data_received_o(cce_data_received),
    .tr_data_received_o(tr_data_received),
    .uncached_data_received_o(uncached_data_received),
    .miss_addr_i(miss_addr_lo),
    .lce_data_cmd_i(lce_data_cmd_i),
    .lce_data_cmd_v_i(lce_data_cmd_v_i),
    .lce_data_cmd_yumi_o(lce_data_cmd_ready_o),
    .data_mem_pkt_v_o(lce_data_cmd_data_mem_pkt_v_lo),
    .data_mem_pkt_o(lce_data_cmd_data_mem_pkt_lo),
    .data_mem_pkt_yumi_i(lce_data_cmd_data_mem_pkt_yumi_li)
  );

  assign N26 = ~timeout_count_r[2];
  assign N27 = timeout_count_r[1] | N26;
  assign N28 = timeout_count_r[0] | N27;
  assign N29 = ~N28;
  assign { N19, N18, N17 } = timeout_count_r + 1'b1;
  assign data_mem_pkt_v_o = (N0)? 1'b1 :
                            (N1)? lce_cmd_data_mem_pkt_v_lo : 1'b0;
  assign N0 = lce_data_cmd_data_mem_pkt_v_lo;
  assign N1 = N7;
  assign data_mem_pkt_o = (N0)? lce_data_cmd_data_mem_pkt_lo :
                          (N1)? lce_cmd_data_mem_pkt_lo : 1'b0;
  assign lce_data_cmd_data_mem_pkt_yumi_li = (N0)? data_mem_pkt_yumi_i :
                                             (N1)? 1'b0 : 1'b0;
  assign lce_cmd_data_mem_pkt_yumi_li = (N0)? 1'b0 :
                                        (N1)? data_mem_pkt_yumi_i : 1'b0;
  assign lce_resp_v_o = (N2)? 1'b1 :
                        (N3)? lce_cmd_to_lce_resp_v_lo : 1'b0;
  assign N2 = lce_req_to_lce_resp_v_lo;
  assign N3 = N8;
  assign lce_resp_o = (N2)? lce_req_to_lce_resp_lo :
                      (N3)? lce_cmd_to_lce_resp_lo : 1'b0;
  assign lce_req_to_lce_resp_yumi_li = (N2)? lce_resp_ready_i :
                                       (N3)? 1'b0 : 1'b0;
  assign lce_cmd_to_lce_resp_yumi_li = (N2)? 1'b0 :
                                       (N3)? N9 : 1'b0;
  assign { N22, N21, N20 } = (N4)? { N19, N18, N17 } :
                             (N16)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N4 = N15;
  assign { N25, N24, N23 } = (N5)? { N22, N21, N20 } :
                             (N13)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N5 = N12;
  assign timeout_count_n = (N6)? { 1'b0, 1'b0, 1'b0 } :
                           (N10)? { N25, N24, N23 } : 1'b0;
  assign N6 = timeout;
  assign N7 = ~lce_data_cmd_data_mem_pkt_v_lo;
  assign N8 = ~lce_req_to_lce_resp_v_lo;
  assign N9 = lce_cmd_to_lce_resp_v_lo & lce_resp_ready_i;
  assign timeout = N29;
  assign N10 = ~timeout;
  assign N11 = N10;
  assign N12 = N30 | stat_mem_pkt_v_o;
  assign N30 = data_mem_pkt_v_o | tag_mem_pkt_v_o;
  assign N13 = ~N12;
  assign N14 = N11 & N12;
  assign N15 = N33 & N34;
  assign N33 = N31 & N32;
  assign N31 = ~data_mem_pkt_yumi_i;
  assign N32 = ~tag_mem_pkt_yumi_i;
  assign N34 = ~stat_mem_pkt_yumi_i;
  assign N16 = ~N15;
  assign ready_o = N36 & N37;
  assign N36 = lce_sync_done_lo & N35;
  assign N35 = ~timeout;
  assign N37 = ~cache_miss_o;

  always @(posedge clk_i) begin
    if(reset_i) begin
      { timeout_count_r[2:0] } <= { 1'b0, 1'b0, 1'b0 };
    end else if(1'b1) begin
      { timeout_count_r[2:0] } <= { timeout_count_n[2:0] };
    end
  end


endmodule



module bsg_mux_width_p32_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [63:0] data_i;
  input [0:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1;
  assign data_o[31] = (N1)? data_i[31] :
                      (N0)? data_i[63] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[30] = (N1)? data_i[30] :
                      (N0)? data_i[62] : 1'b0;
  assign data_o[29] = (N1)? data_i[29] :
                      (N0)? data_i[61] : 1'b0;
  assign data_o[28] = (N1)? data_i[28] :
                      (N0)? data_i[60] : 1'b0;
  assign data_o[27] = (N1)? data_i[27] :
                      (N0)? data_i[59] : 1'b0;
  assign data_o[26] = (N1)? data_i[26] :
                      (N0)? data_i[58] : 1'b0;
  assign data_o[25] = (N1)? data_i[25] :
                      (N0)? data_i[57] : 1'b0;
  assign data_o[24] = (N1)? data_i[24] :
                      (N0)? data_i[56] : 1'b0;
  assign data_o[23] = (N1)? data_i[23] :
                      (N0)? data_i[55] : 1'b0;
  assign data_o[22] = (N1)? data_i[22] :
                      (N0)? data_i[54] : 1'b0;
  assign data_o[21] = (N1)? data_i[21] :
                      (N0)? data_i[53] : 1'b0;
  assign data_o[20] = (N1)? data_i[20] :
                      (N0)? data_i[52] : 1'b0;
  assign data_o[19] = (N1)? data_i[19] :
                      (N0)? data_i[51] : 1'b0;
  assign data_o[18] = (N1)? data_i[18] :
                      (N0)? data_i[50] : 1'b0;
  assign data_o[17] = (N1)? data_i[17] :
                      (N0)? data_i[49] : 1'b0;
  assign data_o[16] = (N1)? data_i[16] :
                      (N0)? data_i[48] : 1'b0;
  assign data_o[15] = (N1)? data_i[15] :
                      (N0)? data_i[47] : 1'b0;
  assign data_o[14] = (N1)? data_i[14] :
                      (N0)? data_i[46] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] :
                      (N0)? data_i[45] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] :
                      (N0)? data_i[44] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] :
                      (N0)? data_i[43] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] :
                      (N0)? data_i[42] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] :
                     (N0)? data_i[41] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] :
                     (N0)? data_i[40] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] :
                     (N0)? data_i[39] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] :
                     (N0)? data_i[38] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] :
                     (N0)? data_i[37] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] :
                     (N0)? data_i[36] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] :
                     (N0)? data_i[35] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] :
                     (N0)? data_i[34] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] :
                     (N0)? data_i[33] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] :
                     (N0)? data_i[32] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_mux_width_p16_els_p4
(
  data_i,
  sel_i,
  data_o
);

  input [63:0] data_i;
  input [1:0] sel_i;
  output [15:0] data_o;
  wire [15:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[15] = (N2)? data_i[15] :
                      (N4)? data_i[31] :
                      (N3)? data_i[47] :
                      (N5)? data_i[63] : 1'b0;
  assign data_o[14] = (N2)? data_i[14] :
                      (N4)? data_i[30] :
                      (N3)? data_i[46] :
                      (N5)? data_i[62] : 1'b0;
  assign data_o[13] = (N2)? data_i[13] :
                      (N4)? data_i[29] :
                      (N3)? data_i[45] :
                      (N5)? data_i[61] : 1'b0;
  assign data_o[12] = (N2)? data_i[12] :
                      (N4)? data_i[28] :
                      (N3)? data_i[44] :
                      (N5)? data_i[60] : 1'b0;
  assign data_o[11] = (N2)? data_i[11] :
                      (N4)? data_i[27] :
                      (N3)? data_i[43] :
                      (N5)? data_i[59] : 1'b0;
  assign data_o[10] = (N2)? data_i[10] :
                      (N4)? data_i[26] :
                      (N3)? data_i[42] :
                      (N5)? data_i[58] : 1'b0;
  assign data_o[9] = (N2)? data_i[9] :
                     (N4)? data_i[25] :
                     (N3)? data_i[41] :
                     (N5)? data_i[57] : 1'b0;
  assign data_o[8] = (N2)? data_i[8] :
                     (N4)? data_i[24] :
                     (N3)? data_i[40] :
                     (N5)? data_i[56] : 1'b0;
  assign data_o[7] = (N2)? data_i[7] :
                     (N4)? data_i[23] :
                     (N3)? data_i[39] :
                     (N5)? data_i[55] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] :
                     (N4)? data_i[22] :
                     (N3)? data_i[38] :
                     (N5)? data_i[54] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] :
                     (N4)? data_i[21] :
                     (N3)? data_i[37] :
                     (N5)? data_i[53] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] :
                     (N4)? data_i[20] :
                     (N3)? data_i[36] :
                     (N5)? data_i[52] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] :
                     (N4)? data_i[19] :
                     (N3)? data_i[35] :
                     (N5)? data_i[51] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] :
                     (N4)? data_i[18] :
                     (N3)? data_i[34] :
                     (N5)? data_i[50] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] :
                     (N4)? data_i[17] :
                     (N3)? data_i[33] :
                     (N5)? data_i[49] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] :
                     (N4)? data_i[16] :
                     (N3)? data_i[32] :
                     (N5)? data_i[48] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_mux_width_p8_els_p8
(
  data_i,
  sel_i,
  data_o
);

  input [63:0] data_i;
  input [2:0] sel_i;
  output [7:0] data_o;
  wire [7:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14;
  assign data_o[7] = (N7)? data_i[7] :
                     (N9)? data_i[15] :
                     (N11)? data_i[23] :
                     (N13)? data_i[31] :
                     (N8)? data_i[39] :
                     (N10)? data_i[47] :
                     (N12)? data_i[55] :
                     (N14)? data_i[63] : 1'b0;
  assign data_o[6] = (N7)? data_i[6] :
                     (N9)? data_i[14] :
                     (N11)? data_i[22] :
                     (N13)? data_i[30] :
                     (N8)? data_i[38] :
                     (N10)? data_i[46] :
                     (N12)? data_i[54] :
                     (N14)? data_i[62] : 1'b0;
  assign data_o[5] = (N7)? data_i[5] :
                     (N9)? data_i[13] :
                     (N11)? data_i[21] :
                     (N13)? data_i[29] :
                     (N8)? data_i[37] :
                     (N10)? data_i[45] :
                     (N12)? data_i[53] :
                     (N14)? data_i[61] : 1'b0;
  assign data_o[4] = (N7)? data_i[4] :
                     (N9)? data_i[12] :
                     (N11)? data_i[20] :
                     (N13)? data_i[28] :
                     (N8)? data_i[36] :
                     (N10)? data_i[44] :
                     (N12)? data_i[52] :
                     (N14)? data_i[60] : 1'b0;
  assign data_o[3] = (N7)? data_i[3] :
                     (N9)? data_i[11] :
                     (N11)? data_i[19] :
                     (N13)? data_i[27] :
                     (N8)? data_i[35] :
                     (N10)? data_i[43] :
                     (N12)? data_i[51] :
                     (N14)? data_i[59] : 1'b0;
  assign data_o[2] = (N7)? data_i[2] :
                     (N9)? data_i[10] :
                     (N11)? data_i[18] :
                     (N13)? data_i[26] :
                     (N8)? data_i[34] :
                     (N10)? data_i[42] :
                     (N12)? data_i[50] :
                     (N14)? data_i[58] : 1'b0;
  assign data_o[1] = (N7)? data_i[1] :
                     (N9)? data_i[9] :
                     (N11)? data_i[17] :
                     (N13)? data_i[25] :
                     (N8)? data_i[33] :
                     (N10)? data_i[41] :
                     (N12)? data_i[49] :
                     (N14)? data_i[57] : 1'b0;
  assign data_o[0] = (N7)? data_i[0] :
                     (N9)? data_i[8] :
                     (N11)? data_i[16] :
                     (N13)? data_i[24] :
                     (N8)? data_i[32] :
                     (N10)? data_i[40] :
                     (N12)? data_i[48] :
                     (N14)? data_i[56] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];
  assign N6 = ~sel_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & sel_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & sel_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & sel_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & sel_i[2];

endmodule



module bsg_decode_with_v_num_out_p8
(
  i,
  v_i,
  o
);

  input [2:0] i;
  output [7:0] o;
  input v_i;
  wire [7:0] o,lo;

  bsg_decode_num_out_p8
  bd
  (
    .i(i),
    .o(lo)
  );

  assign o[7] = v_i & lo[7];
  assign o[6] = v_i & lo[6];
  assign o[5] = v_i & lo[5];
  assign o[4] = v_i & lo[4];
  assign o[3] = v_i & lo[3];
  assign o[2] = v_i & lo[2];
  assign o[1] = v_i & lo[1];
  assign o[0] = v_i & lo[0];

endmodule



module bp_be_dcache_data_width_p64_paddr_width_p22_sets_p64_ways_p8_num_cce_p1_num_lce_p2
(
  clk_i,
  reset_i,
  lce_id_i,
  dcache_pkt_i,
  v_i,
  ready_o,
  data_o,
  v_o,
  tlb_miss_i,
  ptag_i,
  uncached_i,
  cache_miss_o,
  poison_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i
);

  input [0:0] lce_id_i;
  input [79:0] dcache_pkt_i;
  output [63:0] data_o;
  input [9:0] ptag_i;
  output [96:0] lce_req_o;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  input [35:0] lce_cmd_i;
  input [517:0] lce_data_cmd_i;
  output [517:0] lce_data_cmd_o;
  input clk_i;
  input reset_i;
  input v_i;
  input tlb_miss_i;
  input uncached_i;
  input poison_i;
  input lce_req_ready_i;
  input lce_resp_ready_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_v_i;
  input lce_data_cmd_ready_i;
  output ready_o;
  output v_o;
  output cache_miss_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_ready_o;
  output lce_data_cmd_ready_o;
  output lce_data_cmd_v_o;
  wire [63:0] data_o,data_mem_mask_li,bypass_data_lo,ld_data_way_picked,bypass_data_masked;
  wire [96:0] lce_req_o,wbuf_entry_out;
  wire [25:0] lce_resp_o;
  wire [536:0] lce_data_resp_o;
  wire [517:0] lce_data_cmd_o;
  wire ready_o,v_o,cache_miss_o,lce_req_v_o,lce_resp_v_o,lce_data_resp_v_o,
  lce_cmd_ready_o,lce_data_cmd_ready_o,lce_data_cmd_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,
  N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,
  N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,
  N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,load_op,
  signed_op,tl_we,N70,N71,N72,N73,N74,N75,n_0_net_,tag_mem_w_li,tag_mem_v_li,
  n_1_net_,data_mem_w_li,n_2_net_,n_3_net_,n_4_net_,n_5_net_,n_6_net_,n_7_net_,
  n_8_net_,tv_we,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,load_hit,
  store_hit,load_miss_tv,store_miss_tv,uncached_load_req,uncached_store_req,wbuf_v_li,
  wbuf_entry_in_data__63_,wbuf_entry_in_data__62_,wbuf_entry_in_data__61_,
  wbuf_entry_in_data__60_,wbuf_entry_in_data__59_,wbuf_entry_in_data__58_,
  wbuf_entry_in_data__57_,wbuf_entry_in_data__56_,wbuf_entry_in_data__55_,wbuf_entry_in_data__54_,
  wbuf_entry_in_data__53_,wbuf_entry_in_data__52_,wbuf_entry_in_data__51_,
  wbuf_entry_in_data__50_,wbuf_entry_in_data__49_,wbuf_entry_in_data__48_,
  wbuf_entry_in_data__47_,wbuf_entry_in_data__46_,wbuf_entry_in_data__45_,wbuf_entry_in_data__44_,
  wbuf_entry_in_data__43_,wbuf_entry_in_data__42_,wbuf_entry_in_data__41_,
  wbuf_entry_in_data__40_,wbuf_entry_in_data__39_,wbuf_entry_in_data__38_,
  wbuf_entry_in_data__37_,wbuf_entry_in_data__36_,wbuf_entry_in_data__35_,wbuf_entry_in_data__34_,
  wbuf_entry_in_data__33_,wbuf_entry_in_data__32_,wbuf_entry_in_data__31_,
  wbuf_entry_in_data__30_,wbuf_entry_in_data__29_,wbuf_entry_in_data__28_,
  wbuf_entry_in_data__27_,wbuf_entry_in_data__26_,wbuf_entry_in_data__25_,wbuf_entry_in_data__24_,
  wbuf_entry_in_data__23_,wbuf_entry_in_data__22_,wbuf_entry_in_data__21_,
  wbuf_entry_in_data__20_,wbuf_entry_in_data__19_,wbuf_entry_in_data__18_,
  wbuf_entry_in_data__17_,wbuf_entry_in_data__16_,wbuf_entry_in_data__15_,wbuf_entry_in_data__14_,
  wbuf_entry_in_data__13_,wbuf_entry_in_data__12_,wbuf_entry_in_data__11_,
  wbuf_entry_in_data__10_,wbuf_entry_in_data__9_,wbuf_entry_in_data__8_,
  wbuf_entry_in_mask__7_,wbuf_entry_in_mask__6_,wbuf_entry_in_mask__5_,wbuf_entry_in_mask__4_,
  wbuf_entry_in_mask__3_,wbuf_entry_in_mask__2_,wbuf_entry_in_mask__1_,
  wbuf_entry_in_mask__0_,wbuf_v_lo,wbuf_yumi_li,wbuf_empty_lo,bypass_v_li,lce_snoop_match_lo,N90,N91,
  N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,
  N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,n_10_net_,
  stat_mem_w_li,stat_mem_v_li,invalid_exist,N124,lce_data_mem_pkt_v,
  lce_data_mem_pkt_yumi,lce_tag_mem_pkt_v,lce_tag_mem_pkt_yumi,lce_stat_mem_pkt_v,
  lce_stat_mem_pkt_yumi,N125,N126,N127,N128,N129,N130,N131,N132,N133,n_13_net__2_,n_13_net__1_,
  n_13_net__0_,genblk4_word_sigext,genblk4_half_sigext,genblk4_byte_sigext,N134,
  N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,
  N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,
  N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,
  N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,
  N199,N200,N201,N202,N203,N204,N205,N206,N207,n_14_net__2_,n_14_net__1_,
  n_14_net__0_,lce_data_mem_v,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,
  N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,
  N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,
  N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,
  N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,
  N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,
  N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,
  dirty_mask_v_li,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,
  N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,
  N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,
  N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,
  N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,
  N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
  N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,
  N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,
  N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,
  N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,
  N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488;
  wire [5:0] tag_mem_addr_li,stat_mem_addr_li;
  wire [95:0] tag_mem_data_li,tag_mem_mask_li,tag_mem_data_lo;
  wire [71:0] data_mem_addr_li;
  wire [511:0] data_mem_data_li,data_mem_data_lo,lce_data_mem_data_li,lce_data_mem_write_data;
  wire [7:0] data_mem_v_li,tag_match_tv,load_hit_tv,store_hit_tv,bypass_mask_lo,
  genblk4_data_byte_selected,wbuf_data_mem_v,lce_tag_mem_way_one_hot,dirty_mask_lo;
  wire [2:0] load_hit_way,store_hit_way,lru_encode,invalid_way,lce_lru_way_li,
  lru_decode_way_li,dirty_mask_way_li;
  wire [14:0] stat_mem_data_li,stat_mem_mask_li,stat_mem_data_lo;
  wire [522:0] lce_data_mem_pkt;
  wire [22:0] lce_tag_mem_pkt;
  wire [10:0] lce_stat_mem_pkt;
  wire [31:0] genblk4_data_word_selected;
  wire [15:0] genblk4_data_half_selected;
  wire [6:0] lru_decode_data_lo,lru_decode_mask_lo;
  reg [63:0] data_tl_r,data_tv_r,uncached_load_data_r;
  reg v_tl_r,load_op_tl_r,store_op_tl_r,signed_op_tl_r,double_op_tl_r,word_op_tl_r,
  half_op_tl_r,v_tv_r,uncached_tv_r,load_op_tv_r,store_op_tv_r,signed_op_tv_r,
  double_op_tv_r,word_op_tv_r,half_op_tv_r,uncached_load_data_v_r;
  reg [11:0] page_offset_tl_r;
  reg [1:0] size_op_tl_r,size_op_tv_r;
  reg [21:0] paddr_tv_r;
  reg [95:0] tag_info_tv_r;
  reg [511:0] ld_data_tv_r;
  reg [2:0] lce_data_mem_pkt_way_r;

  bsg_mem_1rw_sync_mask_write_bit_width_p96_els_p64
  tag_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(tag_mem_data_li),
    .addr_i(tag_mem_addr_li),
    .v_i(n_0_net_),
    .w_mask_i(tag_mem_mask_li),
    .w_i(tag_mem_w_li),
    .data_o(tag_mem_data_lo)
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_0__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_1_net_),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li[8:0]),
    .data_i(data_mem_data_li[63:0]),
    .write_mask_i(data_mem_mask_li[7:0]),
    .data_o(data_mem_data_lo[63:0])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_1__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_2_net_),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li[17:9]),
    .data_i(data_mem_data_li[127:64]),
    .write_mask_i(data_mem_mask_li[15:8]),
    .data_o(data_mem_data_lo[127:64])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_2__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_3_net_),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li[26:18]),
    .data_i(data_mem_data_li[191:128]),
    .write_mask_i(data_mem_mask_li[23:16]),
    .data_o(data_mem_data_lo[191:128])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_3__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_4_net_),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li[35:27]),
    .data_i(data_mem_data_li[255:192]),
    .write_mask_i(data_mem_mask_li[31:24]),
    .data_o(data_mem_data_lo[255:192])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_4__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_5_net_),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li[44:36]),
    .data_i(data_mem_data_li[319:256]),
    .write_mask_i(data_mem_mask_li[39:32]),
    .data_o(data_mem_data_lo[319:256])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_5__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_6_net_),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li[53:45]),
    .data_i(data_mem_data_li[383:320]),
    .write_mask_i(data_mem_mask_li[47:40]),
    .data_o(data_mem_data_lo[383:320])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_6__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_7_net_),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li[62:54]),
    .data_i(data_mem_data_li[447:384]),
    .write_mask_i(data_mem_mask_li[55:48]),
    .data_o(data_mem_data_lo[447:384])
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p512_data_width_p64
  data_mem_7__data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(n_8_net_),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li[71:63]),
    .data_i(data_mem_data_li[511:448]),
    .write_mask_i(data_mem_mask_li[63:56]),
    .data_o(data_mem_data_lo[511:448])
  );

  assign tag_match_tv[0] = paddr_tv_r[21:12] == tag_info_tv_r[9:0];
  assign tag_match_tv[1] = paddr_tv_r[21:12] == tag_info_tv_r[21:12];
  assign tag_match_tv[2] = paddr_tv_r[21:12] == tag_info_tv_r[33:24];
  assign tag_match_tv[3] = paddr_tv_r[21:12] == tag_info_tv_r[45:36];
  assign tag_match_tv[4] = paddr_tv_r[21:12] == tag_info_tv_r[57:48];
  assign tag_match_tv[5] = paddr_tv_r[21:12] == tag_info_tv_r[69:60];
  assign tag_match_tv[6] = paddr_tv_r[21:12] == tag_info_tv_r[81:72];
  assign tag_match_tv[7] = paddr_tv_r[21:12] == tag_info_tv_r[93:84];

  bsg_priority_encode_width_p8_lo_to_hi_p1
  pe_load_hit
  (
    .i(load_hit_tv),
    .addr_o(load_hit_way),
    .v_o(load_hit)
  );


  bsg_priority_encode_width_p8_lo_to_hi_p1
  pe_store_hit
  (
    .i(store_hit_tv),
    .addr_o(store_hit_way),
    .v_o(store_hit)
  );


  bp_be_dcache_wbuf_data_width_p64_paddr_width_p22_ways_p8_sets_p64
  wbuf
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(wbuf_v_li),
    .wbuf_entry_i({ paddr_tv_r, wbuf_entry_in_data__63_, wbuf_entry_in_data__62_, wbuf_entry_in_data__61_, wbuf_entry_in_data__60_, wbuf_entry_in_data__59_, wbuf_entry_in_data__58_, wbuf_entry_in_data__57_, wbuf_entry_in_data__56_, wbuf_entry_in_data__55_, wbuf_entry_in_data__54_, wbuf_entry_in_data__53_, wbuf_entry_in_data__52_, wbuf_entry_in_data__51_, wbuf_entry_in_data__50_, wbuf_entry_in_data__49_, wbuf_entry_in_data__48_, wbuf_entry_in_data__47_, wbuf_entry_in_data__46_, wbuf_entry_in_data__45_, wbuf_entry_in_data__44_, wbuf_entry_in_data__43_, wbuf_entry_in_data__42_, wbuf_entry_in_data__41_, wbuf_entry_in_data__40_, wbuf_entry_in_data__39_, wbuf_entry_in_data__38_, wbuf_entry_in_data__37_, wbuf_entry_in_data__36_, wbuf_entry_in_data__35_, wbuf_entry_in_data__34_, wbuf_entry_in_data__33_, wbuf_entry_in_data__32_, wbuf_entry_in_data__31_, wbuf_entry_in_data__30_, wbuf_entry_in_data__29_, wbuf_entry_in_data__28_, wbuf_entry_in_data__27_, wbuf_entry_in_data__26_, wbuf_entry_in_data__25_, wbuf_entry_in_data__24_, wbuf_entry_in_data__23_, wbuf_entry_in_data__22_, wbuf_entry_in_data__21_, wbuf_entry_in_data__20_, wbuf_entry_in_data__19_, wbuf_entry_in_data__18_, wbuf_entry_in_data__17_, wbuf_entry_in_data__16_, wbuf_entry_in_data__15_, wbuf_entry_in_data__14_, wbuf_entry_in_data__13_, wbuf_entry_in_data__12_, wbuf_entry_in_data__11_, wbuf_entry_in_data__10_, wbuf_entry_in_data__9_, wbuf_entry_in_data__8_, data_tv_r[7:0], wbuf_entry_in_mask__7_, wbuf_entry_in_mask__6_, wbuf_entry_in_mask__5_, wbuf_entry_in_mask__4_, wbuf_entry_in_mask__3_, wbuf_entry_in_mask__2_, wbuf_entry_in_mask__1_, wbuf_entry_in_mask__0_, store_hit_way }),
    .yumi_i(wbuf_yumi_li),
    .v_o(wbuf_v_lo),
    .wbuf_entry_o(wbuf_entry_out),
    .empty_o(wbuf_empty_lo),
    .bypass_addr_i({ ptag_i, page_offset_tl_r }),
    .bypass_v_i(bypass_v_li),
    .bypass_data_o(bypass_data_lo),
    .bypass_mask_o(bypass_mask_lo),
    .lce_snoop_index_i(lce_data_mem_pkt[522:517]),
    .lce_snoop_way_i(lce_data_mem_pkt[516:514]),
    .lce_snoop_match_o(lce_snoop_match_lo)
  );


  bsg_mem_1rw_sync_mask_write_bit_width_p15_els_p64
  stat_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(stat_mem_data_li),
    .addr_i(stat_mem_addr_li),
    .v_i(n_10_net_),
    .w_mask_i(stat_mem_mask_li),
    .w_i(stat_mem_w_li),
    .data_o(stat_mem_data_lo)
  );


  bsg_lru_pseudo_tree_encode_ways_p8
  lru_encoder
  (
    .lru_i(stat_mem_data_lo[14:8]),
    .way_id_o(lru_encode)
  );


  bsg_priority_encode_width_p8_lo_to_hi_p1
  pe_invalid
  (
    .i({ N354, N356, N358, N360, N362, N364, N366, N368 }),
    .addr_o(invalid_way),
    .v_o(invalid_exist)
  );


  bp_be_dcache_lce_data_width_p64_paddr_width_p22_lce_data_width_p512_sets_p64_ways_p8_num_cce_p1_num_lce_p2
  lce
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .lce_id_i(lce_id_i[0]),
    .ready_o(ready_o),
    .cache_miss_o(cache_miss_o),
    .load_miss_i(load_miss_tv),
    .store_miss_i(store_miss_tv),
    .uncached_load_req_i(uncached_load_req),
    .uncached_store_req_i(uncached_store_req),
    .miss_addr_i(paddr_tv_r),
    .store_data_i(data_tv_r),
    .size_op_i(size_op_tv_r),
    .data_mem_pkt_v_o(lce_data_mem_pkt_v),
    .data_mem_pkt_o(lce_data_mem_pkt),
    .data_mem_data_i(lce_data_mem_data_li),
    .data_mem_pkt_yumi_i(lce_data_mem_pkt_yumi),
    .tag_mem_pkt_v_o(lce_tag_mem_pkt_v),
    .tag_mem_pkt_o(lce_tag_mem_pkt),
    .tag_mem_pkt_yumi_i(lce_tag_mem_pkt_yumi),
    .stat_mem_pkt_v_o(lce_stat_mem_pkt_v),
    .stat_mem_pkt_o(lce_stat_mem_pkt),
    .lru_way_i(lce_lru_way_li),
    .dirty_i(stat_mem_data_lo[7:0]),
    .stat_mem_pkt_yumi_i(lce_stat_mem_pkt_yumi),
    .lce_req_o(lce_req_o),
    .lce_req_v_o(lce_req_v_o),
    .lce_req_ready_i(lce_req_ready_i),
    .lce_resp_o(lce_resp_o),
    .lce_resp_v_o(lce_resp_v_o),
    .lce_resp_ready_i(lce_resp_ready_i),
    .lce_data_resp_o(lce_data_resp_o),
    .lce_data_resp_v_o(lce_data_resp_v_o),
    .lce_data_resp_ready_i(lce_data_resp_ready_i),
    .lce_cmd_i(lce_cmd_i),
    .lce_cmd_v_i(lce_cmd_v_i),
    .lce_cmd_ready_o(lce_cmd_ready_o),
    .lce_data_cmd_i(lce_data_cmd_i),
    .lce_data_cmd_v_i(lce_data_cmd_v_i),
    .lce_data_cmd_ready_o(lce_data_cmd_ready_o),
    .lce_data_cmd_o(lce_data_cmd_o),
    .lce_data_cmd_v_o(lce_data_cmd_v_o),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_i)
  );


  bsg_mux_width_p64_els_p8
  ld_data_set_select_mux
  (
    .data_i(ld_data_tv_r),
    .sel_i({ n_13_net__2_, n_13_net__1_, n_13_net__0_ }),
    .data_o(ld_data_way_picked)
  );


  bsg_mux_segmented_segments_p8_segment_width_p8
  bypass_mux_segmented
  (
    .data0_i(ld_data_way_picked),
    .data1_i(bypass_data_lo),
    .sel_i(bypass_mask_lo),
    .data_o(bypass_data_masked)
  );


  bsg_mux_width_p32_els_p2
  genblk4_word_mux
  (
    .data_i(bypass_data_masked),
    .sel_i(paddr_tv_r[2]),
    .data_o(genblk4_data_word_selected)
  );


  bsg_mux_width_p16_els_p4
  genblk4_half_mux
  (
    .data_i(bypass_data_masked),
    .sel_i(paddr_tv_r[2:1]),
    .data_o(genblk4_data_half_selected)
  );


  bsg_mux_width_p8_els_p8
  genblk4_byte_mux
  (
    .data_i(bypass_data_masked),
    .sel_i(paddr_tv_r[2:0]),
    .data_o(genblk4_data_byte_selected)
  );


  bsg_decode_num_out_p8
  wbuf_data_mem_v_decode
  (
    .i({ n_14_net__2_, n_14_net__1_, n_14_net__0_ }),
    .o(wbuf_data_mem_v)
  );


  bsg_mux_butterfly_width_p64_els_p8
  write_mux_butterfly
  (
    .data_i(lce_data_mem_pkt[513:2]),
    .sel_i(lce_data_mem_pkt[516:514]),
    .data_o(lce_data_mem_write_data)
  );


  bsg_decode_num_out_p8
  lce_tag_mem_way_decode
  (
    .i(lce_tag_mem_pkt[16:14]),
    .o(lce_tag_mem_way_one_hot)
  );

  assign N308 = N306 & N307;
  assign N309 = lce_tag_mem_pkt[1] | N307;
  assign N311 = N306 | lce_tag_mem_pkt[0];
  assign N313 = lce_tag_mem_pkt[1] & lce_tag_mem_pkt[0];

  bsg_lru_pseudo_tree_decode_ways_p8
  lru_decode
  (
    .way_id_i(lru_decode_way_li),
    .data_o(lru_decode_data_lo),
    .mask_o(lru_decode_mask_lo)
  );


  bsg_decode_with_v_num_out_p8
  dirty_mask_decode
  (
    .i(dirty_mask_way_li),
    .v_i(dirty_mask_v_li),
    .o(dirty_mask_lo)
  );


  bsg_mux_butterfly_width_p64_els_p8
  read_mux_butterfly
  (
    .data_i(data_mem_data_lo),
    .sel_i(lce_data_mem_pkt_way_r),
    .data_o(lce_data_mem_data_li)
  );

  assign N353 = tag_info_tv_r[94] | tag_info_tv_r[95];
  assign N354 = ~N353;
  assign N355 = tag_info_tv_r[82] | tag_info_tv_r[83];
  assign N356 = ~N355;
  assign N357 = tag_info_tv_r[70] | tag_info_tv_r[71];
  assign N358 = ~N357;
  assign N359 = tag_info_tv_r[58] | tag_info_tv_r[59];
  assign N360 = ~N359;
  assign N361 = tag_info_tv_r[46] | tag_info_tv_r[47];
  assign N362 = ~N361;
  assign N363 = tag_info_tv_r[34] | tag_info_tv_r[35];
  assign N364 = ~N363;
  assign N365 = tag_info_tv_r[22] | tag_info_tv_r[23];
  assign N366 = ~N365;
  assign N367 = tag_info_tv_r[10] | tag_info_tv_r[11];
  assign N368 = ~N367;
  assign N369 = lce_data_mem_pkt[0] | lce_data_mem_pkt[1];
  assign N370 = ~N369;
  assign N371 = tag_info_tv_r[94] | tag_info_tv_r[95];
  assign N372 = tag_info_tv_r[82] | tag_info_tv_r[83];
  assign N373 = tag_info_tv_r[70] | tag_info_tv_r[71];
  assign N374 = tag_info_tv_r[58] | tag_info_tv_r[59];
  assign N375 = tag_info_tv_r[46] | tag_info_tv_r[47];
  assign N376 = tag_info_tv_r[34] | tag_info_tv_r[35];
  assign N377 = tag_info_tv_r[22] | tag_info_tv_r[23];
  assign N378 = tag_info_tv_r[10] | tag_info_tv_r[11];
  assign N379 = ~tag_info_tv_r[95];
  assign N380 = tag_info_tv_r[94] | N379;
  assign N381 = ~N380;
  assign N382 = ~tag_info_tv_r[83];
  assign N383 = tag_info_tv_r[82] | N382;
  assign N384 = ~N383;
  assign N385 = ~tag_info_tv_r[71];
  assign N386 = tag_info_tv_r[70] | N385;
  assign N387 = ~N386;
  assign N388 = ~tag_info_tv_r[59];
  assign N389 = tag_info_tv_r[58] | N388;
  assign N390 = ~N389;
  assign N391 = ~tag_info_tv_r[47];
  assign N392 = tag_info_tv_r[46] | N391;
  assign N393 = ~N392;
  assign N394 = ~tag_info_tv_r[35];
  assign N395 = tag_info_tv_r[34] | N394;
  assign N396 = ~N395;
  assign N397 = ~tag_info_tv_r[23];
  assign N398 = tag_info_tv_r[22] | N397;
  assign N399 = ~N398;
  assign N400 = ~tag_info_tv_r[11];
  assign N401 = tag_info_tv_r[10] | N400;
  assign N402 = ~N401;
  assign N403 = ~lce_stat_mem_pkt[0];
  assign N404 = N403 | lce_stat_mem_pkt[1];
  assign N405 = ~lce_data_mem_pkt[1];
  assign N406 = lce_data_mem_pkt[0] | N405;
  assign N407 = dcache_pkt_i[76] & dcache_pkt_i[77];
  assign N408 = ~dcache_pkt_i[77];
  assign N409 = dcache_pkt_i[76] | N408;
  assign N410 = ~N409;
  assign N411 = ~dcache_pkt_i[76];
  assign N412 = N411 | dcache_pkt_i[77];
  assign N413 = ~N412;
  assign N414 = ~lce_data_mem_pkt[0];
  assign N415 = N414 | lce_data_mem_pkt[1];
  assign N416 = ~N415;
  assign N417 = lce_data_mem_pkt[0] | N405;
  assign N418 = ~N417;
  assign N419 = lce_data_mem_pkt[0] | N405;
  assign N420 = ~N419;
  assign N73 = (N0)? 1'b0 :
               (N1)? tl_we : 1'b0;
  assign N0 = N71;
  assign N1 = N70;
  assign N74 = (N0)? 1'b0 :
               (N1)? tl_we : 1'b0;
  assign N75 = (N0)? 1'b0 :
               (N1)? N72 : 1'b0;
  assign N80 = (N2)? 1'b0 :
               (N3)? tv_we : 1'b0;
  assign N2 = N77;
  assign N3 = N76;
  assign N81 = (N2)? 1'b0 :
               (N3)? tv_we : 1'b0;
  assign N82 = (N2)? 1'b0 :
               (N3)? tv_we : 1'b0;
  assign { N88, N87, N86, N85, N84, N83 } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                            (N3)? { N78, N78, N78, N78, N78, N78 } : 1'b0;
  assign N89 = (N2)? 1'b0 :
               (N3)? N79 : 1'b0;
  assign { wbuf_entry_in_data__63_, wbuf_entry_in_data__62_, wbuf_entry_in_data__61_, wbuf_entry_in_data__60_, wbuf_entry_in_data__59_, wbuf_entry_in_data__58_, wbuf_entry_in_data__57_, wbuf_entry_in_data__56_, wbuf_entry_in_data__55_, wbuf_entry_in_data__54_, wbuf_entry_in_data__53_, wbuf_entry_in_data__52_, wbuf_entry_in_data__51_, wbuf_entry_in_data__50_, wbuf_entry_in_data__49_, wbuf_entry_in_data__48_, wbuf_entry_in_data__47_, wbuf_entry_in_data__46_, wbuf_entry_in_data__45_, wbuf_entry_in_data__44_, wbuf_entry_in_data__43_, wbuf_entry_in_data__42_, wbuf_entry_in_data__41_, wbuf_entry_in_data__40_, wbuf_entry_in_data__39_, wbuf_entry_in_data__38_, wbuf_entry_in_data__37_, wbuf_entry_in_data__36_, wbuf_entry_in_data__35_, wbuf_entry_in_data__34_, wbuf_entry_in_data__33_, wbuf_entry_in_data__32_, wbuf_entry_in_data__31_, wbuf_entry_in_data__30_, wbuf_entry_in_data__29_, wbuf_entry_in_data__28_, wbuf_entry_in_data__27_, wbuf_entry_in_data__26_, wbuf_entry_in_data__25_, wbuf_entry_in_data__24_, wbuf_entry_in_data__23_, wbuf_entry_in_data__22_, wbuf_entry_in_data__21_, wbuf_entry_in_data__20_, wbuf_entry_in_data__19_, wbuf_entry_in_data__18_, wbuf_entry_in_data__17_, wbuf_entry_in_data__16_, wbuf_entry_in_data__15_, wbuf_entry_in_data__14_, wbuf_entry_in_data__13_, wbuf_entry_in_data__12_, wbuf_entry_in_data__11_, wbuf_entry_in_data__10_, wbuf_entry_in_data__9_, wbuf_entry_in_data__8_ } = (N4)? data_tv_r[63:8] :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N94)? { data_tv_r[31:0], data_tv_r[31:8] } :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N97)? { data_tv_r[15:0], data_tv_r[15:0], data_tv_r[15:0], data_tv_r[15:8] } :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N92)? { data_tv_r[7:0], data_tv_r[7:0], data_tv_r[7:0], data_tv_r[7:0], data_tv_r[7:0], data_tv_r[7:0], data_tv_r[7:0] } : 1'b0;
  assign N4 = double_op_tv_r;
  assign { wbuf_entry_in_mask__7_, wbuf_entry_in_mask__6_, wbuf_entry_in_mask__5_, wbuf_entry_in_mask__4_, wbuf_entry_in_mask__3_, wbuf_entry_in_mask__2_, wbuf_entry_in_mask__1_, wbuf_entry_in_mask__0_ } = (N4)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } :
                                                                                                                                                                                                              (N121)? { paddr_tv_r[2:2], paddr_tv_r[2:2], paddr_tv_r[2:2], paddr_tv_r[2:2], N101, N102, N103, N104 } :
                                                                                                                                                                                                              (N123)? { N105, N106, N107, N108, N109, N110, N111, N112 } :
                                                                                                                                                                                                              (N100)? { N113, N114, N115, N116, N117, N118, N119, N120 } : 1'b0;
  assign lce_lru_way_li = (N5)? invalid_way :
                          (N6)? lru_encode : 1'b0;
  assign N5 = invalid_exist;
  assign N6 = N124;
  assign N129 = (N7)? uncached_load_data_v_r :
                (N133)? N128 :
                (N127)? 1'b0 : 1'b0;
  assign N7 = load_op_tv_r;
  assign N131 = (N8)? N129 :
                (N9)? N130 : 1'b0;
  assign N8 = uncached_tv_r;
  assign N9 = N437;
  assign v_o = (N10)? N131 :
               (N11)? 1'b0 : 1'b0;
  assign N10 = v_tv_r;
  assign N11 = N125;
  assign { N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139 } = (N4)? bypass_data_masked :
                                                                                                                                                                                                                                                                                                                                                                                                              (N205)? { genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_word_sigext, genblk4_data_word_selected } :
                                                                                                                                                                                                                                                                                                                                                                                                              (N207)? { genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_half_sigext, genblk4_data_half_selected } :
                                                                                                                                                                                                                                                                                                                                                                                                              (N138)? { genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_byte_sigext, genblk4_data_byte_selected } : 1'b0;
  assign data_o = (N12)? uncached_load_data_r :
                  (N204)? { N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139 } :
                  (N135)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = uncached_load_data_v_r;
  assign data_mem_v_li = (N13)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } :
                         (N213)? wbuf_data_mem_v :
                         (N211)? { lce_data_mem_v, lce_data_mem_v, lce_data_mem_v, lce_data_mem_v, lce_data_mem_v, lce_data_mem_v, lce_data_mem_v, lce_data_mem_v } : 1'b0;
  assign N13 = N208;
  assign data_mem_addr_li[8:0] = (N14)? dcache_pkt_i[75:67] :
                                 (N219)? wbuf_entry_out[86:78] :
                                 (N217)? lce_data_mem_pkt[522:514] : 1'b0;
  assign N14 = N214;
  assign data_mem_data_li[63:0] = (N15)? wbuf_entry_out[74:11] :
                                  (N16)? lce_data_mem_write_data[63:0] : 1'b0;
  assign N15 = N221;
  assign N16 = N220;
  assign data_mem_mask_li[7:0] = (N17)? wbuf_entry_out[10:3] :
                                 (N18)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N17 = N223;
  assign N18 = N222;
  assign data_mem_addr_li[17:9] = (N19)? dcache_pkt_i[75:67] :
                                  (N230)? wbuf_entry_out[86:78] :
                                  (N227)? { lce_data_mem_pkt[522:515], N228 } : 1'b0;
  assign N19 = N224;
  assign data_mem_data_li[127:64] = (N20)? wbuf_entry_out[74:11] :
                                    (N21)? lce_data_mem_write_data[127:64] : 1'b0;
  assign N20 = N232;
  assign N21 = N231;
  assign data_mem_mask_li[15:8] = (N22)? wbuf_entry_out[10:3] :
                                  (N23)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N22 = N234;
  assign N23 = N233;
  assign data_mem_addr_li[26:18] = (N24)? dcache_pkt_i[75:67] :
                                   (N241)? wbuf_entry_out[86:78] :
                                   (N238)? { lce_data_mem_pkt[522:516], N239, lce_data_mem_pkt[514:514] } : 1'b0;
  assign N24 = N235;
  assign data_mem_data_li[191:128] = (N25)? wbuf_entry_out[74:11] :
                                     (N26)? lce_data_mem_write_data[191:128] : 1'b0;
  assign N25 = N243;
  assign N26 = N242;
  assign data_mem_mask_li[23:16] = (N27)? wbuf_entry_out[10:3] :
                                   (N28)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N27 = N245;
  assign N28 = N244;
  assign data_mem_addr_li[35:27] = (N29)? dcache_pkt_i[75:67] :
                                   (N253)? wbuf_entry_out[86:78] :
                                   (N249)? { lce_data_mem_pkt[522:516], N250, N251 } : 1'b0;
  assign N29 = N246;
  assign data_mem_data_li[255:192] = (N30)? wbuf_entry_out[74:11] :
                                     (N31)? lce_data_mem_write_data[255:192] : 1'b0;
  assign N30 = N255;
  assign N31 = N254;
  assign data_mem_mask_li[31:24] = (N32)? wbuf_entry_out[10:3] :
                                   (N33)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N32 = N257;
  assign N33 = N256;
  assign data_mem_addr_li[44:36] = (N34)? dcache_pkt_i[75:67] :
                                   (N264)? wbuf_entry_out[86:78] :
                                   (N261)? { lce_data_mem_pkt[522:517], N262, lce_data_mem_pkt[515:514] } : 1'b0;
  assign N34 = N258;
  assign data_mem_data_li[319:256] = (N35)? wbuf_entry_out[74:11] :
                                     (N36)? lce_data_mem_write_data[319:256] : 1'b0;
  assign N35 = N266;
  assign N36 = N265;
  assign data_mem_mask_li[39:32] = (N37)? wbuf_entry_out[10:3] :
                                   (N38)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N37 = N268;
  assign N38 = N267;
  assign data_mem_addr_li[53:45] = (N39)? dcache_pkt_i[75:67] :
                                   (N276)? wbuf_entry_out[86:78] :
                                   (N272)? { lce_data_mem_pkt[522:517], N273, lce_data_mem_pkt[515:515], N274 } : 1'b0;
  assign N39 = N269;
  assign data_mem_data_li[383:320] = (N40)? wbuf_entry_out[74:11] :
                                     (N41)? lce_data_mem_write_data[383:320] : 1'b0;
  assign N40 = N278;
  assign N41 = N277;
  assign data_mem_mask_li[47:40] = (N42)? wbuf_entry_out[10:3] :
                                   (N43)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N42 = N280;
  assign N43 = N279;
  assign data_mem_addr_li[62:54] = (N44)? dcache_pkt_i[75:67] :
                                   (N288)? wbuf_entry_out[86:78] :
                                   (N284)? { lce_data_mem_pkt[522:517], N285, N286, lce_data_mem_pkt[514:514] } : 1'b0;
  assign N44 = N281;
  assign data_mem_data_li[447:384] = (N45)? wbuf_entry_out[74:11] :
                                     (N46)? lce_data_mem_write_data[447:384] : 1'b0;
  assign N45 = N290;
  assign N46 = N289;
  assign data_mem_mask_li[55:48] = (N47)? wbuf_entry_out[10:3] :
                                   (N48)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N47 = N292;
  assign N48 = N291;
  assign data_mem_addr_li[71:63] = (N49)? dcache_pkt_i[75:67] :
                                   (N301)? wbuf_entry_out[86:78] :
                                   (N296)? { lce_data_mem_pkt[522:517], N297, N298, N299 } : 1'b0;
  assign N49 = N293;
  assign data_mem_data_li[511:448] = (N50)? wbuf_entry_out[74:11] :
                                     (N51)? lce_data_mem_write_data[511:448] : 1'b0;
  assign N50 = N303;
  assign N51 = N302;
  assign data_mem_mask_li[63:56] = (N52)? wbuf_entry_out[10:3] :
                                   (N53)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N52 = N305;
  assign N53 = N304;
  assign tag_mem_addr_li = (N54)? dcache_pkt_i[75:70] :
                           (N55)? lce_tag_mem_pkt[22:17] : 1'b0;
  assign N54 = tl_we;
  assign N55 = N475;
  assign tag_mem_data_li = (N56)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                           (N57)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                           (N58)? { lce_tag_mem_pkt[13:2], lce_tag_mem_pkt[13:2], lce_tag_mem_pkt[13:2], lce_tag_mem_pkt[13:2], lce_tag_mem_pkt[13:2], lce_tag_mem_pkt[13:2], lce_tag_mem_pkt[13:2], lce_tag_mem_pkt[13:2] } :
                           (N59)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N56 = N308;
  assign N57 = N310;
  assign N58 = N312;
  assign N59 = N313;
  assign tag_mem_mask_li = (N56)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } :
                           (N57)? { lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                           (N58)? { lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:7], lce_tag_mem_way_one_hot[7:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:6], lce_tag_mem_way_one_hot[6:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:5], lce_tag_mem_way_one_hot[5:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:4], lce_tag_mem_way_one_hot[4:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:3], lce_tag_mem_way_one_hot[3:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:2], lce_tag_mem_way_one_hot[2:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:1], lce_tag_mem_way_one_hot[1:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0], lce_tag_mem_way_one_hot[0:0] } :
                           (N59)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stat_mem_w_li = (N10)? N314 :
                         (N11)? N315 : 1'b0;
  assign stat_mem_addr_li = (N10)? paddr_tv_r[11:6] :
                            (N11)? lce_stat_mem_pkt[10:5] : 1'b0;
  assign { N319, N318, N317 } = (N60)? store_hit_way :
                                (N61)? load_hit_way : 1'b0;
  assign N60 = store_op_tv_r;
  assign N61 = N316;
  assign { N328, N327, N326, N325, N324, N323, N322, N321 } = (N62)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } :
                                                              (N63)? dirty_mask_lo : 1'b0;
  assign N62 = N320;
  assign N63 = lce_stat_mem_pkt[1];
  assign { N337, N336, N335, N334, N333, N332, N331, N330, N329 } = (N64)? { N320, N328, N327, N326, N325, N324, N323, N322, N321 } :
                                                                    (N65)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N64 = N403;
  assign N65 = lce_stat_mem_pkt[0];
  assign lru_decode_way_li = (N66)? { N319, N318, N317 } :
                             (N11)? lce_stat_mem_pkt[4:2] : 1'b0;
  assign N66 = stat_mem_data_li[0];
  assign dirty_mask_way_li = (N66)? store_hit_way :
                             (N11)? lce_stat_mem_pkt[4:2] : 1'b0;
  assign dirty_mask_v_li = (N66)? store_op_tv_r :
                           (N11)? 1'b1 : 1'b0;
  assign stat_mem_data_li[14:1] = (N66)? { lru_decode_data_lo, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } :
                                  (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stat_mem_mask_li = (N66)? { lru_decode_mask_lo, dirty_mask_lo } :
                            (N11)? { N337, N337, N337, N337, N337, N337, N337, N336, N335, N334, N333, N332, N331, N330, N329 } : 1'b0;
  assign lce_data_mem_pkt_yumi = (N67)? lce_data_mem_pkt_v :
                                 (N68)? N339 : 1'b0;
  assign N67 = N420;
  assign N68 = N419;
  assign N345 = (N69)? 1'b1 :
                (N349)? 1'b1 :
                (N352)? 1'b1 :
                (N344)? 1'b0 : 1'b0;
  assign N69 = N341;
  assign N346 = (N69)? 1'b0 :
                (N349)? 1'b1 :
                (N352)? 1'b0 : 1'b0;
  assign N347 = (N69)? 1'b0 :
                (N349)? 1'b1 :
                (N352)? 1'b0 :
                (N344)? 1'b0 : 1'b0;
  assign load_op = ~dcache_pkt_i[79];
  assign signed_op = ~dcache_pkt_i[78];
  assign tl_we = N421 & N422;
  assign N421 = v_i & ready_o;
  assign N422 = ~poison_i;
  assign N70 = ~reset_i;
  assign N71 = reset_i;
  assign N72 = tl_we & dcache_pkt_i[79];
  assign n_0_net_ = N423 & tag_mem_v_li;
  assign N423 = ~reset_i;
  assign n_1_net_ = N424 & data_mem_v_li[0];
  assign N424 = ~reset_i;
  assign n_2_net_ = N425 & data_mem_v_li[1];
  assign N425 = ~reset_i;
  assign n_3_net_ = N426 & data_mem_v_li[2];
  assign N426 = ~reset_i;
  assign n_4_net_ = N427 & data_mem_v_li[3];
  assign N427 = ~reset_i;
  assign n_5_net_ = N428 & data_mem_v_li[4];
  assign N428 = ~reset_i;
  assign n_6_net_ = N429 & data_mem_v_li[5];
  assign N429 = ~reset_i;
  assign n_7_net_ = N430 & data_mem_v_li[6];
  assign N430 = ~reset_i;
  assign n_8_net_ = N431 & data_mem_v_li[7];
  assign N431 = ~reset_i;
  assign tv_we = N432 & N433;
  assign N432 = v_tl_r & N422;
  assign N433 = ~tlb_miss_i;
  assign N76 = ~reset_i;
  assign N77 = reset_i;
  assign N78 = tv_we & load_op_tl_r;
  assign N79 = tv_we & store_op_tl_r;
  assign load_hit_tv[0] = tag_match_tv[0] & N378;
  assign store_hit_tv[0] = tag_match_tv[0] & N402;
  assign load_hit_tv[1] = tag_match_tv[1] & N377;
  assign store_hit_tv[1] = tag_match_tv[1] & N399;
  assign load_hit_tv[2] = tag_match_tv[2] & N376;
  assign store_hit_tv[2] = tag_match_tv[2] & N396;
  assign load_hit_tv[3] = tag_match_tv[3] & N375;
  assign store_hit_tv[3] = tag_match_tv[3] & N393;
  assign load_hit_tv[4] = tag_match_tv[4] & N374;
  assign store_hit_tv[4] = tag_match_tv[4] & N390;
  assign load_hit_tv[5] = tag_match_tv[5] & N373;
  assign store_hit_tv[5] = tag_match_tv[5] & N387;
  assign load_hit_tv[6] = tag_match_tv[6] & N372;
  assign store_hit_tv[6] = tag_match_tv[6] & N384;
  assign load_hit_tv[7] = tag_match_tv[7] & N371;
  assign store_hit_tv[7] = tag_match_tv[7] & N381;
  assign load_miss_tv = N436 & N437;
  assign N436 = N435 & load_op_tv_r;
  assign N435 = N434 & v_tv_r;
  assign N434 = ~load_hit;
  assign N437 = ~uncached_tv_r;
  assign store_miss_tv = N440 & N437;
  assign N440 = N439 & store_op_tv_r;
  assign N439 = N438 & v_tv_r;
  assign N438 = ~store_hit;
  assign uncached_load_req = N442 & N443;
  assign N442 = N441 & uncached_tv_r;
  assign N441 = v_tv_r & load_op_tv_r;
  assign N443 = ~uncached_load_data_v_r;
  assign uncached_store_req = N444 & uncached_tv_r;
  assign N444 = v_tv_r & store_op_tv_r;
  assign N90 = word_op_tv_r | double_op_tv_r;
  assign N91 = half_op_tv_r | N90;
  assign N92 = ~N91;
  assign N93 = ~double_op_tv_r;
  assign N94 = word_op_tv_r & N93;
  assign N95 = ~word_op_tv_r;
  assign N96 = N93 & N95;
  assign N97 = half_op_tv_r & N96;
  assign N98 = word_op_tv_r | double_op_tv_r;
  assign N99 = half_op_tv_r | N98;
  assign N100 = ~N99;
  assign N101 = ~paddr_tv_r[2];
  assign N102 = ~paddr_tv_r[2];
  assign N103 = ~paddr_tv_r[2];
  assign N104 = ~paddr_tv_r[2];
  assign N105 = paddr_tv_r[2] & paddr_tv_r[1];
  assign N106 = paddr_tv_r[2] & paddr_tv_r[1];
  assign N107 = paddr_tv_r[2] & N445;
  assign N445 = ~paddr_tv_r[1];
  assign N108 = paddr_tv_r[2] & N446;
  assign N446 = ~paddr_tv_r[1];
  assign N109 = N447 & paddr_tv_r[1];
  assign N447 = ~paddr_tv_r[2];
  assign N110 = N448 & paddr_tv_r[1];
  assign N448 = ~paddr_tv_r[2];
  assign N111 = N449 & N450;
  assign N449 = ~paddr_tv_r[2];
  assign N450 = ~paddr_tv_r[1];
  assign N112 = N451 & N452;
  assign N451 = ~paddr_tv_r[2];
  assign N452 = ~paddr_tv_r[1];
  assign N113 = N453 & paddr_tv_r[0];
  assign N453 = paddr_tv_r[2] & paddr_tv_r[1];
  assign N114 = N454 & N455;
  assign N454 = paddr_tv_r[2] & paddr_tv_r[1];
  assign N455 = ~paddr_tv_r[0];
  assign N115 = N457 & paddr_tv_r[0];
  assign N457 = paddr_tv_r[2] & N456;
  assign N456 = ~paddr_tv_r[1];
  assign N116 = N459 & N460;
  assign N459 = paddr_tv_r[2] & N458;
  assign N458 = ~paddr_tv_r[1];
  assign N460 = ~paddr_tv_r[0];
  assign N117 = N462 & paddr_tv_r[0];
  assign N462 = N461 & paddr_tv_r[1];
  assign N461 = ~paddr_tv_r[2];
  assign N118 = N464 & N465;
  assign N464 = N463 & paddr_tv_r[1];
  assign N463 = ~paddr_tv_r[2];
  assign N465 = ~paddr_tv_r[0];
  assign N119 = N468 & paddr_tv_r[0];
  assign N468 = N466 & N467;
  assign N466 = ~paddr_tv_r[2];
  assign N467 = ~paddr_tv_r[1];
  assign N120 = N471 & N472;
  assign N471 = N469 & N470;
  assign N469 = ~paddr_tv_r[2];
  assign N470 = ~paddr_tv_r[1];
  assign N472 = ~paddr_tv_r[0];
  assign N121 = word_op_tv_r & N93;
  assign N122 = N93 & N95;
  assign N123 = half_op_tv_r & N122;
  assign n_10_net_ = N473 & stat_mem_v_li;
  assign N473 = ~reset_i;
  assign N124 = ~invalid_exist;
  assign N125 = ~v_tv_r;
  assign N126 = store_op_tv_r | load_op_tv_r;
  assign N127 = ~N126;
  assign N128 = ~cache_miss_o;
  assign N130 = v_tv_r & N128;
  assign N132 = ~load_op_tv_r;
  assign N133 = store_op_tv_r & N132;
  assign n_13_net__2_ = load_hit_way[2] ^ paddr_tv_r[5];
  assign n_13_net__1_ = load_hit_way[1] ^ paddr_tv_r[4];
  assign n_13_net__0_ = load_hit_way[0] ^ paddr_tv_r[3];
  assign genblk4_word_sigext = signed_op_tv_r & genblk4_data_word_selected[31];
  assign genblk4_half_sigext = signed_op_tv_r & genblk4_data_half_selected[15];
  assign genblk4_byte_sigext = signed_op_tv_r & genblk4_data_byte_selected[7];
  assign N134 = load_op_tv_r | uncached_load_data_v_r;
  assign N135 = ~N134;
  assign N136 = word_op_tv_r | double_op_tv_r;
  assign N137 = half_op_tv_r | N136;
  assign N138 = ~N137;
  assign N203 = ~uncached_load_data_v_r;
  assign N204 = load_op_tv_r & N203;
  assign N205 = word_op_tv_r & N93;
  assign N206 = N93 & N95;
  assign N207 = half_op_tv_r & N206;
  assign n_14_net__2_ = wbuf_entry_out[2] ^ wbuf_entry_out[80];
  assign n_14_net__1_ = wbuf_entry_out[1] ^ wbuf_entry_out[79];
  assign n_14_net__0_ = wbuf_entry_out[0] ^ wbuf_entry_out[78];
  assign lce_data_mem_v = N406 & lce_data_mem_pkt_yumi;
  assign N208 = load_op & tl_we;
  assign N209 = wbuf_yumi_li;
  assign N210 = N209 | N208;
  assign N211 = ~N210;
  assign N212 = ~N208;
  assign N213 = N209 & N212;
  assign data_mem_w_li = wbuf_yumi_li | N474;
  assign N474 = lce_data_mem_pkt_yumi & N370;
  assign N214 = load_op & tl_we;
  assign N215 = wbuf_yumi_li;
  assign N216 = N215 | N214;
  assign N217 = ~N216;
  assign N218 = ~N214;
  assign N219 = N215 & N218;
  assign N220 = ~wbuf_yumi_li;
  assign N221 = wbuf_yumi_li;
  assign N222 = ~wbuf_yumi_li;
  assign N223 = wbuf_yumi_li;
  assign N224 = load_op & tl_we;
  assign N225 = wbuf_yumi_li;
  assign N226 = N225 | N224;
  assign N227 = ~N226;
  assign N228 = ~lce_data_mem_pkt[514];
  assign N229 = ~N224;
  assign N230 = N225 & N229;
  assign N231 = ~wbuf_yumi_li;
  assign N232 = wbuf_yumi_li;
  assign N233 = ~wbuf_yumi_li;
  assign N234 = wbuf_yumi_li;
  assign N235 = load_op & tl_we;
  assign N236 = wbuf_yumi_li;
  assign N237 = N236 | N235;
  assign N238 = ~N237;
  assign N239 = ~lce_data_mem_pkt[515];
  assign N240 = ~N235;
  assign N241 = N236 & N240;
  assign N242 = ~wbuf_yumi_li;
  assign N243 = wbuf_yumi_li;
  assign N244 = ~wbuf_yumi_li;
  assign N245 = wbuf_yumi_li;
  assign N246 = load_op & tl_we;
  assign N247 = wbuf_yumi_li;
  assign N248 = N247 | N246;
  assign N249 = ~N248;
  assign N250 = ~lce_data_mem_pkt[515];
  assign N251 = ~lce_data_mem_pkt[514];
  assign N252 = ~N246;
  assign N253 = N247 & N252;
  assign N254 = ~wbuf_yumi_li;
  assign N255 = wbuf_yumi_li;
  assign N256 = ~wbuf_yumi_li;
  assign N257 = wbuf_yumi_li;
  assign N258 = load_op & tl_we;
  assign N259 = wbuf_yumi_li;
  assign N260 = N259 | N258;
  assign N261 = ~N260;
  assign N262 = ~lce_data_mem_pkt[516];
  assign N263 = ~N258;
  assign N264 = N259 & N263;
  assign N265 = ~wbuf_yumi_li;
  assign N266 = wbuf_yumi_li;
  assign N267 = ~wbuf_yumi_li;
  assign N268 = wbuf_yumi_li;
  assign N269 = load_op & tl_we;
  assign N270 = wbuf_yumi_li;
  assign N271 = N270 | N269;
  assign N272 = ~N271;
  assign N273 = ~lce_data_mem_pkt[516];
  assign N274 = ~lce_data_mem_pkt[514];
  assign N275 = ~N269;
  assign N276 = N270 & N275;
  assign N277 = ~wbuf_yumi_li;
  assign N278 = wbuf_yumi_li;
  assign N279 = ~wbuf_yumi_li;
  assign N280 = wbuf_yumi_li;
  assign N281 = load_op & tl_we;
  assign N282 = wbuf_yumi_li;
  assign N283 = N282 | N281;
  assign N284 = ~N283;
  assign N285 = ~lce_data_mem_pkt[516];
  assign N286 = ~lce_data_mem_pkt[515];
  assign N287 = ~N281;
  assign N288 = N282 & N287;
  assign N289 = ~wbuf_yumi_li;
  assign N290 = wbuf_yumi_li;
  assign N291 = ~wbuf_yumi_li;
  assign N292 = wbuf_yumi_li;
  assign N293 = load_op & tl_we;
  assign N294 = wbuf_yumi_li;
  assign N295 = N294 | N293;
  assign N296 = ~N295;
  assign N297 = ~lce_data_mem_pkt[516];
  assign N298 = ~lce_data_mem_pkt[515];
  assign N299 = ~lce_data_mem_pkt[514];
  assign N300 = ~N293;
  assign N301 = N294 & N300;
  assign N302 = ~wbuf_yumi_li;
  assign N303 = wbuf_yumi_li;
  assign N304 = ~wbuf_yumi_li;
  assign N305 = wbuf_yumi_li;
  assign tag_mem_v_li = tl_we | lce_tag_mem_pkt_yumi;
  assign tag_mem_w_li = N475 & lce_tag_mem_pkt_v;
  assign N475 = ~tl_we;
  assign N306 = ~lce_tag_mem_pkt[1];
  assign N307 = ~lce_tag_mem_pkt[0];
  assign N310 = ~N309;
  assign N312 = ~N311;
  assign stat_mem_v_li = N476 | lce_stat_mem_pkt_yumi;
  assign N476 = v_tv_r & N437;
  assign N314 = ~N477;
  assign N477 = load_miss_tv | store_miss_tv;
  assign N315 = lce_stat_mem_pkt_yumi & N404;
  assign stat_mem_data_li[0] = v_tv_r;
  assign N316 = ~store_op_tv_r;
  assign N320 = ~lce_stat_mem_pkt[1];
  assign wbuf_v_li = N478 & store_hit;
  assign N478 = v_tv_r & store_op_tv_r;
  assign wbuf_yumi_li = wbuf_v_lo & N480;
  assign N480 = ~N479;
  assign N479 = load_op & tl_we;
  assign bypass_v_li = tv_we & load_op_tl_r;
  assign N338 = lce_data_mem_pkt_yumi & N416;
  assign N339 = N486 & lce_data_mem_pkt_v;
  assign N486 = N484 & N485;
  assign N484 = N482 & N483;
  assign N482 = ~N481;
  assign N481 = load_op & tl_we;
  assign N483 = ~wbuf_v_lo;
  assign N485 = ~lce_snoop_match_lo;
  assign N340 = lce_data_mem_pkt_yumi & N418;
  assign N341 = reset_i;
  assign N342 = N340 | N341;
  assign N343 = v_o | N342;
  assign N344 = ~N343;
  assign N348 = ~N341;
  assign N349 = N340 & N348;
  assign N350 = ~N340;
  assign N351 = N348 & N350;
  assign N352 = v_o & N351;
  assign lce_tag_mem_pkt_yumi = lce_tag_mem_pkt_v & N475;
  assign lce_stat_mem_pkt_yumi = N488 & lce_stat_mem_pkt_v;
  assign N488 = ~N487;
  assign N487 = v_tv_r & N437;

  always @(posedge clk_i) begin
    if(N75) begin
      { data_tl_r[63:0] } <= { dcache_pkt_i[63:0] };
    end
    if(1'b1) begin
      v_tl_r <= N73;
      v_tv_r <= N80;
    end
    if(N74) begin
      { page_offset_tl_r[11:0] } <= { dcache_pkt_i[75:64] };
      load_op_tl_r <= load_op;
      store_op_tl_r <= dcache_pkt_i[79];
      signed_op_tl_r <= signed_op;
      { size_op_tl_r[1:0] } <= { dcache_pkt_i[77:76] };
      double_op_tl_r <= N407;
      word_op_tl_r <= N410;
      half_op_tl_r <= N413;
    end
    if(N89) begin
      { data_tv_r[63:0] } <= { data_tl_r[63:0] };
    end
    if(N81) begin
      uncached_tv_r <= uncached_i;
      load_op_tv_r <= load_op_tl_r;
      { paddr_tv_r[21:20] } <= { ptag_i[9:8] };
      { tag_info_tv_r[95:0] } <= { tag_mem_data_lo[95:0] };
    end
    if(N82) begin
      store_op_tv_r <= store_op_tl_r;
      signed_op_tv_r <= signed_op_tl_r;
      { size_op_tv_r[1:0] } <= { size_op_tl_r[1:0] };
      double_op_tv_r <= double_op_tl_r;
      word_op_tv_r <= word_op_tl_r;
      half_op_tv_r <= half_op_tl_r;
      { paddr_tv_r[19:0] } <= { ptag_i[7:0], page_offset_tl_r[11:0] };
    end
    if(N83) begin
      { ld_data_tv_r[511:413], ld_data_tv_r[0:0] } <= { data_mem_data_lo[511:413], data_mem_data_lo[0:0] };
    end
    if(N84) begin
      { ld_data_tv_r[412:314], ld_data_tv_r[1:1] } <= { data_mem_data_lo[412:314], data_mem_data_lo[1:1] };
    end
    if(N85) begin
      { ld_data_tv_r[313:215], ld_data_tv_r[2:2] } <= { data_mem_data_lo[313:215], data_mem_data_lo[2:2] };
    end
    if(N86) begin
      { ld_data_tv_r[214:116], ld_data_tv_r[3:3] } <= { data_mem_data_lo[214:116], data_mem_data_lo[3:3] };
    end
    if(N87) begin
      { ld_data_tv_r[115:17], ld_data_tv_r[4:4] } <= { data_mem_data_lo[115:17], data_mem_data_lo[4:4] };
    end
    if(N88) begin
      { ld_data_tv_r[16:5] } <= { data_mem_data_lo[16:5] };
    end
    if(N338) begin
      { lce_data_mem_pkt_way_r[2:0] } <= { lce_data_mem_pkt[516:514] };
    end
    if(N347) begin
      { uncached_load_data_r[63:0] } <= { lce_data_mem_pkt[65:2] };
    end
    if(N345) begin
      uncached_load_data_v_r <= N346;
    end
  end


endmodule



module bp_be_mmu_top_vaddr_width_p39_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36_num_cce_p1_num_lce_p2_cce_block_size_in_bytes_p64_lce_assoc_p8_lce_sets_p64
(
  clk_i,
  reset_i,
  mmu_cmd_i,
  mmu_cmd_v_i,
  mmu_cmd_ready_o,
  chk_poison_ex_i,
  mmu_resp_o,
  mmu_resp_v_o,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i,
  dcache_id_i
);

  input [106:0] mmu_cmd_i;
  output [72:0] mmu_resp_o;
  output [96:0] lce_req_o;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  input [35:0] lce_cmd_i;
  input [517:0] lce_data_cmd_i;
  output [517:0] lce_data_cmd_o;
  input [0:0] dcache_id_i;
  input clk_i;
  input reset_i;
  input mmu_cmd_v_i;
  input chk_poison_ex_i;
  input lce_req_ready_i;
  input lce_resp_ready_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_v_i;
  input lce_data_cmd_ready_i;
  output mmu_cmd_ready_o;
  output mmu_resp_v_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_ready_o;
  output lce_data_cmd_ready_o;
  output lce_data_cmd_v_o;
  wire [72:0] mmu_resp_o;
  wire [96:0] lce_req_o;
  wire [25:0] lce_resp_o;
  wire [536:0] lce_data_resp_o;
  wire [517:0] lce_data_cmd_o;
  wire mmu_cmd_ready_o,mmu_resp_v_o,lce_req_v_o,lce_resp_v_o,lce_data_resp_v_o,
  lce_cmd_ready_o,lce_data_cmd_ready_o,lce_data_cmd_v_o,mmu_resp_o_8,mmu_resp_o_7,
  mmu_resp_o_6,mmu_resp_o_5,mmu_resp_o_4,mmu_resp_o_3,mmu_resp_o_2,mmu_resp_o_1,
  dcache_ready,N0;
  reg [9:0] ptag_r;

  bp_be_dcache_data_width_p64_paddr_width_p22_sets_p64_ways_p8_num_cce_p1_num_lce_p2
  dcache
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .lce_id_i(dcache_id_i[0]),
    .dcache_pkt_i({ mmu_cmd_i[106:103], mmu_cmd_i[75:0] }),
    .v_i(mmu_cmd_v_i),
    .ready_o(dcache_ready),
    .data_o(mmu_resp_o[72:9]),
    .v_o(mmu_resp_v_o),
    .tlb_miss_i(1'b0),
    .ptag_i(ptag_r),
    .uncached_i(1'b0),
    .cache_miss_o(mmu_resp_o[0]),
    .poison_i(chk_poison_ex_i),
    .lce_req_o(lce_req_o),
    .lce_req_v_o(lce_req_v_o),
    .lce_req_ready_i(lce_req_ready_i),
    .lce_resp_o(lce_resp_o),
    .lce_resp_v_o(lce_resp_v_o),
    .lce_resp_ready_i(lce_resp_ready_i),
    .lce_data_resp_o(lce_data_resp_o),
    .lce_data_resp_v_o(lce_data_resp_v_o),
    .lce_data_resp_ready_i(lce_data_resp_ready_i),
    .lce_cmd_i(lce_cmd_i),
    .lce_cmd_v_i(lce_cmd_v_i),
    .lce_cmd_ready_o(lce_cmd_ready_o),
    .lce_data_cmd_i(lce_data_cmd_i),
    .lce_data_cmd_v_i(lce_data_cmd_v_i),
    .lce_data_cmd_ready_o(lce_data_cmd_ready_o),
    .lce_data_cmd_o(lce_data_cmd_o),
    .lce_data_cmd_v_o(lce_data_cmd_v_o),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_i)
  );

  assign mmu_cmd_ready_o = dcache_ready & N0;
  assign N0 = ~mmu_resp_o[0];

  always @(posedge clk_i) begin
    if(1'b1) begin
      { ptag_r[9:0] } <= { mmu_cmd_i[85:76] };
    end
  end


endmodule



module bp_be_top_vaddr_width_p39_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36_core_els_p1_trace_p0_num_cce_p1_num_lce_p2_lce_assoc_p8_lce_sets_p64_cce_block_size_in_bytes_p64
(
  clk_i,
  reset_i,
  fe_queue_i,
  fe_queue_v_i,
  fe_queue_ready_o,
  fe_queue_clr_o,
  fe_queue_dequeue_o,
  fe_queue_rollback_o,
  fe_cmd_o,
  fe_cmd_v_o,
  fe_cmd_ready_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i,
  proc_cfg_i,
  cmt_rd_w_v_o,
  cmt_rd_addr_o,
  cmt_mem_w_v_o,
  cmt_mem_addr_o,
  cmt_mem_op_o,
  cmt_data_o
);

  input [133:0] fe_queue_i;
  output [108:0] fe_cmd_o;
  output [96:0] lce_req_o;
  output [25:0] lce_resp_o;
  output [536:0] lce_data_resp_o;
  input [35:0] lce_cmd_i;
  input [517:0] lce_data_cmd_i;
  output [517:0] lce_data_cmd_o;
  input [2:0] proc_cfg_i;
  output [4:0] cmt_rd_addr_o;
  output [63:0] cmt_mem_addr_o;
  output [3:0] cmt_mem_op_o;
  output [63:0] cmt_data_o;
  input clk_i;
  input reset_i;
  input fe_queue_v_i;
  input fe_cmd_ready_i;
  input lce_req_ready_i;
  input lce_resp_ready_i;
  input lce_data_resp_ready_i;
  input lce_cmd_v_i;
  input lce_data_cmd_v_i;
  input lce_data_cmd_ready_i;
  output fe_queue_ready_o;
  output fe_queue_clr_o;
  output fe_queue_dequeue_o;
  output fe_queue_rollback_o;
  output fe_cmd_v_o;
  output lce_req_v_o;
  output lce_resp_v_o;
  output lce_data_resp_v_o;
  output lce_cmd_ready_o;
  output lce_data_cmd_ready_o;
  output lce_data_cmd_v_o;
  output cmt_rd_w_v_o;
  output cmt_mem_w_v_o;
  wire [108:0] fe_cmd_o;
  wire [96:0] lce_req_o;
  wire [25:0] lce_resp_o;
  wire [536:0] lce_data_resp_o;
  wire [517:0] lce_data_cmd_o;
  wire [4:0] cmt_rd_addr_o;
  wire [63:0] cmt_mem_addr_o,cmt_data_o,chk_mtvec_li,chk_mtvec_lo,chk_mepc_li,chk_mepc_lo;
  wire [3:0] cmt_mem_op_o;
  wire fe_queue_ready_o,fe_queue_clr_o,fe_queue_dequeue_o,fe_queue_rollback_o,
  fe_cmd_v_o,lce_req_v_o,lce_resp_v_o,lce_data_resp_v_o,lce_cmd_ready_o,
  lce_data_cmd_ready_o,lce_data_cmd_v_o,cmt_rd_w_v_o,cmt_mem_w_v_o,chk_dispatch_v,chk_roll,
  chk_poison_isd,chk_poison_ex1,chk_poison_ex2,chk_poison_ex3,mmu_cmd_rdy,issue_pkt_v,
  issue_pkt_rdy,chk_mtvec_w_v_li,chk_mepc_w_v_li,mmu_cmd_v,mmu_resp_v,mmu_resp_rdy;
  wire [306:0] calc_status;
  wire [220:0] issue_pkt;
  wire [106:0] mmu_cmd;
  wire [72:0] mmu_resp;

  bp_be_checker_top_vaddr_width_p39_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36_load_to_use_forwarding_p1
  be_checker
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .fe_cmd_o(fe_cmd_o),
    .fe_cmd_v_o(fe_cmd_v_o),
    .fe_cmd_ready_i(fe_cmd_ready_i),
    .fe_queue_i(fe_queue_i),
    .fe_queue_v_i(fe_queue_v_i),
    .fe_queue_ready_o(fe_queue_ready_o),
    .chk_roll_fe_o(fe_queue_rollback_o),
    .chk_flush_fe_o(fe_queue_clr_o),
    .chk_dequeue_fe_o(fe_queue_dequeue_o),
    .issue_pkt_o(issue_pkt),
    .issue_pkt_v_o(issue_pkt_v),
    .issue_pkt_ready_i(issue_pkt_rdy),
    .calc_status_i(calc_status),
    .mmu_cmd_ready_i(mmu_cmd_rdy),
    .chk_dispatch_v_o(chk_dispatch_v),
    .chk_roll_o(chk_roll),
    .chk_poison_isd_o(chk_poison_isd),
    .chk_poison_ex1_o(chk_poison_ex1),
    .chk_poison_ex2_o(chk_poison_ex2),
    .chk_poison_ex3_o(chk_poison_ex3),
    .mtvec_i(chk_mtvec_li),
    .mtvec_w_v_i(chk_mtvec_w_v_li),
    .mtvec_o(chk_mtvec_lo),
    .mepc_i(chk_mepc_li),
    .mepc_w_v_i(chk_mepc_w_v_li),
    .mepc_o(chk_mepc_lo)
  );


  bp_be_calculator_top_vaddr_width_p39_paddr_width_p22_asid_width_p10_core_els_p1_num_lce_p2_lce_sets_p64_trace_p0_debug_p0_debug_file_pinv
  be_calculator
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .proc_cfg_i(proc_cfg_i),
    .issue_pkt_i(issue_pkt),
    .issue_pkt_v_i(issue_pkt_v),
    .issue_pkt_ready_o(issue_pkt_rdy),
    .chk_dispatch_v_i(chk_dispatch_v),
    .chk_roll_i(chk_roll),
    .chk_poison_isd_i(chk_poison_isd),
    .chk_poison_ex1_i(chk_poison_ex1),
    .chk_poison_ex2_i(chk_poison_ex2),
    .chk_poison_ex3_i(chk_poison_ex3),
    .calc_status_o(calc_status),
    .mmu_cmd_o(mmu_cmd),
    .mmu_cmd_v_o(mmu_cmd_v),
    .mmu_cmd_ready_i(mmu_cmd_rdy),
    .mmu_resp_i(mmu_resp),
    .mmu_resp_v_i(mmu_resp_v),
    .mmu_resp_ready_o(mmu_resp_rdy),
    .mtvec_o(chk_mtvec_li),
    .mtvec_w_v_o(chk_mtvec_w_v_li),
    .mtvec_i(chk_mtvec_lo),
    .mepc_o(chk_mepc_li),
    .mepc_w_v_o(chk_mepc_w_v_li),
    .mepc_i(chk_mepc_lo),
    .cmt_rd_w_v_o(cmt_rd_w_v_o),
    .cmt_rd_addr_o(cmt_rd_addr_o),
    .cmt_mem_w_v_o(cmt_mem_w_v_o),
    .cmt_mem_addr_o(cmt_mem_addr_o),
    .cmt_mem_op_o(cmt_mem_op_o),
    .cmt_data_o(cmt_data_o)
  );


  bp_be_mmu_top_vaddr_width_p39_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36_num_cce_p1_num_lce_p2_cce_block_size_in_bytes_p64_lce_assoc_p8_lce_sets_p64
  be_mmu
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .mmu_cmd_i(mmu_cmd),
    .mmu_cmd_v_i(mmu_cmd_v),
    .mmu_cmd_ready_o(mmu_cmd_rdy),
    .chk_poison_ex_i(chk_poison_ex2),
    .mmu_resp_o(mmu_resp),
    .mmu_resp_v_o(mmu_resp_v),
    .lce_req_o(lce_req_o),
    .lce_req_v_o(lce_req_v_o),
    .lce_req_ready_i(lce_req_ready_i),
    .lce_resp_o(lce_resp_o),
    .lce_resp_v_o(lce_resp_v_o),
    .lce_resp_ready_i(lce_resp_ready_i),
    .lce_data_resp_o(lce_data_resp_o),
    .lce_data_resp_v_o(lce_data_resp_v_o),
    .lce_data_resp_ready_i(lce_data_resp_ready_i),
    .lce_cmd_i(lce_cmd_i),
    .lce_cmd_v_i(lce_cmd_v_i),
    .lce_cmd_ready_o(lce_cmd_ready_o),
    .lce_data_cmd_i(lce_data_cmd_i),
    .lce_data_cmd_v_i(lce_data_cmd_v_i),
    .lce_data_cmd_ready_o(lce_data_cmd_ready_o),
    .lce_data_cmd_o(lce_data_cmd_o),
    .lce_data_cmd_v_o(lce_data_cmd_v_o),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_i),
    .dcache_id_i(proc_cfg_i[0])
  );


endmodule



module bp_core_core_els_p1_num_lce_p2_num_cce_p1_lce_assoc_p8_lce_sets_p64_cce_block_size_in_bytes_p64_data_width_p64_vaddr_width_p39_paddr_width_p22_branch_metadata_fwd_width_p36_asid_width_p10_btb_indx_width_p9_bht_indx_width_p5_ras_addr_width_p22_trace_p0
(
  clk_i,
  reset_i,
  proc_cfg_i,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i,
  cmt_rd_w_v_o,
  cmt_rd_addr_o,
  cmt_mem_w_v_o,
  cmt_mem_addr_o,
  cmt_mem_op_o,
  cmt_data_o
);

  input [2:0] proc_cfg_i;
  output [193:0] lce_req_o;
  output [1:0] lce_req_v_o;
  input [1:0] lce_req_ready_i;
  output [51:0] lce_resp_o;
  output [1:0] lce_resp_v_o;
  input [1:0] lce_resp_ready_i;
  output [1073:0] lce_data_resp_o;
  output [1:0] lce_data_resp_v_o;
  input [1:0] lce_data_resp_ready_i;
  input [71:0] lce_cmd_i;
  input [1:0] lce_cmd_v_i;
  output [1:0] lce_cmd_ready_o;
  input [1035:0] lce_data_cmd_i;
  input [1:0] lce_data_cmd_v_i;
  output [1:0] lce_data_cmd_ready_o;
  output [1035:0] lce_data_cmd_o;
  output [1:0] lce_data_cmd_v_o;
  input [1:0] lce_data_cmd_ready_i;
  output [4:0] cmt_rd_addr_o;
  output [63:0] cmt_mem_addr_o;
  output [3:0] cmt_mem_op_o;
  output [63:0] cmt_data_o;
  input clk_i;
  input reset_i;
  output cmt_rd_w_v_o;
  output cmt_mem_w_v_o;
  wire [193:0] lce_req_o;
  wire [1:0] lce_req_v_o,lce_resp_v_o,lce_data_resp_v_o,lce_cmd_ready_o,lce_data_cmd_ready_o,
  lce_data_cmd_v_o;
  wire [51:0] lce_resp_o;
  wire [1073:0] lce_data_resp_o;
  wire [1035:0] lce_data_cmd_o;
  wire [4:0] cmt_rd_addr_o;
  wire [63:0] cmt_mem_addr_o,cmt_data_o;
  wire [3:0] cmt_mem_op_o;
  wire cmt_rd_w_v_o,cmt_mem_w_v_o,fe_fe_queue_v,fe_fe_queue_ready,be_fe_queue_v,
  be_fe_queue_ready;
  wire [133:0] fe_fe_queue,be_fe_queue;
  wire [108:0] fe_fe_cmd,be_fe_cmd;
  wire [0:0] fe_fe_cmd_v,fe_fe_cmd_ready,fe_queue_clr,fe_queue_dequeue,fe_queue_rollback,
  be_fe_cmd_v,be_fe_cmd_ready;

  bp_fe_top_39_22_1_2_8_64_64_9_5_22_10_80000124
  fe
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .icache_id_i(proc_cfg_i[1]),
    .fe_cmd_i(fe_fe_cmd),
    .fe_cmd_v_i(fe_fe_cmd_v[0]),
    .fe_cmd_ready_o(fe_fe_cmd_ready[0]),
    .fe_queue_o(fe_fe_queue),
    .fe_queue_v_o(fe_fe_queue_v),
    .fe_queue_ready_i(fe_fe_queue_ready),
    .lce_req_o(lce_req_o[96:0]),
    .lce_req_v_o(lce_req_v_o[0]),
    .lce_req_ready_i(lce_req_ready_i[0]),
    .lce_resp_o(lce_resp_o[25:0]),
    .lce_resp_v_o(lce_resp_v_o[0]),
    .lce_resp_ready_i(lce_resp_ready_i[0]),
    .lce_data_resp_o(lce_data_resp_o[536:0]),
    .lce_data_resp_v_o(lce_data_resp_v_o[0]),
    .lce_data_resp_ready_i(lce_data_resp_ready_i[0]),
    .lce_cmd_i(lce_cmd_i[35:0]),
    .lce_cmd_v_i(lce_cmd_v_i[0]),
    .lce_cmd_ready_o(lce_cmd_ready_o[0]),
    .lce_data_cmd_i(lce_data_cmd_i[517:0]),
    .lce_data_cmd_v_i(lce_data_cmd_v_i[0]),
    .lce_data_cmd_ready_o(lce_data_cmd_ready_o[0]),
    .lce_data_cmd_o(lce_data_cmd_o[517:0]),
    .lce_data_cmd_v_o(lce_data_cmd_v_o[0]),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_i[0])
  );


  bsg_fifo_1r1w_rolly_width_p134_els_p8_ready_THEN_valid_p1
  fe_queue_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clr_v_i(fe_queue_clr[0]),
    .ckpt_v_i(fe_queue_dequeue[0]),
    .roll_v_i(fe_queue_rollback[0]),
    .data_i(fe_fe_queue),
    .v_i(fe_fe_queue_v),
    .ready_o(fe_fe_queue_ready),
    .data_o(be_fe_queue),
    .v_o(be_fe_queue_v),
    .yumi_i(be_fe_queue_ready)
  );


  bsg_fifo_1r1w_small_width_p109_els_p2_ready_THEN_valid_p1
  fe_cmd_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(be_fe_cmd_v[0]),
    .ready_o(be_fe_cmd_ready[0]),
    .data_i(be_fe_cmd),
    .v_o(fe_fe_cmd_v[0]),
    .data_o(fe_fe_cmd),
    .yumi_i(fe_fe_cmd_ready[0])
  );


  bp_be_top_vaddr_width_p39_paddr_width_p22_asid_width_p10_branch_metadata_fwd_width_p36_core_els_p1_trace_p0_num_cce_p1_num_lce_p2_lce_assoc_p8_lce_sets_p64_cce_block_size_in_bytes_p64
  be
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .fe_queue_i(be_fe_queue),
    .fe_queue_v_i(be_fe_queue_v),
    .fe_queue_ready_o(be_fe_queue_ready),
    .fe_queue_clr_o(fe_queue_clr[0]),
    .fe_queue_dequeue_o(fe_queue_dequeue[0]),
    .fe_queue_rollback_o(fe_queue_rollback[0]),
    .fe_cmd_o(be_fe_cmd),
    .fe_cmd_v_o(be_fe_cmd_v[0]),
    .fe_cmd_ready_i(be_fe_cmd_ready[0]),
    .lce_req_o(lce_req_o[193:97]),
    .lce_req_v_o(lce_req_v_o[1]),
    .lce_req_ready_i(lce_req_ready_i[1]),
    .lce_resp_o(lce_resp_o[51:26]),
    .lce_resp_v_o(lce_resp_v_o[1]),
    .lce_resp_ready_i(lce_resp_ready_i[1]),
    .lce_data_resp_o(lce_data_resp_o[1073:537]),
    .lce_data_resp_v_o(lce_data_resp_v_o[1]),
    .lce_data_resp_ready_i(lce_data_resp_ready_i[1]),
    .lce_cmd_i(lce_cmd_i[71:36]),
    .lce_cmd_v_i(lce_cmd_v_i[1]),
    .lce_cmd_ready_o(lce_cmd_ready_o[1]),
    .lce_data_cmd_i(lce_data_cmd_i[1035:518]),
    .lce_data_cmd_v_i(lce_data_cmd_v_i[1]),
    .lce_data_cmd_ready_o(lce_data_cmd_ready_o[1]),
    .lce_data_cmd_o(lce_data_cmd_o[1035:518]),
    .lce_data_cmd_v_o(lce_data_cmd_v_o[1]),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_i[1]),
    .proc_cfg_i(proc_cfg_i),
    .cmt_rd_w_v_o(cmt_rd_w_v_o),
    .cmt_rd_addr_o(cmt_rd_addr_o),
    .cmt_mem_w_v_o(cmt_mem_w_v_o),
    .cmt_mem_addr_o(cmt_mem_addr_o),
    .cmt_mem_op_o(cmt_mem_op_o),
    .cmt_data_o(cmt_data_o)
  );


endmodule



module bsg_mem_p38
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [37:0] w_data_i;
  input [0:0] r_addr_i;
  output [37:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [37:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  reg [75:0] mem;
  assign r_data_o[37] = (N3)? mem[37] :
                        (N0)? mem[75] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[36] = (N3)? mem[36] :
                        (N0)? mem[74] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] :
                        (N0)? mem[73] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] :
                        (N0)? mem[72] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] :
                        (N0)? mem[71] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] :
                        (N0)? mem[70] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] :
                        (N0)? mem[69] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] :
                        (N0)? mem[68] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] :
                        (N0)? mem[67] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] :
                        (N0)? mem[66] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] :
                        (N0)? mem[65] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] :
                        (N0)? mem[64] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] :
                        (N0)? mem[63] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] :
                        (N0)? mem[62] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] :
                        (N0)? mem[61] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] :
                        (N0)? mem[60] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] :
                        (N0)? mem[59] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] :
                        (N0)? mem[58] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] :
                        (N0)? mem[57] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] :
                        (N0)? mem[56] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] :
                        (N0)? mem[55] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] :
                        (N0)? mem[54] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] :
                        (N0)? mem[53] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] :
                        (N0)? mem[52] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] :
                        (N0)? mem[51] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] :
                        (N0)? mem[50] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] :
                        (N0)? mem[49] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] :
                        (N0)? mem[48] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] :
                       (N0)? mem[47] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] :
                       (N0)? mem[46] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] :
                       (N0)? mem[45] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] :
                       (N0)? mem[44] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] :
                       (N0)? mem[43] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] :
                       (N0)? mem[42] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] :
                       (N0)? mem[41] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] :
                       (N0)? mem[40] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] :
                       (N0)? mem[39] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] :
                       (N0)? mem[38] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } :
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      { mem[75:38] } <= { w_data_i[37:0] };
    end
    if(N7) begin
      { mem[37:0] } <= { w_data_i[37:0] };
    end
  end


endmodule



module bsg_mem_1r1w_width_p38_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [37:0] w_data_i;
  input [0:0] r_addr_i;
  output [37:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [37:0] r_data_o;

  bsg_mem_p38
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p38
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [37:0] data_i;
  output [37:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [37:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p38_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 :
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 :
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 :
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 :
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 :
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 :
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end
    if(N9) begin
      tail_r <= N10;
    end
    if(N11) begin
      head_r <= N12;
    end
  end


endmodule



module bsg_mesh_router_dor_decoder_x_cord_width_p1_y_cord_width_p1_dirs_lp5_XY_order_p0
(
  clk_i,
  v_i,
  x_dirs_i,
  y_dirs_i,
  my_x_i,
  my_y_i,
  req_o
);

  input [4:0] v_i;
  input [4:0] x_dirs_i;
  input [4:0] y_dirs_i;
  input [0:0] my_x_i;
  input [0:0] my_y_i;
  output [24:0] req_o;
  input clk_i;
  wire [24:0] req_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,y_gt_0,x_lt_0,
  y_lt_0,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,
  N37,N38,N39,N40,N41,N42;
  wire [4:0] x_eq,y_eq,x_gt;
  wire [4:3] y_gt;
  wire [4:2] x_lt;
  wire [4:4] y_lt;
  assign req_o[12] = 1'b0;
  assign req_o[6] = 1'b0;
  assign req_o[24] = 1'b0;
  assign req_o[18] = 1'b0;
  assign req_o[14] = 1'b0;
  assign req_o[13] = 1'b0;
  assign req_o[9] = 1'b0;
  assign req_o[8] = 1'b0;
  assign N0 = x_dirs_i[0] ^ my_x_i[0];
  assign x_eq[0] = ~N0;
  assign N1 = y_dirs_i[0] ^ my_y_i[0];
  assign y_eq[0] = ~N1;
  assign x_gt[0] = x_dirs_i[0] & N2;
  assign N2 = ~my_x_i[0];
  assign y_gt_0 = y_dirs_i[0] & N3;
  assign N3 = ~my_y_i[0];
  assign N4 = x_dirs_i[1] ^ my_x_i[0];
  assign x_eq[1] = ~N4;
  assign N5 = y_dirs_i[1] ^ my_y_i[0];
  assign y_eq[1] = ~N5;
  assign x_gt[1] = x_dirs_i[1] & N6;
  assign N6 = ~my_x_i[0];
  assign N7 = x_dirs_i[2] ^ my_x_i[0];
  assign x_eq[2] = ~N7;
  assign N8 = y_dirs_i[2] ^ my_y_i[0];
  assign y_eq[2] = ~N8;
  assign x_gt[2] = x_dirs_i[2] & N9;
  assign N9 = ~my_x_i[0];
  assign N10 = x_dirs_i[3] ^ my_x_i[0];
  assign x_eq[3] = ~N10;
  assign N11 = y_dirs_i[3] ^ my_y_i[0];
  assign y_eq[3] = ~N11;
  assign x_gt[3] = x_dirs_i[3] & N12;
  assign N12 = ~my_x_i[0];
  assign y_gt[3] = y_dirs_i[3] & N13;
  assign N13 = ~my_y_i[0];
  assign N14 = x_dirs_i[4] ^ my_x_i[0];
  assign x_eq[4] = ~N14;
  assign N15 = y_dirs_i[4] ^ my_y_i[0];
  assign y_eq[4] = ~N15;
  assign x_gt[4] = x_dirs_i[4] & N16;
  assign N16 = ~my_x_i[0];
  assign y_gt[4] = y_dirs_i[4] & N17;
  assign N17 = ~my_y_i[0];
  assign x_lt_0 = N18 & N19;
  assign N18 = ~x_gt[0];
  assign N19 = ~x_eq[0];
  assign y_lt_0 = N20 & N21;
  assign N20 = ~y_gt_0;
  assign N21 = ~y_eq[0];
  assign x_lt[2] = N22 & N23;
  assign N22 = ~x_gt[2];
  assign N23 = ~x_eq[2];
  assign x_lt[3] = N24 & N25;
  assign N24 = ~x_gt[3];
  assign N25 = ~x_eq[3];
  assign x_lt[4] = N26 & N27;
  assign N26 = ~x_gt[4];
  assign N27 = ~x_eq[4];
  assign y_lt[4] = N28 & N29;
  assign N28 = ~y_gt[4];
  assign N29 = ~y_eq[4];
  assign req_o[16] = N30 & x_lt[3];
  assign N30 = v_i[3] & y_eq[3];
  assign req_o[17] = N31 & x_gt[3];
  assign N31 = v_i[3] & y_eq[3];
  assign req_o[21] = N32 & x_lt[4];
  assign N32 = v_i[4] & y_eq[4];
  assign req_o[22] = N33 & x_gt[4];
  assign N33 = v_i[4] & y_eq[4];
  assign req_o[19] = v_i[3] & y_gt[3];
  assign req_o[23] = v_i[4] & y_lt[4];
  assign req_o[7] = N34 & x_gt[1];
  assign N34 = v_i[1] & y_eq[1];
  assign req_o[11] = N35 & x_lt[2];
  assign N35 = v_i[2] & y_eq[2];
  assign req_o[4] = v_i[0] & y_gt_0;
  assign req_o[3] = v_i[0] & y_lt_0;
  assign req_o[0] = N36 & y_eq[0];
  assign N36 = v_i[0] & x_eq[0];
  assign req_o[2] = N37 & x_gt[0];
  assign N37 = v_i[0] & y_eq[0];
  assign req_o[1] = N38 & x_lt_0;
  assign N38 = v_i[0] & y_eq[0];
  assign req_o[5] = N39 & y_eq[1];
  assign N39 = v_i[1] & x_eq[1];
  assign req_o[10] = N40 & y_eq[2];
  assign N40 = v_i[2] & x_eq[2];
  assign req_o[15] = N41 & y_eq[3];
  assign N41 = v_i[3] & x_eq[3];
  assign req_o[20] = N42 & y_eq[4];
  assign N42 = v_i[4] & x_eq[4];

endmodule



module bsg_round_robin_arb_inputs_p4
(
  clk_i,
  reset_i,
  grants_en_i,
  reqs_i,
  grants_o,
  sel_one_hot_o,
  v_o,
  tag_o,
  yumi_i
);

  input [3:0] reqs_i;
  output [3:0] grants_o;
  output [3:0] sel_one_hot_o;
  output [1:0] tag_o;
  input clk_i;
  input reset_i;
  input grants_en_i;
  input yumi_i;
  output v_o;
  wire [3:0] grants_o,sel_one_hot_o;
  wire [1:0] tag_o;
  wire v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,
  N101,N102,N103;
  reg [1:0] last_r;
  assign N79 = N0 & N1 & (N2 & N3);
  assign N0 = ~reqs_i[1];
  assign N1 = ~reqs_i[2];
  assign N2 = ~reqs_i[0];
  assign N3 = ~reqs_i[3];
  assign N80 = reqs_i[1] & N4 & N5;
  assign N4 = ~last_r[0];
  assign N5 = ~last_r[1];
  assign N81 = N6 & reqs_i[2] & (N7 & N8);
  assign N6 = ~reqs_i[1];
  assign N7 = ~last_r[0];
  assign N8 = ~last_r[1];
  assign N82 = N9 & N10 & (reqs_i[3] & N11) & N12;
  assign N9 = ~reqs_i[1];
  assign N10 = ~reqs_i[2];
  assign N11 = ~last_r[0];
  assign N12 = ~last_r[1];
  assign N13 = N17 & N18;
  assign N14 = N13 & reqs_i[0];
  assign N15 = N14 & N19;
  assign N16 = N15 & N20;
  assign N83 = N16 & N21;
  assign N17 = ~reqs_i[1];
  assign N18 = ~reqs_i[2];
  assign N19 = ~reqs_i[3];
  assign N20 = ~last_r[0];
  assign N21 = ~last_r[1];
  assign N84 = reqs_i[2] & last_r[0] & N22;
  assign N22 = ~last_r[1];
  assign N85 = N23 & reqs_i[3] & (last_r[0] & N24);
  assign N23 = ~reqs_i[2];
  assign N24 = ~last_r[1];
  assign N86 = N25 & reqs_i[0] & (N26 & last_r[0]) & N27;
  assign N25 = ~reqs_i[2];
  assign N26 = ~reqs_i[3];
  assign N27 = ~last_r[1];
  assign N28 = reqs_i[1] & N32;
  assign N29 = N28 & N33;
  assign N30 = N29 & N34;
  assign N31 = N30 & last_r[0];
  assign N87 = N31 & N35;
  assign N32 = ~reqs_i[2];
  assign N33 = ~reqs_i[0];
  assign N34 = ~reqs_i[3];
  assign N35 = ~last_r[1];
  assign N88 = reqs_i[3] & N36 & last_r[1];
  assign N36 = ~last_r[0];
  assign N89 = reqs_i[0] & N37 & (N38 & last_r[1]);
  assign N37 = ~reqs_i[3];
  assign N38 = ~last_r[0];
  assign N90 = reqs_i[1] & N39 & (N40 & N41) & last_r[1];
  assign N39 = ~reqs_i[0];
  assign N40 = ~reqs_i[3];
  assign N41 = ~last_r[0];
  assign N42 = N46 & reqs_i[2];
  assign N43 = N42 & N47;
  assign N44 = N43 & N48;
  assign N45 = N44 & N49;
  assign N91 = N45 & last_r[1];
  assign N46 = ~reqs_i[1];
  assign N47 = ~reqs_i[0];
  assign N48 = ~reqs_i[3];
  assign N49 = ~last_r[0];
  assign N92 = reqs_i[0] & last_r[0] & last_r[1];
  assign N93 = reqs_i[1] & N50 & (last_r[0] & last_r[1]);
  assign N50 = ~reqs_i[0];
  assign N94 = N51 & reqs_i[2] & (N52 & last_r[0]) & last_r[1];
  assign N51 = ~reqs_i[1];
  assign N52 = ~reqs_i[0];
  assign N53 = N57 & N58;
  assign N54 = N53 & N59;
  assign N55 = N54 & reqs_i[3];
  assign N56 = N55 & last_r[0];
  assign N95 = N56 & last_r[1];
  assign N57 = ~reqs_i[1];
  assign N58 = ~reqs_i[2];
  assign N59 = ~reqs_i[0];
  assign sel_one_hot_o = (N60)? { 1'b0, 1'b0, 1'b0, 1'b0 } :
                         (N61)? { 1'b0, 1'b0, 1'b1, 1'b0 } :
                         (N62)? { 1'b0, 1'b1, 1'b0, 1'b0 } :
                         (N63)? { 1'b1, 1'b0, 1'b0, 1'b0 } :
                         (N64)? { 1'b0, 1'b0, 1'b0, 1'b1 } :
                         (N65)? { 1'b0, 1'b1, 1'b0, 1'b0 } :
                         (N66)? { 1'b1, 1'b0, 1'b0, 1'b0 } :
                         (N67)? { 1'b0, 1'b0, 1'b0, 1'b1 } :
                         (N68)? { 1'b0, 1'b0, 1'b1, 1'b0 } :
                         (N69)? { 1'b1, 1'b0, 1'b0, 1'b0 } :
                         (N70)? { 1'b0, 1'b0, 1'b0, 1'b1 } :
                         (N71)? { 1'b0, 1'b0, 1'b1, 1'b0 } :
                         (N72)? { 1'b0, 1'b1, 1'b0, 1'b0 } :
                         (N73)? { 1'b0, 1'b0, 1'b0, 1'b1 } :
                         (N74)? { 1'b0, 1'b0, 1'b1, 1'b0 } :
                         (N75)? { 1'b0, 1'b1, 1'b0, 1'b0 } :
                         (N76)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N60 = N79;
  assign N61 = N80;
  assign N62 = N81;
  assign N63 = N82;
  assign N64 = N83;
  assign N65 = N84;
  assign N66 = N85;
  assign N67 = N86;
  assign N68 = N87;
  assign N69 = N88;
  assign N70 = N89;
  assign N71 = N90;
  assign N72 = N91;
  assign N73 = N92;
  assign N74 = N93;
  assign N75 = N94;
  assign N76 = N95;
  assign tag_o = (N60)? { 1'b0, 1'b0 } :
                 (N61)? { 1'b0, 1'b1 } :
                 (N62)? { 1'b1, 1'b0 } :
                 (N63)? { 1'b1, 1'b1 } :
                 (N64)? { 1'b0, 1'b0 } :
                 (N65)? { 1'b1, 1'b0 } :
                 (N66)? { 1'b1, 1'b1 } :
                 (N67)? { 1'b0, 1'b0 } :
                 (N68)? { 1'b0, 1'b1 } :
                 (N69)? { 1'b1, 1'b1 } :
                 (N70)? { 1'b0, 1'b0 } :
                 (N71)? { 1'b0, 1'b1 } :
                 (N72)? { 1'b1, 1'b0 } :
                 (N73)? { 1'b0, 1'b0 } :
                 (N74)? { 1'b0, 1'b1 } :
                 (N75)? { 1'b1, 1'b0 } :
                 (N76)? { 1'b1, 1'b1 } : 1'b0;
  assign { N99, N98 } = (N77)? { 1'b0, 1'b0 } :
                        (N78)? tag_o : 1'b0;
  assign N77 = reset_i;
  assign N78 = N97;
  assign grants_o[3] = sel_one_hot_o[3] & grants_en_i;
  assign grants_o[2] = sel_one_hot_o[2] & grants_en_i;
  assign grants_o[1] = sel_one_hot_o[1] & grants_en_i;
  assign grants_o[0] = sel_one_hot_o[0] & grants_en_i;
  assign v_o = N103 | reqs_i[0];
  assign N103 = N102 | reqs_i[1];
  assign N102 = reqs_i[3] | reqs_i[2];
  assign N96 = ~yumi_i;
  assign N97 = ~reset_i;
  assign N100 = N96 & N97;
  assign N101 = ~N100;

  always @(posedge clk_i) begin
    if(N101) begin
      { last_r[1:0] } <= { N99, N98 };
    end
  end


endmodule



module bsg_mux_one_hot_width_p38_els_p4
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [151:0] data_i;
  input [3:0] sel_one_hot_i;
  output [37:0] data_o;
  wire [37:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75;
  wire [151:0] data_masked;
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[1];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[1];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[1];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[1];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[1];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[1];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[1];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[1];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[1];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[1];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[1];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[1];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[1];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[1];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[1];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[1];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[1];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[1];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[1];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[1];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[1];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[1];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[1];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[1];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[1];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[2];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[2];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[2];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[2];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[2];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[2];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[2];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[2];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[2];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[2];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[2];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[2];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[2];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[2];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[2];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[2];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[2];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[2];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[2];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[2];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[2];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[2];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[2];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[2];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[2];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[2];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[2];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[2];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[2];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[2];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[2];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[2];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[2];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[2];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[2];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[2];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[2];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[2];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[3];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[3];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[3];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[3];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[3];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[3];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[3];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[3];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[3];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[3];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[3];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[3];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[3];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[3];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[3];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[3];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[3];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[3];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[3];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[3];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[3];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[3];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[3];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[3];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[3];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[3];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[3];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[3];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[3];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[3];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[3];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[3];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[3];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[3];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[3];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[3];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[3];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[3];
  assign data_o[0] = N1 | data_masked[0];
  assign N1 = N0 | data_masked[38];
  assign N0 = data_masked[114] | data_masked[76];
  assign data_o[1] = N3 | data_masked[1];
  assign N3 = N2 | data_masked[39];
  assign N2 = data_masked[115] | data_masked[77];
  assign data_o[2] = N5 | data_masked[2];
  assign N5 = N4 | data_masked[40];
  assign N4 = data_masked[116] | data_masked[78];
  assign data_o[3] = N7 | data_masked[3];
  assign N7 = N6 | data_masked[41];
  assign N6 = data_masked[117] | data_masked[79];
  assign data_o[4] = N9 | data_masked[4];
  assign N9 = N8 | data_masked[42];
  assign N8 = data_masked[118] | data_masked[80];
  assign data_o[5] = N11 | data_masked[5];
  assign N11 = N10 | data_masked[43];
  assign N10 = data_masked[119] | data_masked[81];
  assign data_o[6] = N13 | data_masked[6];
  assign N13 = N12 | data_masked[44];
  assign N12 = data_masked[120] | data_masked[82];
  assign data_o[7] = N15 | data_masked[7];
  assign N15 = N14 | data_masked[45];
  assign N14 = data_masked[121] | data_masked[83];
  assign data_o[8] = N17 | data_masked[8];
  assign N17 = N16 | data_masked[46];
  assign N16 = data_masked[122] | data_masked[84];
  assign data_o[9] = N19 | data_masked[9];
  assign N19 = N18 | data_masked[47];
  assign N18 = data_masked[123] | data_masked[85];
  assign data_o[10] = N21 | data_masked[10];
  assign N21 = N20 | data_masked[48];
  assign N20 = data_masked[124] | data_masked[86];
  assign data_o[11] = N23 | data_masked[11];
  assign N23 = N22 | data_masked[49];
  assign N22 = data_masked[125] | data_masked[87];
  assign data_o[12] = N25 | data_masked[12];
  assign N25 = N24 | data_masked[50];
  assign N24 = data_masked[126] | data_masked[88];
  assign data_o[13] = N27 | data_masked[13];
  assign N27 = N26 | data_masked[51];
  assign N26 = data_masked[127] | data_masked[89];
  assign data_o[14] = N29 | data_masked[14];
  assign N29 = N28 | data_masked[52];
  assign N28 = data_masked[128] | data_masked[90];
  assign data_o[15] = N31 | data_masked[15];
  assign N31 = N30 | data_masked[53];
  assign N30 = data_masked[129] | data_masked[91];
  assign data_o[16] = N33 | data_masked[16];
  assign N33 = N32 | data_masked[54];
  assign N32 = data_masked[130] | data_masked[92];
  assign data_o[17] = N35 | data_masked[17];
  assign N35 = N34 | data_masked[55];
  assign N34 = data_masked[131] | data_masked[93];
  assign data_o[18] = N37 | data_masked[18];
  assign N37 = N36 | data_masked[56];
  assign N36 = data_masked[132] | data_masked[94];
  assign data_o[19] = N39 | data_masked[19];
  assign N39 = N38 | data_masked[57];
  assign N38 = data_masked[133] | data_masked[95];
  assign data_o[20] = N41 | data_masked[20];
  assign N41 = N40 | data_masked[58];
  assign N40 = data_masked[134] | data_masked[96];
  assign data_o[21] = N43 | data_masked[21];
  assign N43 = N42 | data_masked[59];
  assign N42 = data_masked[135] | data_masked[97];
  assign data_o[22] = N45 | data_masked[22];
  assign N45 = N44 | data_masked[60];
  assign N44 = data_masked[136] | data_masked[98];
  assign data_o[23] = N47 | data_masked[23];
  assign N47 = N46 | data_masked[61];
  assign N46 = data_masked[137] | data_masked[99];
  assign data_o[24] = N49 | data_masked[24];
  assign N49 = N48 | data_masked[62];
  assign N48 = data_masked[138] | data_masked[100];
  assign data_o[25] = N51 | data_masked[25];
  assign N51 = N50 | data_masked[63];
  assign N50 = data_masked[139] | data_masked[101];
  assign data_o[26] = N53 | data_masked[26];
  assign N53 = N52 | data_masked[64];
  assign N52 = data_masked[140] | data_masked[102];
  assign data_o[27] = N55 | data_masked[27];
  assign N55 = N54 | data_masked[65];
  assign N54 = data_masked[141] | data_masked[103];
  assign data_o[28] = N57 | data_masked[28];
  assign N57 = N56 | data_masked[66];
  assign N56 = data_masked[142] | data_masked[104];
  assign data_o[29] = N59 | data_masked[29];
  assign N59 = N58 | data_masked[67];
  assign N58 = data_masked[143] | data_masked[105];
  assign data_o[30] = N61 | data_masked[30];
  assign N61 = N60 | data_masked[68];
  assign N60 = data_masked[144] | data_masked[106];
  assign data_o[31] = N63 | data_masked[31];
  assign N63 = N62 | data_masked[69];
  assign N62 = data_masked[145] | data_masked[107];
  assign data_o[32] = N65 | data_masked[32];
  assign N65 = N64 | data_masked[70];
  assign N64 = data_masked[146] | data_masked[108];
  assign data_o[33] = N67 | data_masked[33];
  assign N67 = N66 | data_masked[71];
  assign N66 = data_masked[147] | data_masked[109];
  assign data_o[34] = N69 | data_masked[34];
  assign N69 = N68 | data_masked[72];
  assign N68 = data_masked[148] | data_masked[110];
  assign data_o[35] = N71 | data_masked[35];
  assign N71 = N70 | data_masked[73];
  assign N70 = data_masked[149] | data_masked[111];
  assign data_o[36] = N73 | data_masked[36];
  assign N73 = N72 | data_masked[74];
  assign N72 = data_masked[150] | data_masked[112];
  assign data_o[37] = N75 | data_masked[37];
  assign N75 = N74 | data_masked[75];
  assign N74 = data_masked[151] | data_masked[113];

endmodule



module bsg_round_robin_arb_inputs_p2
(
  clk_i,
  reset_i,
  grants_en_i,
  reqs_i,
  grants_o,
  sel_one_hot_o,
  v_o,
  tag_o,
  yumi_i
);

  input [1:0] reqs_i;
  output [1:0] grants_o;
  output [1:0] sel_one_hot_o;
  output [0:0] tag_o;
  input clk_i;
  input reset_i;
  input grants_en_i;
  input yumi_i;
  output v_o;
  wire [1:0] grants_o,sel_one_hot_o;
  wire [0:0] tag_o;
  wire v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22;
  reg [0:0] last_r;
  assign N13 = N0 & N1;
  assign N0 = ~reqs_i[1];
  assign N1 = ~reqs_i[0];
  assign N14 = reqs_i[1] & N2;
  assign N2 = ~last_r[0];
  assign N15 = N3 & reqs_i[0] & N4;
  assign N3 = ~reqs_i[1];
  assign N4 = ~last_r[0];
  assign N16 = reqs_i[0] & last_r[0];
  assign N17 = reqs_i[1] & N5 & last_r[0];
  assign N5 = ~reqs_i[0];
  assign sel_one_hot_o = (N6)? { 1'b0, 1'b0 } :
                         (N7)? { 1'b1, 1'b0 } :
                         (N8)? { 1'b0, 1'b1 } :
                         (N9)? { 1'b0, 1'b1 } :
                         (N10)? { 1'b1, 1'b0 } : 1'b0;
  assign N6 = N13;
  assign N7 = N14;
  assign N8 = N15;
  assign N9 = N16;
  assign N10 = N17;
  assign tag_o[0] = (N6)? 1'b0 :
                    (N7)? 1'b1 :
                    (N8)? 1'b0 :
                    (N9)? 1'b0 :
                    (N10)? 1'b1 : 1'b0;
  assign N20 = (N11)? 1'b0 :
               (N12)? tag_o[0] : 1'b0;
  assign N11 = reset_i;
  assign N12 = N19;
  assign grants_o[1] = sel_one_hot_o[1] & grants_en_i;
  assign grants_o[0] = sel_one_hot_o[0] & grants_en_i;
  assign v_o = reqs_i[1] | reqs_i[0];
  assign N18 = ~yumi_i;
  assign N19 = ~reset_i;
  assign N21 = N18 & N19;
  assign N22 = ~N21;

  always @(posedge clk_i) begin
    if(N22) begin
      { last_r[0:0] } <= { N20 };
    end
  end


endmodule



module bsg_mux_one_hot_width_p38_els_p2
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [75:0] data_i;
  input [1:0] sel_one_hot_i;
  output [37:0] data_o;
  wire [37:0] data_o;
  wire [75:0] data_masked;
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[1];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[1];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[1];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[1];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[1];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[1];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[1];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[1];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[1];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[1];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[1];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[1];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[1];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[1];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[1];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[1];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[1];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[1];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[1];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[1];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[1];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[1];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[1];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[1];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[1];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[1];
  assign data_o[0] = data_masked[38] | data_masked[0];
  assign data_o[1] = data_masked[39] | data_masked[1];
  assign data_o[2] = data_masked[40] | data_masked[2];
  assign data_o[3] = data_masked[41] | data_masked[3];
  assign data_o[4] = data_masked[42] | data_masked[4];
  assign data_o[5] = data_masked[43] | data_masked[5];
  assign data_o[6] = data_masked[44] | data_masked[6];
  assign data_o[7] = data_masked[45] | data_masked[7];
  assign data_o[8] = data_masked[46] | data_masked[8];
  assign data_o[9] = data_masked[47] | data_masked[9];
  assign data_o[10] = data_masked[48] | data_masked[10];
  assign data_o[11] = data_masked[49] | data_masked[11];
  assign data_o[12] = data_masked[50] | data_masked[12];
  assign data_o[13] = data_masked[51] | data_masked[13];
  assign data_o[14] = data_masked[52] | data_masked[14];
  assign data_o[15] = data_masked[53] | data_masked[15];
  assign data_o[16] = data_masked[54] | data_masked[16];
  assign data_o[17] = data_masked[55] | data_masked[17];
  assign data_o[18] = data_masked[56] | data_masked[18];
  assign data_o[19] = data_masked[57] | data_masked[19];
  assign data_o[20] = data_masked[58] | data_masked[20];
  assign data_o[21] = data_masked[59] | data_masked[21];
  assign data_o[22] = data_masked[60] | data_masked[22];
  assign data_o[23] = data_masked[61] | data_masked[23];
  assign data_o[24] = data_masked[62] | data_masked[24];
  assign data_o[25] = data_masked[63] | data_masked[25];
  assign data_o[26] = data_masked[64] | data_masked[26];
  assign data_o[27] = data_masked[65] | data_masked[27];
  assign data_o[28] = data_masked[66] | data_masked[28];
  assign data_o[29] = data_masked[67] | data_masked[29];
  assign data_o[30] = data_masked[68] | data_masked[30];
  assign data_o[31] = data_masked[69] | data_masked[31];
  assign data_o[32] = data_masked[70] | data_masked[32];
  assign data_o[33] = data_masked[71] | data_masked[33];
  assign data_o[34] = data_masked[72] | data_masked[34];
  assign data_o[35] = data_masked[73] | data_masked[35];
  assign data_o[36] = data_masked[74] | data_masked[36];
  assign data_o[37] = data_masked[75] | data_masked[37];

endmodule



module bsg_round_robin_arb_inputs_p5
(
  clk_i,
  reset_i,
  grants_en_i,
  reqs_i,
  grants_o,
  sel_one_hot_o,
  v_o,
  tag_o,
  yumi_i
);

  input [4:0] reqs_i;
  output [4:0] grants_o;
  output [4:0] sel_one_hot_o;
  output [2:0] tag_o;
  input clk_i;
  input reset_i;
  input grants_en_i;
  input yumi_i;
  output v_o;
  wire [4:0] grants_o,sel_one_hot_o;
  wire [2:0] tag_o;
  wire v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,
  N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,
  N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,
  N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,
  N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,
  N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,
  N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195;
  reg [2:0] last_r;
  assign N21 = N19 & N88;
  assign N22 = N21 & N37;
  assign N23 = N22 & N20;
  assign N27 = N24 & N25;
  assign N28 = N26 & reqs_i[1];
  assign N29 = N27 & N28;
  assign N31 = N24 & N25;
  assign N32 = N26 & reqs_i[2];
  assign N33 = N31 & N32;
  assign N34 = N33 & N30;
  assign N35 = N24 & N25;
  assign N36 = N26 & reqs_i[3];
  assign N37 = N56 & N30;
  assign N38 = N35 & N36;
  assign N39 = N38 & N37;
  assign N40 = last_r[2] | last_r[1];
  assign N41 = last_r[0] | N19;
  assign N42 = N40 | N41;
  assign N43 = N63 | reqs_i[1];
  assign N44 = N42 | N43;
  assign N46 = last_r[2] | last_r[1];
  assign N47 = last_r[0] | reqs_i[4];
  assign N48 = reqs_i[1] | N20;
  assign N49 = N46 | N47;
  assign N50 = N63 | N48;
  assign N51 = N49 | N50;
  assign N53 = N24 & N25;
  assign N54 = last_r[0] & reqs_i[2];
  assign N55 = N53 & N54;
  assign N57 = N24 & N25;
  assign N58 = last_r[0] & reqs_i[3];
  assign N59 = N57 & N58;
  assign N60 = N59 & N56;
  assign N61 = last_r[2] | last_r[1];
  assign N62 = N26 | N19;
  assign N63 = reqs_i[3] | reqs_i[2];
  assign N64 = N61 | N62;
  assign N65 = N64 | N63;
  assign N67 = N24 & N25;
  assign N68 = last_r[0] & N19;
  assign N69 = N88 & N56;
  assign N70 = N67 & N68;
  assign N71 = N69 & reqs_i[0];
  assign N72 = N70 & N71;
  assign N73 = last_r[2] | last_r[1];
  assign N74 = N26 | reqs_i[4];
  assign N75 = N30 | reqs_i[0];
  assign N76 = N73 | N74;
  assign N77 = N63 | N75;
  assign N78 = N76 | N77;
  assign N80 = N24 & last_r[1];
  assign N81 = N26 & reqs_i[3];
  assign N82 = N80 & N81;
  assign N83 = last_r[2] | N25;
  assign N84 = last_r[0] | N19;
  assign N85 = N83 | N84;
  assign N86 = N85 | reqs_i[3];
  assign N89 = N24 & last_r[1];
  assign N90 = N26 & N19;
  assign N91 = N88 & reqs_i[0];
  assign N92 = N89 & N90;
  assign N93 = N92 & N91;
  assign N94 = N24 & last_r[1];
  assign N95 = N26 & N19;
  assign N96 = N88 & reqs_i[1];
  assign N97 = N94 & N95;
  assign N98 = N96 & N20;
  assign N99 = N97 & N98;
  assign N100 = last_r[2] | N25;
  assign N101 = last_r[0] | reqs_i[4];
  assign N102 = reqs_i[3] | N56;
  assign N103 = reqs_i[1] | reqs_i[0];
  assign N104 = N100 | N101;
  assign N105 = N102 | N103;
  assign N106 = N104 | N105;
  assign N108 = last_r[2] | N25;
  assign N109 = N26 | N19;
  assign N110 = N108 | N109;
  assign N112 = N24 & last_r[1];
  assign N113 = last_r[0] & N19;
  assign N114 = N112 & N113;
  assign N115 = N114 & reqs_i[0];
  assign N116 = N24 & last_r[1];
  assign N117 = last_r[0] & N19;
  assign N118 = reqs_i[1] & N20;
  assign N119 = N116 & N117;
  assign N120 = N119 & N118;
  assign N121 = N24 & last_r[1];
  assign N122 = last_r[0] & N19;
  assign N123 = reqs_i[2] & N30;
  assign N124 = N121 & N122;
  assign N125 = N123 & N20;
  assign N126 = N124 & N125;
  assign N127 = last_r[2] | N25;
  assign N128 = N26 | reqs_i[4];
  assign N129 = N88 | reqs_i[2];
  assign N130 = N127 | N128;
  assign N131 = N129 | N103;
  assign N132 = N130 | N131;
  assign N134 = last_r[2] & N25;
  assign N135 = N26 & reqs_i[0];
  assign N136 = N134 & N135;
  assign N137 = last_r[2] & N25;
  assign N138 = N26 & reqs_i[1];
  assign N139 = N137 & N138;
  assign N140 = N139 & N20;
  assign N141 = last_r[2] & N25;
  assign N142 = N26 & reqs_i[2];
  assign N143 = N30 & N20;
  assign N144 = N141 & N142;
  assign N145 = N144 & N143;
  assign N146 = last_r[2] & N25;
  assign N147 = N26 & reqs_i[3];
  assign N148 = N146 & N147;
  assign N149 = N37 & N20;
  assign N150 = N148 & N149;
  assign N151 = N24 | last_r[1];
  assign N152 = last_r[0] | N19;
  assign N153 = N151 | N152;
  assign N154 = N63 | N103;
  assign N155 = N153 | N154;
  assign N157 = last_r[2] & last_r[0];
  assign N158 = N157 & reqs_i[2];
  assign N159 = last_r[2] & last_r[0];
  assign N160 = N159 & reqs_i[3];
  assign N161 = last_r[2] & last_r[0];
  assign N162 = N161 & reqs_i[4];
  assign N163 = last_r[2] & last_r[0];
  assign N164 = N163 & reqs_i[0];
  assign N165 = last_r[2] & last_r[0];
  assign N166 = N165 & reqs_i[1];
  assign N167 = last_r[2] & last_r[1];
  assign N168 = N167 & reqs_i[3];
  assign N169 = last_r[2] & last_r[1];
  assign N170 = N169 & reqs_i[4];
  assign N171 = last_r[2] & last_r[1];
  assign N172 = N171 & reqs_i[0];
  assign N173 = last_r[2] & last_r[1];
  assign N174 = N173 & reqs_i[1];
  assign N175 = last_r[2] & last_r[1];
  assign N176 = N175 & reqs_i[2];
  assign sel_one_hot_o = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                         (N1)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } :
                         (N2)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } :
                         (N3)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } :
                         (N45)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } :
                         (N52)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } :
                         (N4)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } :
                         (N5)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } :
                         (N66)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } :
                         (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } :
                         (N79)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } :
                         (N7)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } :
                         (N87)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } :
                         (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } :
                         (N9)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } :
                         (N107)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } :
                         (N111)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } :
                         (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } :
                         (N11)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } :
                         (N12)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } :
                         (N133)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } :
                         (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } :
                         (N14)? { 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } :
                         (N15)? { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } :
                         (N16)? { 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } :
                         (N156)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N23;
  assign N1 = N29;
  assign N2 = N34;
  assign N3 = N39;
  assign N4 = N55;
  assign N5 = N60;
  assign N6 = N72;
  assign N7 = N82;
  assign N8 = N93;
  assign N9 = N99;
  assign N10 = N115;
  assign N11 = N120;
  assign N12 = N126;
  assign N13 = N136;
  assign N14 = N140;
  assign N15 = N145;
  assign N16 = N150;
  assign tag_o = (N0)? { 1'b0, 1'b0, 1'b0 } :
                 (N1)? { 1'b0, 1'b0, 1'b1 } :
                 (N2)? { 1'b0, 1'b1, 1'b0 } :
                 (N3)? { 1'b0, 1'b1, 1'b1 } :
                 (N45)? { 1'b1, 1'b0, 1'b0 } :
                 (N52)? { 1'b0, 1'b0, 1'b0 } :
                 (N4)? { 1'b0, 1'b1, 1'b0 } :
                 (N5)? { 1'b0, 1'b1, 1'b1 } :
                 (N66)? { 1'b1, 1'b0, 1'b0 } :
                 (N6)? { 1'b0, 1'b0, 1'b0 } :
                 (N79)? { 1'b0, 1'b0, 1'b1 } :
                 (N7)? { 1'b0, 1'b1, 1'b1 } :
                 (N87)? { 1'b1, 1'b0, 1'b0 } :
                 (N8)? { 1'b0, 1'b0, 1'b0 } :
                 (N9)? { 1'b0, 1'b0, 1'b1 } :
                 (N107)? { 1'b0, 1'b1, 1'b0 } :
                 (N111)? { 1'b1, 1'b0, 1'b0 } :
                 (N10)? { 1'b0, 1'b0, 1'b0 } :
                 (N11)? { 1'b0, 1'b0, 1'b1 } :
                 (N12)? { 1'b0, 1'b1, 1'b0 } :
                 (N133)? { 1'b0, 1'b1, 1'b1 } :
                 (N13)? { 1'b0, 1'b0, 1'b0 } :
                 (N14)? { 1'b0, 1'b0, 1'b1 } :
                 (N15)? { 1'b0, 1'b1, 1'b0 } :
                 (N16)? { 1'b0, 1'b1, 1'b1 } :
                 (N156)? { 1'b1, 1'b0, 1'b0 } :
                 (N177)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N182, N181, N180 } = (N17)? { 1'b0, 1'b0, 1'b0 } :
                                (N18)? tag_o : 1'b0;
  assign N17 = reset_i;
  assign N18 = N179;
  assign N19 = ~reqs_i[4];
  assign N20 = ~reqs_i[0];
  assign N24 = ~last_r[2];
  assign N25 = ~last_r[1];
  assign N26 = ~last_r[0];
  assign N30 = ~reqs_i[1];
  assign N45 = ~N44;
  assign N52 = ~N51;
  assign N56 = ~reqs_i[2];
  assign N66 = ~N65;
  assign N79 = ~N78;
  assign N87 = ~N86;
  assign N88 = ~reqs_i[3];
  assign N107 = ~N106;
  assign N111 = ~N110;
  assign N133 = ~N132;
  assign N156 = ~N155;
  assign N177 = N158 | N192;
  assign N192 = N160 | N191;
  assign N191 = N162 | N190;
  assign N190 = N164 | N189;
  assign N189 = N166 | N188;
  assign N188 = N168 | N187;
  assign N187 = N170 | N186;
  assign N186 = N172 | N185;
  assign N185 = N174 | N176;
  assign grants_o[4] = sel_one_hot_o[4] & grants_en_i;
  assign grants_o[3] = sel_one_hot_o[3] & grants_en_i;
  assign grants_o[2] = sel_one_hot_o[2] & grants_en_i;
  assign grants_o[1] = sel_one_hot_o[1] & grants_en_i;
  assign grants_o[0] = sel_one_hot_o[0] & grants_en_i;
  assign v_o = N195 | reqs_i[0];
  assign N195 = N194 | reqs_i[1];
  assign N194 = N193 | reqs_i[2];
  assign N193 = reqs_i[4] | reqs_i[3];
  assign N178 = ~yumi_i;
  assign N179 = ~reset_i;
  assign N183 = N178 & N179;
  assign N184 = ~N183;

  always @(posedge clk_i) begin
    if(N184) begin
      { last_r[2:0] } <= { N182, N181, N180 };
    end
  end


endmodule



module bsg_mux_one_hot_width_p38_els_p5
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [189:0] data_i;
  input [4:0] sel_one_hot_i;
  output [37:0] data_o;
  wire [37:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113;
  wire [189:0] data_masked;
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[1];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[1];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[1];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[1];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[1];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[1];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[1];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[1];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[1];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[1];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[1];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[1];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[1];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[1];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[1];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[1];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[1];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[1];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[1];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[1];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[1];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[1];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[1];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[1];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[1];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[2];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[2];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[2];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[2];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[2];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[2];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[2];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[2];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[2];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[2];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[2];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[2];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[2];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[2];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[2];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[2];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[2];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[2];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[2];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[2];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[2];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[2];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[2];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[2];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[2];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[2];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[2];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[2];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[2];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[2];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[2];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[2];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[2];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[2];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[2];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[2];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[2];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[2];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[3];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[3];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[3];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[3];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[3];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[3];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[3];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[3];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[3];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[3];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[3];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[3];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[3];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[3];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[3];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[3];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[3];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[3];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[3];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[3];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[3];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[3];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[3];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[3];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[3];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[3];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[3];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[3];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[3];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[3];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[3];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[3];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[3];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[3];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[3];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[3];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[3];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[3];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[4];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[4];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[4];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[4];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[4];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[4];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[4];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[4];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[4];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[4];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[4];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[4];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[4];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[4];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[4];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[4];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[4];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[4];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[4];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[4];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[4];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[4];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[4];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[4];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[4];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[4];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[4];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[4];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[4];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[4];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[4];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[4];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[4];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[4];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[4];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[4];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[4];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[4];
  assign data_o[0] = N2 | data_masked[0];
  assign N2 = N1 | data_masked[38];
  assign N1 = N0 | data_masked[76];
  assign N0 = data_masked[152] | data_masked[114];
  assign data_o[1] = N5 | data_masked[1];
  assign N5 = N4 | data_masked[39];
  assign N4 = N3 | data_masked[77];
  assign N3 = data_masked[153] | data_masked[115];
  assign data_o[2] = N8 | data_masked[2];
  assign N8 = N7 | data_masked[40];
  assign N7 = N6 | data_masked[78];
  assign N6 = data_masked[154] | data_masked[116];
  assign data_o[3] = N11 | data_masked[3];
  assign N11 = N10 | data_masked[41];
  assign N10 = N9 | data_masked[79];
  assign N9 = data_masked[155] | data_masked[117];
  assign data_o[4] = N14 | data_masked[4];
  assign N14 = N13 | data_masked[42];
  assign N13 = N12 | data_masked[80];
  assign N12 = data_masked[156] | data_masked[118];
  assign data_o[5] = N17 | data_masked[5];
  assign N17 = N16 | data_masked[43];
  assign N16 = N15 | data_masked[81];
  assign N15 = data_masked[157] | data_masked[119];
  assign data_o[6] = N20 | data_masked[6];
  assign N20 = N19 | data_masked[44];
  assign N19 = N18 | data_masked[82];
  assign N18 = data_masked[158] | data_masked[120];
  assign data_o[7] = N23 | data_masked[7];
  assign N23 = N22 | data_masked[45];
  assign N22 = N21 | data_masked[83];
  assign N21 = data_masked[159] | data_masked[121];
  assign data_o[8] = N26 | data_masked[8];
  assign N26 = N25 | data_masked[46];
  assign N25 = N24 | data_masked[84];
  assign N24 = data_masked[160] | data_masked[122];
  assign data_o[9] = N29 | data_masked[9];
  assign N29 = N28 | data_masked[47];
  assign N28 = N27 | data_masked[85];
  assign N27 = data_masked[161] | data_masked[123];
  assign data_o[10] = N32 | data_masked[10];
  assign N32 = N31 | data_masked[48];
  assign N31 = N30 | data_masked[86];
  assign N30 = data_masked[162] | data_masked[124];
  assign data_o[11] = N35 | data_masked[11];
  assign N35 = N34 | data_masked[49];
  assign N34 = N33 | data_masked[87];
  assign N33 = data_masked[163] | data_masked[125];
  assign data_o[12] = N38 | data_masked[12];
  assign N38 = N37 | data_masked[50];
  assign N37 = N36 | data_masked[88];
  assign N36 = data_masked[164] | data_masked[126];
  assign data_o[13] = N41 | data_masked[13];
  assign N41 = N40 | data_masked[51];
  assign N40 = N39 | data_masked[89];
  assign N39 = data_masked[165] | data_masked[127];
  assign data_o[14] = N44 | data_masked[14];
  assign N44 = N43 | data_masked[52];
  assign N43 = N42 | data_masked[90];
  assign N42 = data_masked[166] | data_masked[128];
  assign data_o[15] = N47 | data_masked[15];
  assign N47 = N46 | data_masked[53];
  assign N46 = N45 | data_masked[91];
  assign N45 = data_masked[167] | data_masked[129];
  assign data_o[16] = N50 | data_masked[16];
  assign N50 = N49 | data_masked[54];
  assign N49 = N48 | data_masked[92];
  assign N48 = data_masked[168] | data_masked[130];
  assign data_o[17] = N53 | data_masked[17];
  assign N53 = N52 | data_masked[55];
  assign N52 = N51 | data_masked[93];
  assign N51 = data_masked[169] | data_masked[131];
  assign data_o[18] = N56 | data_masked[18];
  assign N56 = N55 | data_masked[56];
  assign N55 = N54 | data_masked[94];
  assign N54 = data_masked[170] | data_masked[132];
  assign data_o[19] = N59 | data_masked[19];
  assign N59 = N58 | data_masked[57];
  assign N58 = N57 | data_masked[95];
  assign N57 = data_masked[171] | data_masked[133];
  assign data_o[20] = N62 | data_masked[20];
  assign N62 = N61 | data_masked[58];
  assign N61 = N60 | data_masked[96];
  assign N60 = data_masked[172] | data_masked[134];
  assign data_o[21] = N65 | data_masked[21];
  assign N65 = N64 | data_masked[59];
  assign N64 = N63 | data_masked[97];
  assign N63 = data_masked[173] | data_masked[135];
  assign data_o[22] = N68 | data_masked[22];
  assign N68 = N67 | data_masked[60];
  assign N67 = N66 | data_masked[98];
  assign N66 = data_masked[174] | data_masked[136];
  assign data_o[23] = N71 | data_masked[23];
  assign N71 = N70 | data_masked[61];
  assign N70 = N69 | data_masked[99];
  assign N69 = data_masked[175] | data_masked[137];
  assign data_o[24] = N74 | data_masked[24];
  assign N74 = N73 | data_masked[62];
  assign N73 = N72 | data_masked[100];
  assign N72 = data_masked[176] | data_masked[138];
  assign data_o[25] = N77 | data_masked[25];
  assign N77 = N76 | data_masked[63];
  assign N76 = N75 | data_masked[101];
  assign N75 = data_masked[177] | data_masked[139];
  assign data_o[26] = N80 | data_masked[26];
  assign N80 = N79 | data_masked[64];
  assign N79 = N78 | data_masked[102];
  assign N78 = data_masked[178] | data_masked[140];
  assign data_o[27] = N83 | data_masked[27];
  assign N83 = N82 | data_masked[65];
  assign N82 = N81 | data_masked[103];
  assign N81 = data_masked[179] | data_masked[141];
  assign data_o[28] = N86 | data_masked[28];
  assign N86 = N85 | data_masked[66];
  assign N85 = N84 | data_masked[104];
  assign N84 = data_masked[180] | data_masked[142];
  assign data_o[29] = N89 | data_masked[29];
  assign N89 = N88 | data_masked[67];
  assign N88 = N87 | data_masked[105];
  assign N87 = data_masked[181] | data_masked[143];
  assign data_o[30] = N92 | data_masked[30];
  assign N92 = N91 | data_masked[68];
  assign N91 = N90 | data_masked[106];
  assign N90 = data_masked[182] | data_masked[144];
  assign data_o[31] = N95 | data_masked[31];
  assign N95 = N94 | data_masked[69];
  assign N94 = N93 | data_masked[107];
  assign N93 = data_masked[183] | data_masked[145];
  assign data_o[32] = N98 | data_masked[32];
  assign N98 = N97 | data_masked[70];
  assign N97 = N96 | data_masked[108];
  assign N96 = data_masked[184] | data_masked[146];
  assign data_o[33] = N101 | data_masked[33];
  assign N101 = N100 | data_masked[71];
  assign N100 = N99 | data_masked[109];
  assign N99 = data_masked[185] | data_masked[147];
  assign data_o[34] = N104 | data_masked[34];
  assign N104 = N103 | data_masked[72];
  assign N103 = N102 | data_masked[110];
  assign N102 = data_masked[186] | data_masked[148];
  assign data_o[35] = N107 | data_masked[35];
  assign N107 = N106 | data_masked[73];
  assign N106 = N105 | data_masked[111];
  assign N105 = data_masked[187] | data_masked[149];
  assign data_o[36] = N110 | data_masked[36];
  assign N110 = N109 | data_masked[74];
  assign N109 = N108 | data_masked[112];
  assign N108 = data_masked[188] | data_masked[150];
  assign data_o[37] = N113 | data_masked[37];
  assign N113 = N112 | data_masked[75];
  assign N112 = N111 | data_masked[113];
  assign N111 = data_masked[189] | data_masked[151];

endmodule



module bsg_mesh_router_38_1_1_0_0a_0
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  yumi_o,
  ready_i,
  data_o,
  v_o,
  my_x_i,
  my_y_i
);

  input [189:0] data_i;
  input [4:0] v_i;
  output [4:0] yumi_o;
  input [4:0] ready_i;
  output [189:0] data_o;
  output [4:0] v_o;
  input [0:0] my_x_i;
  input [0:0] my_y_i;
  input clk_i;
  input reset_i;
  wire [4:0] yumi_o,v_o;
  wire [189:0] data_o;
  wire n_3_net_,W_sel_e,W_sel_p,W_sel_n,W_sel_s,W_gnt_e,W_gnt_p,W_gnt_n,W_gnt_s,
  n_9_net_,E_sel_w,E_sel_p,E_sel_n,E_sel_s,E_gnt_w,E_gnt_p,E_gnt_n,E_gnt_s,n_15_net_,
  N_sel_s,N_sel_p,N_gnt_s,N_gnt_p,n_21_net_,S_sel_n,S_sel_p,S_gnt_n,S_gnt_p,n_27_net_,
  P_sel_s,P_sel_n,P_sel_e,P_sel_w,P_sel_p,P_gnt_s,P_gnt_n,P_gnt_e,P_gnt_w,P_gnt_p,
  N0,N1,N2,N3,N4,N5,N6,SV2V_UNCONNECTED_1,SV2V_UNCONNECTED_2,
  SV2V_UNCONNECTED_3,SV2V_UNCONNECTED_4,SV2V_UNCONNECTED_5,SV2V_UNCONNECTED_6,
  SV2V_UNCONNECTED_7,SV2V_UNCONNECTED_8,SV2V_UNCONNECTED_9;
  wire [24:0] req;

  bsg_mesh_router_dor_decoder_x_cord_width_p1_y_cord_width_p1_dirs_lp5_XY_order_p0
  dor_decoder
  (
    .clk_i(clk_i),
    .v_i({ v_i[4:4], 1'b0, v_i[2:2], 1'b0, v_i[0:0] }),
    .x_dirs_i({ data_i[152:152], data_i[114:114], data_i[76:76], data_i[38:38], data_i[0:0] }),
    .y_dirs_i({ data_i[153:153], data_i[115:115], data_i[77:77], data_i[39:39], data_i[1:1] }),
    .my_x_i(my_x_i[0]),
    .my_y_i(my_y_i[0]),
    .req_o(req)
  );


  bsg_round_robin_arb_inputs_p4
  genblk2_west_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ req[11:11], req[1:1], req[16:16], req[21:21] }),
    .grants_o({ W_gnt_e, W_gnt_p, W_gnt_n, W_gnt_s }),
    .sel_one_hot_o({ W_sel_e, W_sel_p, W_sel_n, W_sel_s }),
    .v_o(v_o[1]),
    .tag_o({ SV2V_UNCONNECTED_1, SV2V_UNCONNECTED_2 }),
    .yumi_i(n_3_net_)
  );


  bsg_mux_one_hot_width_p38_els_p4
  genblk2_mux_data_west
  (
    .data_i({ data_i[37:0], data_i[113:76], data_i[151:114], data_i[189:152] }),
    .sel_one_hot_i({ W_sel_p, W_sel_e, W_sel_n, W_sel_s }),
    .data_o(data_o[75:38])
  );


  bsg_round_robin_arb_inputs_p4
  genblk3_east_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[2]),
    .reqs_i({ req[7:7], req[2:2], req[17:17], req[22:22] }),
    .grants_o({ E_gnt_w, E_gnt_p, E_gnt_n, E_gnt_s }),
    .sel_one_hot_o({ E_sel_w, E_sel_p, E_sel_n, E_sel_s }),
    .v_o(v_o[2]),
    .tag_o({ SV2V_UNCONNECTED_3, SV2V_UNCONNECTED_4 }),
    .yumi_i(n_9_net_)
  );


  bsg_mux_one_hot_width_p38_els_p4
  genblk3_mux_data_east
  (
    .data_i({ data_i[37:0], data_i[75:38], data_i[151:114], data_i[189:152] }),
    .sel_one_hot_i({ E_sel_p, E_sel_w, E_sel_n, E_sel_s }),
    .data_o(data_o[113:76])
  );


  bsg_round_robin_arb_inputs_p2
  genblk4_north_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ req[23:23], req[3:3] }),
    .grants_o({ N_gnt_s, N_gnt_p }),
    .sel_one_hot_o({ N_sel_s, N_sel_p }),
    .v_o(v_o[3]),
    .tag_o(SV2V_UNCONNECTED_5),
    .yumi_i(n_15_net_)
  );


  bsg_mux_one_hot_width_p38_els_p2
  genblk4_mux_data_north
  (
    .data_i({ data_i[37:0], data_i[189:152] }),
    .sel_one_hot_i({ N_sel_p, N_sel_s }),
    .data_o(data_o[151:114])
  );


  bsg_round_robin_arb_inputs_p2
  genblk5_south_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[4]),
    .reqs_i({ req[19:19], req[4:4] }),
    .grants_o({ S_gnt_n, S_gnt_p }),
    .sel_one_hot_o({ S_sel_n, S_sel_p }),
    .v_o(v_o[4]),
    .tag_o(SV2V_UNCONNECTED_6),
    .yumi_i(n_21_net_)
  );


  bsg_mux_one_hot_width_p38_els_p2
  genblk5_mux_data_south
  (
    .data_i({ data_i[37:0], data_i[151:114] }),
    .sel_one_hot_i({ S_sel_p, S_sel_n }),
    .data_o(data_o[189:152])
  );


  bsg_round_robin_arb_inputs_p5
  proc_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[0]),
    .reqs_i({ req[20:20], req[15:15], req[10:10], req[5:5], req[0:0] }),
    .grants_o({ P_gnt_s, P_gnt_n, P_gnt_e, P_gnt_w, P_gnt_p }),
    .sel_one_hot_o({ P_sel_s, P_sel_n, P_sel_e, P_sel_w, P_sel_p }),
    .v_o(v_o[0]),
    .tag_o({ SV2V_UNCONNECTED_7, SV2V_UNCONNECTED_8, SV2V_UNCONNECTED_9 }),
    .yumi_i(n_27_net_)
  );


  bsg_mux_one_hot_width_p38_els_p5
  mux_data_proc
  (
    .data_i({ data_i[37:0], data_i[113:76], data_i[189:152], data_i[75:38], data_i[151:114] }),
    .sel_one_hot_i({ P_sel_p, P_sel_e, P_sel_s, P_sel_w, P_sel_n }),
    .data_o(data_o[37:0])
  );

  assign n_3_net_ = v_o[1] & 1'b1;
  assign n_9_net_ = v_o[2] & ready_i[2];
  assign n_15_net_ = v_o[3] & 1'b1;
  assign n_21_net_ = v_o[4] & ready_i[4];
  assign n_27_net_ = v_o[0] & ready_i[0];
  assign yumi_o[0] = N2 | W_gnt_p;
  assign N2 = N1 | P_gnt_p;
  assign N1 = N0 | S_gnt_p;
  assign N0 = E_gnt_p | N_gnt_p;
  assign yumi_o[1] = E_gnt_w | P_gnt_w;
  assign yumi_o[2] = W_gnt_e | P_gnt_e;
  assign yumi_o[3] = N4 | P_gnt_n;
  assign N4 = N3 | E_gnt_n;
  assign N3 = S_gnt_n | W_gnt_n;
  assign yumi_o[4] = N6 | P_gnt_s;
  assign N6 = N5 | E_gnt_s;
  assign N5 = N_gnt_s | W_gnt_s;

endmodule



module bsg_mesh_router_buffered_38_1_1_0_5_0a_0_40_00
(
  clk_i,
  reset_i,
  link_i,
  link_o,
  my_x_i,
  my_y_i
);

  input [199:0] link_i;
  output [199:0] link_o;
  input [0:0] my_x_i;
  input [0:0] my_y_i;
  input clk_i;
  input reset_i;
  wire [199:0] link_o;
  wire fifo_valid_2,fifo_valid_0,fifo_data_4__37_,fifo_data_4__36_,fifo_data_4__35_,
  fifo_data_4__34_,fifo_data_4__33_,fifo_data_4__32_,fifo_data_4__31_,
  fifo_data_4__30_,fifo_data_4__29_,fifo_data_4__28_,fifo_data_4__27_,fifo_data_4__26_,
  fifo_data_4__25_,fifo_data_4__24_,fifo_data_4__23_,fifo_data_4__22_,fifo_data_4__21_,
  fifo_data_4__20_,fifo_data_4__19_,fifo_data_4__18_,fifo_data_4__17_,fifo_data_4__16_,
  fifo_data_4__15_,fifo_data_4__14_,fifo_data_4__13_,fifo_data_4__12_,
  fifo_data_4__11_,fifo_data_4__10_,fifo_data_4__9_,fifo_data_4__8_,fifo_data_4__7_,
  fifo_data_4__6_,fifo_data_4__5_,fifo_data_4__4_,fifo_data_4__3_,fifo_data_4__2_,
  fifo_data_4__1_,fifo_data_4__0_,fifo_data_2__37_,fifo_data_2__36_,fifo_data_2__35_,
  fifo_data_2__34_,fifo_data_2__33_,fifo_data_2__32_,fifo_data_2__31_,fifo_data_2__30_,
  fifo_data_2__29_,fifo_data_2__28_,fifo_data_2__27_,fifo_data_2__26_,
  fifo_data_2__25_,fifo_data_2__24_,fifo_data_2__23_,fifo_data_2__22_,fifo_data_2__21_,
  fifo_data_2__20_,fifo_data_2__19_,fifo_data_2__18_,fifo_data_2__17_,fifo_data_2__16_,
  fifo_data_2__15_,fifo_data_2__14_,fifo_data_2__13_,fifo_data_2__12_,
  fifo_data_2__11_,fifo_data_2__10_,fifo_data_2__9_,fifo_data_2__8_,fifo_data_2__7_,
  fifo_data_2__6_,fifo_data_2__5_,fifo_data_2__4_,fifo_data_2__3_,fifo_data_2__2_,
  fifo_data_2__1_,fifo_data_2__0_,fifo_data_0__37_,fifo_data_0__36_,fifo_data_0__35_,
  fifo_data_0__34_,fifo_data_0__33_,fifo_data_0__32_,fifo_data_0__31_,fifo_data_0__30_,
  fifo_data_0__29_,fifo_data_0__28_,fifo_data_0__27_,fifo_data_0__26_,fifo_data_0__25_,
  fifo_data_0__24_,fifo_data_0__23_,fifo_data_0__22_,fifo_data_0__21_,
  fifo_data_0__20_,fifo_data_0__19_,fifo_data_0__18_,fifo_data_0__17_,fifo_data_0__16_,
  fifo_data_0__15_,fifo_data_0__14_,fifo_data_0__13_,fifo_data_0__12_,fifo_data_0__11_,
  fifo_data_0__10_,fifo_data_0__9_,fifo_data_0__8_,fifo_data_0__7_,fifo_data_0__6_,
  fifo_data_0__5_,fifo_data_0__4_,fifo_data_0__3_,fifo_data_0__2_,fifo_data_0__1_,
  fifo_data_0__0_;
  wire [4:4] fifo_valid;
  wire [4:0] fifo_yumi;
  assign link_o[78] = 1'b0;
  assign link_o[158] = 1'b0;

  bsg_two_fifo_width_p38
  rof_0__fi_twofer
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(link_o[38]),
    .data_i(link_i[37:0]),
    .v_i(link_i[39]),
    .v_o(fifo_valid_0),
    .data_o({ fifo_data_0__37_, fifo_data_0__36_, fifo_data_0__35_, fifo_data_0__34_, fifo_data_0__33_, fifo_data_0__32_, fifo_data_0__31_, fifo_data_0__30_, fifo_data_0__29_, fifo_data_0__28_, fifo_data_0__27_, fifo_data_0__26_, fifo_data_0__25_, fifo_data_0__24_, fifo_data_0__23_, fifo_data_0__22_, fifo_data_0__21_, fifo_data_0__20_, fifo_data_0__19_, fifo_data_0__18_, fifo_data_0__17_, fifo_data_0__16_, fifo_data_0__15_, fifo_data_0__14_, fifo_data_0__13_, fifo_data_0__12_, fifo_data_0__11_, fifo_data_0__10_, fifo_data_0__9_, fifo_data_0__8_, fifo_data_0__7_, fifo_data_0__6_, fifo_data_0__5_, fifo_data_0__4_, fifo_data_0__3_, fifo_data_0__2_, fifo_data_0__1_, fifo_data_0__0_ }),
    .yumi_i(fifo_yumi[0])
  );


  bsg_two_fifo_width_p38
  rof_2__fi_twofer
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(link_o[118]),
    .data_i(link_i[117:80]),
    .v_i(link_i[119]),
    .v_o(fifo_valid_2),
    .data_o({ fifo_data_2__37_, fifo_data_2__36_, fifo_data_2__35_, fifo_data_2__34_, fifo_data_2__33_, fifo_data_2__32_, fifo_data_2__31_, fifo_data_2__30_, fifo_data_2__29_, fifo_data_2__28_, fifo_data_2__27_, fifo_data_2__26_, fifo_data_2__25_, fifo_data_2__24_, fifo_data_2__23_, fifo_data_2__22_, fifo_data_2__21_, fifo_data_2__20_, fifo_data_2__19_, fifo_data_2__18_, fifo_data_2__17_, fifo_data_2__16_, fifo_data_2__15_, fifo_data_2__14_, fifo_data_2__13_, fifo_data_2__12_, fifo_data_2__11_, fifo_data_2__10_, fifo_data_2__9_, fifo_data_2__8_, fifo_data_2__7_, fifo_data_2__6_, fifo_data_2__5_, fifo_data_2__4_, fifo_data_2__3_, fifo_data_2__2_, fifo_data_2__1_, fifo_data_2__0_ }),
    .yumi_i(fifo_yumi[2])
  );


  bsg_two_fifo_width_p38
  rof_4__fi_twofer
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(link_o[198]),
    .data_i(link_i[197:160]),
    .v_i(link_i[199]),
    .v_o(fifo_valid[4]),
    .data_o({ fifo_data_4__37_, fifo_data_4__36_, fifo_data_4__35_, fifo_data_4__34_, fifo_data_4__33_, fifo_data_4__32_, fifo_data_4__31_, fifo_data_4__30_, fifo_data_4__29_, fifo_data_4__28_, fifo_data_4__27_, fifo_data_4__26_, fifo_data_4__25_, fifo_data_4__24_, fifo_data_4__23_, fifo_data_4__22_, fifo_data_4__21_, fifo_data_4__20_, fifo_data_4__19_, fifo_data_4__18_, fifo_data_4__17_, fifo_data_4__16_, fifo_data_4__15_, fifo_data_4__14_, fifo_data_4__13_, fifo_data_4__12_, fifo_data_4__11_, fifo_data_4__10_, fifo_data_4__9_, fifo_data_4__8_, fifo_data_4__7_, fifo_data_4__6_, fifo_data_4__5_, fifo_data_4__4_, fifo_data_4__3_, fifo_data_4__2_, fifo_data_4__1_, fifo_data_4__0_ }),
    .yumi_i(fifo_yumi[4])
  );


  bsg_mesh_router_38_1_1_0_0a_0
  bmr
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ fifo_data_4__37_, fifo_data_4__36_, fifo_data_4__35_, fifo_data_4__34_, fifo_data_4__33_, fifo_data_4__32_, fifo_data_4__31_, fifo_data_4__30_, fifo_data_4__29_, fifo_data_4__28_, fifo_data_4__27_, fifo_data_4__26_, fifo_data_4__25_, fifo_data_4__24_, fifo_data_4__23_, fifo_data_4__22_, fifo_data_4__21_, fifo_data_4__20_, fifo_data_4__19_, fifo_data_4__18_, fifo_data_4__17_, fifo_data_4__16_, fifo_data_4__15_, fifo_data_4__14_, fifo_data_4__13_, fifo_data_4__12_, fifo_data_4__11_, fifo_data_4__10_, fifo_data_4__9_, fifo_data_4__8_, fifo_data_4__7_, fifo_data_4__6_, fifo_data_4__5_, fifo_data_4__4_, fifo_data_4__3_, fifo_data_4__2_, fifo_data_4__1_, fifo_data_4__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_2__37_, fifo_data_2__36_, fifo_data_2__35_, fifo_data_2__34_, fifo_data_2__33_, fifo_data_2__32_, fifo_data_2__31_, fifo_data_2__30_, fifo_data_2__29_, fifo_data_2__28_, fifo_data_2__27_, fifo_data_2__26_, fifo_data_2__25_, fifo_data_2__24_, fifo_data_2__23_, fifo_data_2__22_, fifo_data_2__21_, fifo_data_2__20_, fifo_data_2__19_, fifo_data_2__18_, fifo_data_2__17_, fifo_data_2__16_, fifo_data_2__15_, fifo_data_2__14_, fifo_data_2__13_, fifo_data_2__12_, fifo_data_2__11_, fifo_data_2__10_, fifo_data_2__9_, fifo_data_2__8_, fifo_data_2__7_, fifo_data_2__6_, fifo_data_2__5_, fifo_data_2__4_, fifo_data_2__3_, fifo_data_2__2_, fifo_data_2__1_, fifo_data_2__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_0__37_, fifo_data_0__36_, fifo_data_0__35_, fifo_data_0__34_, fifo_data_0__33_, fifo_data_0__32_, fifo_data_0__31_, fifo_data_0__30_, fifo_data_0__29_, fifo_data_0__28_, fifo_data_0__27_, fifo_data_0__26_, fifo_data_0__25_, fifo_data_0__24_, fifo_data_0__23_, fifo_data_0__22_, fifo_data_0__21_, fifo_data_0__20_, fifo_data_0__19_, fifo_data_0__18_, fifo_data_0__17_, fifo_data_0__16_, fifo_data_0__15_, fifo_data_0__14_, fifo_data_0__13_, fifo_data_0__12_, fifo_data_0__11_, fifo_data_0__10_, fifo_data_0__9_, fifo_data_0__8_, fifo_data_0__7_, fifo_data_0__6_, fifo_data_0__5_, fifo_data_0__4_, fifo_data_0__3_, fifo_data_0__2_, fifo_data_0__1_, fifo_data_0__0_ }),
    .v_i({ fifo_valid[4:4], 1'b0, fifo_valid_2, 1'b0, fifo_valid_0 }),
    .yumi_o(fifo_yumi),
    .ready_i({ link_i[198:198], link_i[158:158], link_i[118:118], link_i[78:78], link_i[38:38] }),
    .data_o({ link_o[197:160], link_o[157:120], link_o[117:80], link_o[77:40], link_o[37:0] }),
    .v_o({ link_o[199:199], link_o[159:159], link_o[119:119], link_o[79:79], link_o[39:39] }),
    .my_x_i(my_x_i[0]),
    .my_y_i(my_y_i[0])
  );


endmodule



module bsg_mesh_router_38_1_1_0_1c_0
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  yumi_o,
  ready_i,
  data_o,
  v_o,
  my_x_i,
  my_y_i
);

  input [189:0] data_i;
  input [4:0] v_i;
  output [4:0] yumi_o;
  input [4:0] ready_i;
  output [189:0] data_o;
  output [4:0] v_o;
  input [0:0] my_x_i;
  input [0:0] my_y_i;
  input clk_i;
  input reset_i;
  wire [4:0] yumi_o,v_o;
  wire [189:0] data_o;
  wire n_3_net_,W_sel_e,W_sel_p,W_sel_n,W_sel_s,W_gnt_e,W_gnt_p,W_gnt_n,W_gnt_s,
  n_9_net_,E_sel_w,E_sel_p,E_sel_n,E_sel_s,E_gnt_w,E_gnt_p,E_gnt_n,E_gnt_s,n_15_net_,
  N_sel_s,N_sel_p,N_gnt_s,N_gnt_p,n_21_net_,S_sel_n,S_sel_p,S_gnt_n,S_gnt_p,n_27_net_,
  P_sel_s,P_sel_n,P_sel_e,P_sel_w,P_sel_p,P_gnt_s,P_gnt_n,P_gnt_e,P_gnt_w,P_gnt_p,
  N0,N1,N2,N3,N4,N5,N6,SV2V_UNCONNECTED_1,SV2V_UNCONNECTED_2,
  SV2V_UNCONNECTED_3,SV2V_UNCONNECTED_4,SV2V_UNCONNECTED_5,SV2V_UNCONNECTED_6,
  SV2V_UNCONNECTED_7,SV2V_UNCONNECTED_8,SV2V_UNCONNECTED_9;
  wire [24:0] req;

  bsg_mesh_router_dor_decoder_x_cord_width_p1_y_cord_width_p1_dirs_lp5_XY_order_p0
  dor_decoder
  (
    .clk_i(clk_i),
    .v_i({ 1'b0, 1'b0, 1'b0, v_i[1:0] }),
    .x_dirs_i({ data_i[152:152], data_i[114:114], data_i[76:76], data_i[38:38], data_i[0:0] }),
    .y_dirs_i({ data_i[153:153], data_i[115:115], data_i[77:77], data_i[39:39], data_i[1:1] }),
    .my_x_i(my_x_i[0]),
    .my_y_i(my_y_i[0]),
    .req_o(req)
  );


  bsg_round_robin_arb_inputs_p4
  genblk2_west_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[1]),
    .reqs_i({ req[11:11], req[1:1], req[16:16], req[21:21] }),
    .grants_o({ W_gnt_e, W_gnt_p, W_gnt_n, W_gnt_s }),
    .sel_one_hot_o({ W_sel_e, W_sel_p, W_sel_n, W_sel_s }),
    .v_o(v_o[1]),
    .tag_o({ SV2V_UNCONNECTED_1, SV2V_UNCONNECTED_2 }),
    .yumi_i(n_3_net_)
  );


  bsg_mux_one_hot_width_p38_els_p4
  genblk2_mux_data_west
  (
    .data_i({ data_i[37:0], data_i[113:76], data_i[151:114], data_i[189:152] }),
    .sel_one_hot_i({ W_sel_p, W_sel_e, W_sel_n, W_sel_s }),
    .data_o(data_o[75:38])
  );


  bsg_round_robin_arb_inputs_p4
  genblk3_east_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ req[7:7], req[2:2], req[17:17], req[22:22] }),
    .grants_o({ E_gnt_w, E_gnt_p, E_gnt_n, E_gnt_s }),
    .sel_one_hot_o({ E_sel_w, E_sel_p, E_sel_n, E_sel_s }),
    .v_o(v_o[2]),
    .tag_o({ SV2V_UNCONNECTED_3, SV2V_UNCONNECTED_4 }),
    .yumi_i(n_9_net_)
  );


  bsg_mux_one_hot_width_p38_els_p4
  genblk3_mux_data_east
  (
    .data_i({ data_i[37:0], data_i[75:38], data_i[151:114], data_i[189:152] }),
    .sel_one_hot_i({ E_sel_p, E_sel_w, E_sel_n, E_sel_s }),
    .data_o(data_o[113:76])
  );


  bsg_round_robin_arb_inputs_p2
  genblk4_north_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ req[23:23], req[3:3] }),
    .grants_o({ N_gnt_s, N_gnt_p }),
    .sel_one_hot_o({ N_sel_s, N_sel_p }),
    .v_o(v_o[3]),
    .tag_o(SV2V_UNCONNECTED_5),
    .yumi_i(n_15_net_)
  );


  bsg_mux_one_hot_width_p38_els_p2
  genblk4_mux_data_north
  (
    .data_i({ data_i[37:0], data_i[189:152] }),
    .sel_one_hot_i({ N_sel_p, N_sel_s }),
    .data_o(data_o[151:114])
  );


  bsg_round_robin_arb_inputs_p2
  genblk5_south_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ req[19:19], req[4:4] }),
    .grants_o({ S_gnt_n, S_gnt_p }),
    .sel_one_hot_o({ S_sel_n, S_sel_p }),
    .v_o(v_o[4]),
    .tag_o(SV2V_UNCONNECTED_6),
    .yumi_i(n_21_net_)
  );


  bsg_mux_one_hot_width_p38_els_p2
  genblk5_mux_data_south
  (
    .data_i({ data_i[37:0], data_i[151:114] }),
    .sel_one_hot_i({ S_sel_p, S_sel_n }),
    .data_o(data_o[189:152])
  );


  bsg_round_robin_arb_inputs_p5
  proc_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[0]),
    .reqs_i({ req[20:20], req[15:15], req[10:10], req[5:5], req[0:0] }),
    .grants_o({ P_gnt_s, P_gnt_n, P_gnt_e, P_gnt_w, P_gnt_p }),
    .sel_one_hot_o({ P_sel_s, P_sel_n, P_sel_e, P_sel_w, P_sel_p }),
    .v_o(v_o[0]),
    .tag_o({ SV2V_UNCONNECTED_7, SV2V_UNCONNECTED_8, SV2V_UNCONNECTED_9 }),
    .yumi_i(n_27_net_)
  );


  bsg_mux_one_hot_width_p38_els_p5
  mux_data_proc
  (
    .data_i({ data_i[37:0], data_i[113:76], data_i[189:152], data_i[75:38], data_i[151:114] }),
    .sel_one_hot_i({ P_sel_p, P_sel_e, P_sel_s, P_sel_w, P_sel_n }),
    .data_o(data_o[37:0])
  );

  assign n_3_net_ = v_o[1] & ready_i[1];
  assign n_9_net_ = v_o[2] & 1'b1;
  assign n_15_net_ = v_o[3] & 1'b1;
  assign n_21_net_ = v_o[4] & 1'b1;
  assign n_27_net_ = v_o[0] & ready_i[0];
  assign yumi_o[0] = N2 | W_gnt_p;
  assign N2 = N1 | P_gnt_p;
  assign N1 = N0 | S_gnt_p;
  assign N0 = E_gnt_p | N_gnt_p;
  assign yumi_o[1] = E_gnt_w | P_gnt_w;
  assign yumi_o[2] = W_gnt_e | P_gnt_e;
  assign yumi_o[3] = N4 | P_gnt_n;
  assign N4 = N3 | E_gnt_n;
  assign N3 = S_gnt_n | W_gnt_n;
  assign yumi_o[4] = N6 | P_gnt_s;
  assign N6 = N5 | E_gnt_s;
  assign N5 = N_gnt_s | W_gnt_s;

endmodule



module bsg_mesh_router_buffered_38_1_1_0_5_1c_0_40_00
(
  clk_i,
  reset_i,
  link_i,
  link_o,
  my_x_i,
  my_y_i
);

  input [199:0] link_i;
  output [199:0] link_o;
  input [0:0] my_x_i;
  input [0:0] my_y_i;
  input clk_i;
  input reset_i;
  wire [199:0] link_o;
  wire fifo_data_1__37_,fifo_data_1__36_,fifo_data_1__35_,fifo_data_1__34_,
  fifo_data_1__33_,fifo_data_1__32_,fifo_data_1__31_,fifo_data_1__30_,fifo_data_1__29_,
  fifo_data_1__28_,fifo_data_1__27_,fifo_data_1__26_,fifo_data_1__25_,fifo_data_1__24_,
  fifo_data_1__23_,fifo_data_1__22_,fifo_data_1__21_,fifo_data_1__20_,
  fifo_data_1__19_,fifo_data_1__18_,fifo_data_1__17_,fifo_data_1__16_,fifo_data_1__15_,
  fifo_data_1__14_,fifo_data_1__13_,fifo_data_1__12_,fifo_data_1__11_,fifo_data_1__10_,
  fifo_data_1__9_,fifo_data_1__8_,fifo_data_1__7_,fifo_data_1__6_,fifo_data_1__5_,
  fifo_data_1__4_,fifo_data_1__3_,fifo_data_1__2_,fifo_data_1__1_,fifo_data_1__0_,
  fifo_data_0__37_,fifo_data_0__36_,fifo_data_0__35_,fifo_data_0__34_,
  fifo_data_0__33_,fifo_data_0__32_,fifo_data_0__31_,fifo_data_0__30_,fifo_data_0__29_,
  fifo_data_0__28_,fifo_data_0__27_,fifo_data_0__26_,fifo_data_0__25_,fifo_data_0__24_,
  fifo_data_0__23_,fifo_data_0__22_,fifo_data_0__21_,fifo_data_0__20_,fifo_data_0__19_,
  fifo_data_0__18_,fifo_data_0__17_,fifo_data_0__16_,fifo_data_0__15_,
  fifo_data_0__14_,fifo_data_0__13_,fifo_data_0__12_,fifo_data_0__11_,fifo_data_0__10_,
  fifo_data_0__9_,fifo_data_0__8_,fifo_data_0__7_,fifo_data_0__6_,fifo_data_0__5_,
  fifo_data_0__4_,fifo_data_0__3_,fifo_data_0__2_,fifo_data_0__1_,fifo_data_0__0_;
  wire [1:0] fifo_valid;
  wire [4:0] fifo_yumi;
  assign link_o[118] = 1'b0;
  assign link_o[158] = 1'b0;
  assign link_o[198] = 1'b0;

  bsg_two_fifo_width_p38
  rof_0__fi_twofer
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(link_o[38]),
    .data_i(link_i[37:0]),
    .v_i(link_i[39]),
    .v_o(fifo_valid[0]),
    .data_o({ fifo_data_0__37_, fifo_data_0__36_, fifo_data_0__35_, fifo_data_0__34_, fifo_data_0__33_, fifo_data_0__32_, fifo_data_0__31_, fifo_data_0__30_, fifo_data_0__29_, fifo_data_0__28_, fifo_data_0__27_, fifo_data_0__26_, fifo_data_0__25_, fifo_data_0__24_, fifo_data_0__23_, fifo_data_0__22_, fifo_data_0__21_, fifo_data_0__20_, fifo_data_0__19_, fifo_data_0__18_, fifo_data_0__17_, fifo_data_0__16_, fifo_data_0__15_, fifo_data_0__14_, fifo_data_0__13_, fifo_data_0__12_, fifo_data_0__11_, fifo_data_0__10_, fifo_data_0__9_, fifo_data_0__8_, fifo_data_0__7_, fifo_data_0__6_, fifo_data_0__5_, fifo_data_0__4_, fifo_data_0__3_, fifo_data_0__2_, fifo_data_0__1_, fifo_data_0__0_ }),
    .yumi_i(fifo_yumi[0])
  );


  bsg_two_fifo_width_p38
  rof_1__fi_twofer
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(link_o[78]),
    .data_i(link_i[77:40]),
    .v_i(link_i[79]),
    .v_o(fifo_valid[1]),
    .data_o({ fifo_data_1__37_, fifo_data_1__36_, fifo_data_1__35_, fifo_data_1__34_, fifo_data_1__33_, fifo_data_1__32_, fifo_data_1__31_, fifo_data_1__30_, fifo_data_1__29_, fifo_data_1__28_, fifo_data_1__27_, fifo_data_1__26_, fifo_data_1__25_, fifo_data_1__24_, fifo_data_1__23_, fifo_data_1__22_, fifo_data_1__21_, fifo_data_1__20_, fifo_data_1__19_, fifo_data_1__18_, fifo_data_1__17_, fifo_data_1__16_, fifo_data_1__15_, fifo_data_1__14_, fifo_data_1__13_, fifo_data_1__12_, fifo_data_1__11_, fifo_data_1__10_, fifo_data_1__9_, fifo_data_1__8_, fifo_data_1__7_, fifo_data_1__6_, fifo_data_1__5_, fifo_data_1__4_, fifo_data_1__3_, fifo_data_1__2_, fifo_data_1__1_, fifo_data_1__0_ }),
    .yumi_i(fifo_yumi[1])
  );


  bsg_mesh_router_38_1_1_0_1c_0
  bmr
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_1__37_, fifo_data_1__36_, fifo_data_1__35_, fifo_data_1__34_, fifo_data_1__33_, fifo_data_1__32_, fifo_data_1__31_, fifo_data_1__30_, fifo_data_1__29_, fifo_data_1__28_, fifo_data_1__27_, fifo_data_1__26_, fifo_data_1__25_, fifo_data_1__24_, fifo_data_1__23_, fifo_data_1__22_, fifo_data_1__21_, fifo_data_1__20_, fifo_data_1__19_, fifo_data_1__18_, fifo_data_1__17_, fifo_data_1__16_, fifo_data_1__15_, fifo_data_1__14_, fifo_data_1__13_, fifo_data_1__12_, fifo_data_1__11_, fifo_data_1__10_, fifo_data_1__9_, fifo_data_1__8_, fifo_data_1__7_, fifo_data_1__6_, fifo_data_1__5_, fifo_data_1__4_, fifo_data_1__3_, fifo_data_1__2_, fifo_data_1__1_, fifo_data_1__0_, fifo_data_0__37_, fifo_data_0__36_, fifo_data_0__35_, fifo_data_0__34_, fifo_data_0__33_, fifo_data_0__32_, fifo_data_0__31_, fifo_data_0__30_, fifo_data_0__29_, fifo_data_0__28_, fifo_data_0__27_, fifo_data_0__26_, fifo_data_0__25_, fifo_data_0__24_, fifo_data_0__23_, fifo_data_0__22_, fifo_data_0__21_, fifo_data_0__20_, fifo_data_0__19_, fifo_data_0__18_, fifo_data_0__17_, fifo_data_0__16_, fifo_data_0__15_, fifo_data_0__14_, fifo_data_0__13_, fifo_data_0__12_, fifo_data_0__11_, fifo_data_0__10_, fifo_data_0__9_, fifo_data_0__8_, fifo_data_0__7_, fifo_data_0__6_, fifo_data_0__5_, fifo_data_0__4_, fifo_data_0__3_, fifo_data_0__2_, fifo_data_0__1_, fifo_data_0__0_ }),
    .v_i({ 1'b0, 1'b0, 1'b0, fifo_valid }),
    .yumi_o(fifo_yumi),
    .ready_i({ link_i[198:198], link_i[158:158], link_i[118:118], link_i[78:78], link_i[38:38] }),
    .data_o({ link_o[197:160], link_o[157:120], link_o[117:80], link_o[77:40], link_o[37:0] }),
    .v_o({ link_o[199:199], link_o[159:159], link_o[119:119], link_o[79:79], link_o[39:39] }),
    .my_x_i(my_x_i[0]),
    .my_y_i(my_y_i[0])
  );


endmodule



module bp_me_network_channel_mesh_packet_width_p36_num_src_p1_num_dst_p2_debug_p0
(
  clk_i,
  reset_i,
  src_data_i,
  src_v_i,
  src_ready_o,
  dst_data_o,
  dst_v_o,
  dst_ready_i
);

  input [35:0] src_data_i;
  input [0:0] src_v_i;
  output [0:0] src_ready_o;
  output [71:0] dst_data_o;
  output [1:0] dst_v_o;
  input [1:0] dst_ready_i;
  input clk_i;
  input reset_i;
  wire [0:0] src_ready_o;
  wire [71:0] dst_data_o;
  wire [1:0] dst_v_o;
  wire link_i_stitch_0__2__v_,link_i_stitch_0__2__ready_then_rev_,
  link_i_stitch_0__2__data__37_,link_i_stitch_0__2__data__36_,link_i_stitch_0__2__data__35_,
  link_i_stitch_0__2__data__34_,link_i_stitch_0__2__data__33_,link_i_stitch_0__2__data__32_,
  link_i_stitch_0__2__data__31_,link_i_stitch_0__2__data__30_,
  link_i_stitch_0__2__data__29_,link_i_stitch_0__2__data__28_,link_i_stitch_0__2__data__27_,
  link_i_stitch_0__2__data__26_,link_i_stitch_0__2__data__25_,link_i_stitch_0__2__data__24_,
  link_i_stitch_0__2__data__23_,link_i_stitch_0__2__data__22_,
  link_i_stitch_0__2__data__21_,link_i_stitch_0__2__data__20_,link_i_stitch_0__2__data__19_,
  link_i_stitch_0__2__data__18_,link_i_stitch_0__2__data__17_,link_i_stitch_0__2__data__16_,
  link_i_stitch_0__2__data__15_,link_i_stitch_0__2__data__14_,
  link_i_stitch_0__2__data__13_,link_i_stitch_0__2__data__12_,link_i_stitch_0__2__data__11_,
  link_i_stitch_0__2__data__10_,link_i_stitch_0__2__data__9_,link_i_stitch_0__2__data__8_,
  link_i_stitch_0__2__data__7_,link_i_stitch_0__2__data__6_,
  link_i_stitch_0__2__data__5_,link_i_stitch_0__2__data__4_,link_i_stitch_0__2__data__3_,
  link_i_stitch_0__2__data__2_,link_i_stitch_0__2__data__1_,link_i_stitch_0__2__data__0_,
  link_o_stitch_1__4__v_,link_o_stitch_1__4__ready_then_rev_,link_o_stitch_1__4__data__37_,
  link_o_stitch_1__4__data__36_,link_o_stitch_1__4__data__35_,
  link_o_stitch_1__4__data__34_,link_o_stitch_1__4__data__33_,link_o_stitch_1__4__data__32_,
  link_o_stitch_1__4__data__31_,link_o_stitch_1__4__data__30_,link_o_stitch_1__4__data__29_,
  link_o_stitch_1__4__data__28_,link_o_stitch_1__4__data__27_,
  link_o_stitch_1__4__data__26_,link_o_stitch_1__4__data__25_,link_o_stitch_1__4__data__24_,
  link_o_stitch_1__4__data__23_,link_o_stitch_1__4__data__22_,link_o_stitch_1__4__data__21_,
  link_o_stitch_1__4__data__20_,link_o_stitch_1__4__data__19_,
  link_o_stitch_1__4__data__18_,link_o_stitch_1__4__data__17_,link_o_stitch_1__4__data__16_,
  link_o_stitch_1__4__data__15_,link_o_stitch_1__4__data__14_,link_o_stitch_1__4__data__13_,
  link_o_stitch_1__4__data__12_,link_o_stitch_1__4__data__11_,
  link_o_stitch_1__4__data__10_,link_o_stitch_1__4__data__9_,link_o_stitch_1__4__data__8_,
  link_o_stitch_1__4__data__7_,link_o_stitch_1__4__data__6_,link_o_stitch_1__4__data__5_,
  link_o_stitch_1__4__data__4_,link_o_stitch_1__4__data__3_,link_o_stitch_1__4__data__2_,
  link_o_stitch_1__4__data__1_,link_o_stitch_1__4__data__0_,
  link_o_stitch_1__3__v_,link_o_stitch_1__3__ready_then_rev_,link_o_stitch_1__3__data__37_,
  link_o_stitch_1__3__data__36_,link_o_stitch_1__3__data__35_,link_o_stitch_1__3__data__34_,
  link_o_stitch_1__3__data__33_,link_o_stitch_1__3__data__32_,
  link_o_stitch_1__3__data__31_,link_o_stitch_1__3__data__30_,link_o_stitch_1__3__data__29_,
  link_o_stitch_1__3__data__28_,link_o_stitch_1__3__data__27_,link_o_stitch_1__3__data__26_,
  link_o_stitch_1__3__data__25_,link_o_stitch_1__3__data__24_,
  link_o_stitch_1__3__data__23_,link_o_stitch_1__3__data__22_,link_o_stitch_1__3__data__21_,
  link_o_stitch_1__3__data__20_,link_o_stitch_1__3__data__19_,link_o_stitch_1__3__data__18_,
  link_o_stitch_1__3__data__17_,link_o_stitch_1__3__data__16_,
  link_o_stitch_1__3__data__15_,link_o_stitch_1__3__data__14_,link_o_stitch_1__3__data__13_,
  link_o_stitch_1__3__data__12_,link_o_stitch_1__3__data__11_,link_o_stitch_1__3__data__10_,
  link_o_stitch_1__3__data__9_,link_o_stitch_1__3__data__8_,
  link_o_stitch_1__3__data__7_,link_o_stitch_1__3__data__6_,link_o_stitch_1__3__data__5_,
  link_o_stitch_1__3__data__4_,link_o_stitch_1__3__data__3_,link_o_stitch_1__3__data__2_,
  link_o_stitch_1__3__data__1_,link_o_stitch_1__3__data__0_,link_o_stitch_1__2__v_,
  link_o_stitch_1__2__ready_then_rev_,link_o_stitch_1__2__data__37_,
  link_o_stitch_1__2__data__36_,link_o_stitch_1__2__data__35_,link_o_stitch_1__2__data__34_,
  link_o_stitch_1__2__data__33_,link_o_stitch_1__2__data__32_,link_o_stitch_1__2__data__31_,
  link_o_stitch_1__2__data__30_,link_o_stitch_1__2__data__29_,
  link_o_stitch_1__2__data__28_,link_o_stitch_1__2__data__27_,link_o_stitch_1__2__data__26_,
  link_o_stitch_1__2__data__25_,link_o_stitch_1__2__data__24_,link_o_stitch_1__2__data__23_,
  link_o_stitch_1__2__data__22_,link_o_stitch_1__2__data__21_,
  link_o_stitch_1__2__data__20_,link_o_stitch_1__2__data__19_,link_o_stitch_1__2__data__18_,
  link_o_stitch_1__2__data__17_,link_o_stitch_1__2__data__16_,link_o_stitch_1__2__data__15_,
  link_o_stitch_1__2__data__14_,link_o_stitch_1__2__data__13_,
  link_o_stitch_1__2__data__12_,link_o_stitch_1__2__data__11_,link_o_stitch_1__2__data__10_,
  link_o_stitch_1__2__data__9_,link_o_stitch_1__2__data__8_,link_o_stitch_1__2__data__7_,
  link_o_stitch_1__2__data__6_,link_o_stitch_1__2__data__5_,link_o_stitch_1__2__data__4_,
  link_o_stitch_1__2__data__3_,link_o_stitch_1__2__data__2_,
  link_o_stitch_1__2__data__1_,link_o_stitch_1__2__data__0_,link_o_stitch_1__0__ready_then_rev_,
  link_o_stitch_1__0__data__1_,link_o_stitch_1__0__data__0_,link_o_stitch_0__4__v_,
  link_o_stitch_0__4__data__37_,link_o_stitch_0__4__data__36_,
  link_o_stitch_0__4__data__35_,link_o_stitch_0__4__data__34_,link_o_stitch_0__4__data__33_,
  link_o_stitch_0__4__data__32_,link_o_stitch_0__4__data__31_,link_o_stitch_0__4__data__30_,
  link_o_stitch_0__4__data__29_,link_o_stitch_0__4__data__28_,
  link_o_stitch_0__4__data__27_,link_o_stitch_0__4__data__26_,link_o_stitch_0__4__data__25_,
  link_o_stitch_0__4__data__24_,link_o_stitch_0__4__data__23_,link_o_stitch_0__4__data__22_,
  link_o_stitch_0__4__data__21_,link_o_stitch_0__4__data__20_,
  link_o_stitch_0__4__data__19_,link_o_stitch_0__4__data__18_,link_o_stitch_0__4__data__17_,
  link_o_stitch_0__4__data__16_,link_o_stitch_0__4__data__15_,link_o_stitch_0__4__data__14_,
  link_o_stitch_0__4__data__13_,link_o_stitch_0__4__data__12_,
  link_o_stitch_0__4__data__11_,link_o_stitch_0__4__data__10_,link_o_stitch_0__4__data__9_,
  link_o_stitch_0__4__data__8_,link_o_stitch_0__4__data__7_,link_o_stitch_0__4__data__6_,
  link_o_stitch_0__4__data__5_,link_o_stitch_0__4__data__4_,link_o_stitch_0__4__data__3_,
  link_o_stitch_0__4__data__2_,link_o_stitch_0__4__data__1_,
  link_o_stitch_0__4__data__0_,link_o_stitch_0__3__v_,link_o_stitch_0__3__ready_then_rev_,
  link_o_stitch_0__3__data__37_,link_o_stitch_0__3__data__36_,link_o_stitch_0__3__data__35_,
  link_o_stitch_0__3__data__34_,link_o_stitch_0__3__data__33_,
  link_o_stitch_0__3__data__32_,link_o_stitch_0__3__data__31_,link_o_stitch_0__3__data__30_,
  link_o_stitch_0__3__data__29_,link_o_stitch_0__3__data__28_,link_o_stitch_0__3__data__27_,
  link_o_stitch_0__3__data__26_,link_o_stitch_0__3__data__25_,
  link_o_stitch_0__3__data__24_,link_o_stitch_0__3__data__23_,link_o_stitch_0__3__data__22_,
  link_o_stitch_0__3__data__21_,link_o_stitch_0__3__data__20_,link_o_stitch_0__3__data__19_,
  link_o_stitch_0__3__data__18_,link_o_stitch_0__3__data__17_,
  link_o_stitch_0__3__data__16_,link_o_stitch_0__3__data__15_,link_o_stitch_0__3__data__14_,
  link_o_stitch_0__3__data__13_,link_o_stitch_0__3__data__12_,link_o_stitch_0__3__data__11_,
  link_o_stitch_0__3__data__10_,link_o_stitch_0__3__data__9_,link_o_stitch_0__3__data__8_,
  link_o_stitch_0__3__data__7_,link_o_stitch_0__3__data__6_,
  link_o_stitch_0__3__data__5_,link_o_stitch_0__3__data__4_,link_o_stitch_0__3__data__3_,
  link_o_stitch_0__3__data__2_,link_o_stitch_0__3__data__1_,link_o_stitch_0__3__data__0_,
  link_o_stitch_0__2__v_,link_o_stitch_0__2__ready_then_rev_,
  link_o_stitch_0__2__data__37_,link_o_stitch_0__2__data__36_,link_o_stitch_0__2__data__35_,
  link_o_stitch_0__2__data__34_,link_o_stitch_0__2__data__33_,link_o_stitch_0__2__data__32_,
  link_o_stitch_0__2__data__31_,link_o_stitch_0__2__data__30_,
  link_o_stitch_0__2__data__29_,link_o_stitch_0__2__data__28_,link_o_stitch_0__2__data__27_,
  link_o_stitch_0__2__data__26_,link_o_stitch_0__2__data__25_,link_o_stitch_0__2__data__24_,
  link_o_stitch_0__2__data__23_,link_o_stitch_0__2__data__22_,
  link_o_stitch_0__2__data__21_,link_o_stitch_0__2__data__20_,link_o_stitch_0__2__data__19_,
  link_o_stitch_0__2__data__18_,link_o_stitch_0__2__data__17_,link_o_stitch_0__2__data__16_,
  link_o_stitch_0__2__data__15_,link_o_stitch_0__2__data__14_,
  link_o_stitch_0__2__data__13_,link_o_stitch_0__2__data__12_,link_o_stitch_0__2__data__11_,
  link_o_stitch_0__2__data__10_,link_o_stitch_0__2__data__9_,link_o_stitch_0__2__data__8_,
  link_o_stitch_0__2__data__7_,link_o_stitch_0__2__data__6_,link_o_stitch_0__2__data__5_,
  link_o_stitch_0__2__data__4_,link_o_stitch_0__2__data__3_,
  link_o_stitch_0__2__data__2_,link_o_stitch_0__2__data__1_,link_o_stitch_0__2__data__0_,
  link_o_stitch_0__1__v_,link_o_stitch_0__1__ready_then_rev_,link_o_stitch_0__1__data__37_,
  link_o_stitch_0__1__data__36_,link_o_stitch_0__1__data__35_,link_o_stitch_0__1__data__34_,
  link_o_stitch_0__1__data__33_,link_o_stitch_0__1__data__32_,
  link_o_stitch_0__1__data__31_,link_o_stitch_0__1__data__30_,link_o_stitch_0__1__data__29_,
  link_o_stitch_0__1__data__28_,link_o_stitch_0__1__data__27_,link_o_stitch_0__1__data__26_,
  link_o_stitch_0__1__data__25_,link_o_stitch_0__1__data__24_,
  link_o_stitch_0__1__data__23_,link_o_stitch_0__1__data__22_,link_o_stitch_0__1__data__21_,
  link_o_stitch_0__1__data__20_,link_o_stitch_0__1__data__19_,link_o_stitch_0__1__data__18_,
  link_o_stitch_0__1__data__17_,link_o_stitch_0__1__data__16_,
  link_o_stitch_0__1__data__15_,link_o_stitch_0__1__data__14_,link_o_stitch_0__1__data__13_,
  link_o_stitch_0__1__data__12_,link_o_stitch_0__1__data__11_,link_o_stitch_0__1__data__10_,
  link_o_stitch_0__1__data__9_,link_o_stitch_0__1__data__8_,
  link_o_stitch_0__1__data__7_,link_o_stitch_0__1__data__6_,link_o_stitch_0__1__data__5_,
  link_o_stitch_0__1__data__4_,link_o_stitch_0__1__data__3_,link_o_stitch_0__1__data__2_,
  link_o_stitch_0__1__data__1_,link_o_stitch_0__1__data__0_,
  link_o_stitch_0__0__ready_then_rev_,link_o_stitch_0__0__data__1_,link_o_stitch_0__0__data__0_;

  bsg_mesh_router_buffered_38_1_1_0_5_0a_0_40_00
  rof_0__fi2_efi3_coherence_network_channel_node
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .link_i({ src_v_i[0:0], 1'b0, src_data_i, 1'b1, src_data_i[35:35], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, link_i_stitch_0__2__v_, link_i_stitch_0__2__ready_then_rev_, link_i_stitch_0__2__data__37_, link_i_stitch_0__2__data__36_, link_i_stitch_0__2__data__35_, link_i_stitch_0__2__data__34_, link_i_stitch_0__2__data__33_, link_i_stitch_0__2__data__32_, link_i_stitch_0__2__data__31_, link_i_stitch_0__2__data__30_, link_i_stitch_0__2__data__29_, link_i_stitch_0__2__data__28_, link_i_stitch_0__2__data__27_, link_i_stitch_0__2__data__26_, link_i_stitch_0__2__data__25_, link_i_stitch_0__2__data__24_, link_i_stitch_0__2__data__23_, link_i_stitch_0__2__data__22_, link_i_stitch_0__2__data__21_, link_i_stitch_0__2__data__20_, link_i_stitch_0__2__data__19_, link_i_stitch_0__2__data__18_, link_i_stitch_0__2__data__17_, link_i_stitch_0__2__data__16_, link_i_stitch_0__2__data__15_, link_i_stitch_0__2__data__14_, link_i_stitch_0__2__data__13_, link_i_stitch_0__2__data__12_, link_i_stitch_0__2__data__11_, link_i_stitch_0__2__data__10_, link_i_stitch_0__2__data__9_, link_i_stitch_0__2__data__8_, link_i_stitch_0__2__data__7_, link_i_stitch_0__2__data__6_, link_i_stitch_0__2__data__5_, link_i_stitch_0__2__data__4_, link_i_stitch_0__2__data__3_, link_i_stitch_0__2__data__2_, link_i_stitch_0__2__data__1_, link_i_stitch_0__2__data__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, dst_ready_i[0:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .link_o({ link_o_stitch_0__4__v_, src_ready_o[0:0], link_o_stitch_0__4__data__37_, link_o_stitch_0__4__data__36_, link_o_stitch_0__4__data__35_, link_o_stitch_0__4__data__34_, link_o_stitch_0__4__data__33_, link_o_stitch_0__4__data__32_, link_o_stitch_0__4__data__31_, link_o_stitch_0__4__data__30_, link_o_stitch_0__4__data__29_, link_o_stitch_0__4__data__28_, link_o_stitch_0__4__data__27_, link_o_stitch_0__4__data__26_, link_o_stitch_0__4__data__25_, link_o_stitch_0__4__data__24_, link_o_stitch_0__4__data__23_, link_o_stitch_0__4__data__22_, link_o_stitch_0__4__data__21_, link_o_stitch_0__4__data__20_, link_o_stitch_0__4__data__19_, link_o_stitch_0__4__data__18_, link_o_stitch_0__4__data__17_, link_o_stitch_0__4__data__16_, link_o_stitch_0__4__data__15_, link_o_stitch_0__4__data__14_, link_o_stitch_0__4__data__13_, link_o_stitch_0__4__data__12_, link_o_stitch_0__4__data__11_, link_o_stitch_0__4__data__10_, link_o_stitch_0__4__data__9_, link_o_stitch_0__4__data__8_, link_o_stitch_0__4__data__7_, link_o_stitch_0__4__data__6_, link_o_stitch_0__4__data__5_, link_o_stitch_0__4__data__4_, link_o_stitch_0__4__data__3_, link_o_stitch_0__4__data__2_, link_o_stitch_0__4__data__1_, link_o_stitch_0__4__data__0_, link_o_stitch_0__3__v_, link_o_stitch_0__3__ready_then_rev_, link_o_stitch_0__3__data__37_, link_o_stitch_0__3__data__36_, link_o_stitch_0__3__data__35_, link_o_stitch_0__3__data__34_, link_o_stitch_0__3__data__33_, link_o_stitch_0__3__data__32_, link_o_stitch_0__3__data__31_, link_o_stitch_0__3__data__30_, link_o_stitch_0__3__data__29_, link_o_stitch_0__3__data__28_, link_o_stitch_0__3__data__27_, link_o_stitch_0__3__data__26_, link_o_stitch_0__3__data__25_, link_o_stitch_0__3__data__24_, link_o_stitch_0__3__data__23_, link_o_stitch_0__3__data__22_, link_o_stitch_0__3__data__21_, link_o_stitch_0__3__data__20_, link_o_stitch_0__3__data__19_, link_o_stitch_0__3__data__18_, link_o_stitch_0__3__data__17_, link_o_stitch_0__3__data__16_, link_o_stitch_0__3__data__15_, link_o_stitch_0__3__data__14_, link_o_stitch_0__3__data__13_, link_o_stitch_0__3__data__12_, link_o_stitch_0__3__data__11_, link_o_stitch_0__3__data__10_, link_o_stitch_0__3__data__9_, link_o_stitch_0__3__data__8_, link_o_stitch_0__3__data__7_, link_o_stitch_0__3__data__6_, link_o_stitch_0__3__data__5_, link_o_stitch_0__3__data__4_, link_o_stitch_0__3__data__3_, link_o_stitch_0__3__data__2_, link_o_stitch_0__3__data__1_, link_o_stitch_0__3__data__0_, link_o_stitch_0__2__v_, link_o_stitch_0__2__ready_then_rev_, link_o_stitch_0__2__data__37_, link_o_stitch_0__2__data__36_, link_o_stitch_0__2__data__35_, link_o_stitch_0__2__data__34_, link_o_stitch_0__2__data__33_, link_o_stitch_0__2__data__32_, link_o_stitch_0__2__data__31_, link_o_stitch_0__2__data__30_, link_o_stitch_0__2__data__29_, link_o_stitch_0__2__data__28_, link_o_stitch_0__2__data__27_, link_o_stitch_0__2__data__26_, link_o_stitch_0__2__data__25_, link_o_stitch_0__2__data__24_, link_o_stitch_0__2__data__23_, link_o_stitch_0__2__data__22_, link_o_stitch_0__2__data__21_, link_o_stitch_0__2__data__20_, link_o_stitch_0__2__data__19_, link_o_stitch_0__2__data__18_, link_o_stitch_0__2__data__17_, link_o_stitch_0__2__data__16_, link_o_stitch_0__2__data__15_, link_o_stitch_0__2__data__14_, link_o_stitch_0__2__data__13_, link_o_stitch_0__2__data__12_, link_o_stitch_0__2__data__11_, link_o_stitch_0__2__data__10_, link_o_stitch_0__2__data__9_, link_o_stitch_0__2__data__8_, link_o_stitch_0__2__data__7_, link_o_stitch_0__2__data__6_, link_o_stitch_0__2__data__5_, link_o_stitch_0__2__data__4_, link_o_stitch_0__2__data__3_, link_o_stitch_0__2__data__2_, link_o_stitch_0__2__data__1_, link_o_stitch_0__2__data__0_, link_o_stitch_0__1__v_, link_o_stitch_0__1__ready_then_rev_, link_o_stitch_0__1__data__37_, link_o_stitch_0__1__data__36_, link_o_stitch_0__1__data__35_, link_o_stitch_0__1__data__34_, link_o_stitch_0__1__data__33_, link_o_stitch_0__1__data__32_, link_o_stitch_0__1__data__31_, link_o_stitch_0__1__data__30_, link_o_stitch_0__1__data__29_, link_o_stitch_0__1__data__28_, link_o_stitch_0__1__data__27_, link_o_stitch_0__1__data__26_, link_o_stitch_0__1__data__25_, link_o_stitch_0__1__data__24_, link_o_stitch_0__1__data__23_, link_o_stitch_0__1__data__22_, link_o_stitch_0__1__data__21_, link_o_stitch_0__1__data__20_, link_o_stitch_0__1__data__19_, link_o_stitch_0__1__data__18_, link_o_stitch_0__1__data__17_, link_o_stitch_0__1__data__16_, link_o_stitch_0__1__data__15_, link_o_stitch_0__1__data__14_, link_o_stitch_0__1__data__13_, link_o_stitch_0__1__data__12_, link_o_stitch_0__1__data__11_, link_o_stitch_0__1__data__10_, link_o_stitch_0__1__data__9_, link_o_stitch_0__1__data__8_, link_o_stitch_0__1__data__7_, link_o_stitch_0__1__data__6_, link_o_stitch_0__1__data__5_, link_o_stitch_0__1__data__4_, link_o_stitch_0__1__data__3_, link_o_stitch_0__1__data__2_, link_o_stitch_0__1__data__1_, link_o_stitch_0__1__data__0_, dst_v_o[0:0], link_o_stitch_0__0__ready_then_rev_, dst_data_o[35:0], link_o_stitch_0__0__data__1_, link_o_stitch_0__0__data__0_ }),
    .my_x_i(1'b0),
    .my_y_i(1'b1)
  );


  bsg_mesh_router_buffered_38_1_1_0_5_1c_0_40_00
  rof_1__efi2_fi9_coherence_network_channel_node
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .link_i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, link_o_stitch_0__2__v_, link_o_stitch_0__2__ready_then_rev_, link_o_stitch_0__2__data__37_, link_o_stitch_0__2__data__36_, link_o_stitch_0__2__data__35_, link_o_stitch_0__2__data__34_, link_o_stitch_0__2__data__33_, link_o_stitch_0__2__data__32_, link_o_stitch_0__2__data__31_, link_o_stitch_0__2__data__30_, link_o_stitch_0__2__data__29_, link_o_stitch_0__2__data__28_, link_o_stitch_0__2__data__27_, link_o_stitch_0__2__data__26_, link_o_stitch_0__2__data__25_, link_o_stitch_0__2__data__24_, link_o_stitch_0__2__data__23_, link_o_stitch_0__2__data__22_, link_o_stitch_0__2__data__21_, link_o_stitch_0__2__data__20_, link_o_stitch_0__2__data__19_, link_o_stitch_0__2__data__18_, link_o_stitch_0__2__data__17_, link_o_stitch_0__2__data__16_, link_o_stitch_0__2__data__15_, link_o_stitch_0__2__data__14_, link_o_stitch_0__2__data__13_, link_o_stitch_0__2__data__12_, link_o_stitch_0__2__data__11_, link_o_stitch_0__2__data__10_, link_o_stitch_0__2__data__9_, link_o_stitch_0__2__data__8_, link_o_stitch_0__2__data__7_, link_o_stitch_0__2__data__6_, link_o_stitch_0__2__data__5_, link_o_stitch_0__2__data__4_, link_o_stitch_0__2__data__3_, link_o_stitch_0__2__data__2_, link_o_stitch_0__2__data__1_, link_o_stitch_0__2__data__0_, 1'b0, dst_ready_i[1:1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .link_o({ link_o_stitch_1__4__v_, link_o_stitch_1__4__ready_then_rev_, link_o_stitch_1__4__data__37_, link_o_stitch_1__4__data__36_, link_o_stitch_1__4__data__35_, link_o_stitch_1__4__data__34_, link_o_stitch_1__4__data__33_, link_o_stitch_1__4__data__32_, link_o_stitch_1__4__data__31_, link_o_stitch_1__4__data__30_, link_o_stitch_1__4__data__29_, link_o_stitch_1__4__data__28_, link_o_stitch_1__4__data__27_, link_o_stitch_1__4__data__26_, link_o_stitch_1__4__data__25_, link_o_stitch_1__4__data__24_, link_o_stitch_1__4__data__23_, link_o_stitch_1__4__data__22_, link_o_stitch_1__4__data__21_, link_o_stitch_1__4__data__20_, link_o_stitch_1__4__data__19_, link_o_stitch_1__4__data__18_, link_o_stitch_1__4__data__17_, link_o_stitch_1__4__data__16_, link_o_stitch_1__4__data__15_, link_o_stitch_1__4__data__14_, link_o_stitch_1__4__data__13_, link_o_stitch_1__4__data__12_, link_o_stitch_1__4__data__11_, link_o_stitch_1__4__data__10_, link_o_stitch_1__4__data__9_, link_o_stitch_1__4__data__8_, link_o_stitch_1__4__data__7_, link_o_stitch_1__4__data__6_, link_o_stitch_1__4__data__5_, link_o_stitch_1__4__data__4_, link_o_stitch_1__4__data__3_, link_o_stitch_1__4__data__2_, link_o_stitch_1__4__data__1_, link_o_stitch_1__4__data__0_, link_o_stitch_1__3__v_, link_o_stitch_1__3__ready_then_rev_, link_o_stitch_1__3__data__37_, link_o_stitch_1__3__data__36_, link_o_stitch_1__3__data__35_, link_o_stitch_1__3__data__34_, link_o_stitch_1__3__data__33_, link_o_stitch_1__3__data__32_, link_o_stitch_1__3__data__31_, link_o_stitch_1__3__data__30_, link_o_stitch_1__3__data__29_, link_o_stitch_1__3__data__28_, link_o_stitch_1__3__data__27_, link_o_stitch_1__3__data__26_, link_o_stitch_1__3__data__25_, link_o_stitch_1__3__data__24_, link_o_stitch_1__3__data__23_, link_o_stitch_1__3__data__22_, link_o_stitch_1__3__data__21_, link_o_stitch_1__3__data__20_, link_o_stitch_1__3__data__19_, link_o_stitch_1__3__data__18_, link_o_stitch_1__3__data__17_, link_o_stitch_1__3__data__16_, link_o_stitch_1__3__data__15_, link_o_stitch_1__3__data__14_, link_o_stitch_1__3__data__13_, link_o_stitch_1__3__data__12_, link_o_stitch_1__3__data__11_, link_o_stitch_1__3__data__10_, link_o_stitch_1__3__data__9_, link_o_stitch_1__3__data__8_, link_o_stitch_1__3__data__7_, link_o_stitch_1__3__data__6_, link_o_stitch_1__3__data__5_, link_o_stitch_1__3__data__4_, link_o_stitch_1__3__data__3_, link_o_stitch_1__3__data__2_, link_o_stitch_1__3__data__1_, link_o_stitch_1__3__data__0_, link_o_stitch_1__2__v_, link_o_stitch_1__2__ready_then_rev_, link_o_stitch_1__2__data__37_, link_o_stitch_1__2__data__36_, link_o_stitch_1__2__data__35_, link_o_stitch_1__2__data__34_, link_o_stitch_1__2__data__33_, link_o_stitch_1__2__data__32_, link_o_stitch_1__2__data__31_, link_o_stitch_1__2__data__30_, link_o_stitch_1__2__data__29_, link_o_stitch_1__2__data__28_, link_o_stitch_1__2__data__27_, link_o_stitch_1__2__data__26_, link_o_stitch_1__2__data__25_, link_o_stitch_1__2__data__24_, link_o_stitch_1__2__data__23_, link_o_stitch_1__2__data__22_, link_o_stitch_1__2__data__21_, link_o_stitch_1__2__data__20_, link_o_stitch_1__2__data__19_, link_o_stitch_1__2__data__18_, link_o_stitch_1__2__data__17_, link_o_stitch_1__2__data__16_, link_o_stitch_1__2__data__15_, link_o_stitch_1__2__data__14_, link_o_stitch_1__2__data__13_, link_o_stitch_1__2__data__12_, link_o_stitch_1__2__data__11_, link_o_stitch_1__2__data__10_, link_o_stitch_1__2__data__9_, link_o_stitch_1__2__data__8_, link_o_stitch_1__2__data__7_, link_o_stitch_1__2__data__6_, link_o_stitch_1__2__data__5_, link_o_stitch_1__2__data__4_, link_o_stitch_1__2__data__3_, link_o_stitch_1__2__data__2_, link_o_stitch_1__2__data__1_, link_o_stitch_1__2__data__0_, link_i_stitch_0__2__v_, link_i_stitch_0__2__ready_then_rev_, link_i_stitch_0__2__data__37_, link_i_stitch_0__2__data__36_, link_i_stitch_0__2__data__35_, link_i_stitch_0__2__data__34_, link_i_stitch_0__2__data__33_, link_i_stitch_0__2__data__32_, link_i_stitch_0__2__data__31_, link_i_stitch_0__2__data__30_, link_i_stitch_0__2__data__29_, link_i_stitch_0__2__data__28_, link_i_stitch_0__2__data__27_, link_i_stitch_0__2__data__26_, link_i_stitch_0__2__data__25_, link_i_stitch_0__2__data__24_, link_i_stitch_0__2__data__23_, link_i_stitch_0__2__data__22_, link_i_stitch_0__2__data__21_, link_i_stitch_0__2__data__20_, link_i_stitch_0__2__data__19_, link_i_stitch_0__2__data__18_, link_i_stitch_0__2__data__17_, link_i_stitch_0__2__data__16_, link_i_stitch_0__2__data__15_, link_i_stitch_0__2__data__14_, link_i_stitch_0__2__data__13_, link_i_stitch_0__2__data__12_, link_i_stitch_0__2__data__11_, link_i_stitch_0__2__data__10_, link_i_stitch_0__2__data__9_, link_i_stitch_0__2__data__8_, link_i_stitch_0__2__data__7_, link_i_stitch_0__2__data__6_, link_i_stitch_0__2__data__5_, link_i_stitch_0__2__data__4_, link_i_stitch_0__2__data__3_, link_i_stitch_0__2__data__2_, link_i_stitch_0__2__data__1_, link_i_stitch_0__2__data__0_, dst_v_o[1:1], link_o_stitch_1__0__ready_then_rev_, dst_data_o[71:36], link_o_stitch_1__0__data__1_, link_o_stitch_1__0__data__0_ }),
    .my_x_i(1'b1),
    .my_y_i(1'b1)
  );


endmodule



module bsg_mem_p99
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [98:0] w_data_i;
  input [0:0] r_addr_i;
  output [98:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [98:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  reg [197:0] mem;
  assign r_data_o[98] = (N3)? mem[98] :
                        (N0)? mem[197] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[97] = (N3)? mem[97] :
                        (N0)? mem[196] : 1'b0;
  assign r_data_o[96] = (N3)? mem[96] :
                        (N0)? mem[195] : 1'b0;
  assign r_data_o[95] = (N3)? mem[95] :
                        (N0)? mem[194] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] :
                        (N0)? mem[193] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] :
                        (N0)? mem[192] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] :
                        (N0)? mem[191] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] :
                        (N0)? mem[190] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] :
                        (N0)? mem[189] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] :
                        (N0)? mem[188] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] :
                        (N0)? mem[187] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] :
                        (N0)? mem[186] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] :
                        (N0)? mem[185] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] :
                        (N0)? mem[184] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] :
                        (N0)? mem[183] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] :
                        (N0)? mem[182] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] :
                        (N0)? mem[181] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] :
                        (N0)? mem[180] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] :
                        (N0)? mem[179] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] :
                        (N0)? mem[178] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] :
                        (N0)? mem[177] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] :
                        (N0)? mem[176] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] :
                        (N0)? mem[175] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] :
                        (N0)? mem[174] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] :
                        (N0)? mem[173] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] :
                        (N0)? mem[172] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] :
                        (N0)? mem[171] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] :
                        (N0)? mem[170] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] :
                        (N0)? mem[169] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] :
                        (N0)? mem[168] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] :
                        (N0)? mem[167] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] :
                        (N0)? mem[166] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] :
                        (N0)? mem[165] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] :
                        (N0)? mem[164] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] :
                        (N0)? mem[163] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] :
                        (N0)? mem[162] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] :
                        (N0)? mem[161] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] :
                        (N0)? mem[160] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] :
                        (N0)? mem[159] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] :
                        (N0)? mem[158] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] :
                        (N0)? mem[157] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] :
                        (N0)? mem[156] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] :
                        (N0)? mem[155] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] :
                        (N0)? mem[154] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] :
                        (N0)? mem[153] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] :
                        (N0)? mem[152] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] :
                        (N0)? mem[151] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] :
                        (N0)? mem[150] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] :
                        (N0)? mem[149] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] :
                        (N0)? mem[148] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] :
                        (N0)? mem[147] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] :
                        (N0)? mem[146] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] :
                        (N0)? mem[145] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] :
                        (N0)? mem[144] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] :
                        (N0)? mem[143] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] :
                        (N0)? mem[142] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] :
                        (N0)? mem[141] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] :
                        (N0)? mem[140] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] :
                        (N0)? mem[139] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] :
                        (N0)? mem[138] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] :
                        (N0)? mem[137] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] :
                        (N0)? mem[136] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] :
                        (N0)? mem[135] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] :
                        (N0)? mem[134] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] :
                        (N0)? mem[133] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] :
                        (N0)? mem[132] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] :
                        (N0)? mem[131] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] :
                        (N0)? mem[130] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] :
                        (N0)? mem[129] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] :
                        (N0)? mem[128] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] :
                        (N0)? mem[127] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] :
                        (N0)? mem[126] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] :
                        (N0)? mem[125] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] :
                        (N0)? mem[124] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] :
                        (N0)? mem[123] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] :
                        (N0)? mem[122] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] :
                        (N0)? mem[121] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] :
                        (N0)? mem[120] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] :
                        (N0)? mem[119] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] :
                        (N0)? mem[118] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] :
                        (N0)? mem[117] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] :
                        (N0)? mem[116] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] :
                        (N0)? mem[115] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] :
                        (N0)? mem[114] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] :
                        (N0)? mem[113] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] :
                        (N0)? mem[112] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] :
                        (N0)? mem[111] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] :
                        (N0)? mem[110] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] :
                        (N0)? mem[109] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] :
                       (N0)? mem[108] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] :
                       (N0)? mem[107] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] :
                       (N0)? mem[106] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] :
                       (N0)? mem[105] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] :
                       (N0)? mem[104] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] :
                       (N0)? mem[103] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] :
                       (N0)? mem[102] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] :
                       (N0)? mem[101] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] :
                       (N0)? mem[100] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] :
                       (N0)? mem[99] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } :
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      { mem[197:99] } <= { w_data_i[98:0] };
    end
    if(N7) begin
      { mem[98:0] } <= { w_data_i[98:0] };
    end
  end


endmodule



module bsg_mem_1r1w_width_p99_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [98:0] w_data_i;
  input [0:0] r_addr_i;
  output [98:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [98:0] r_data_o;

  bsg_mem_p99
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p99
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [98:0] data_i;
  output [98:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [98:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p99_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 :
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 :
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 :
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 :
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 :
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 :
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end
    if(N9) begin
      tail_r <= N10;
    end
    if(N11) begin
      head_r <= N12;
    end
  end


endmodule



module bsg_mux_one_hot_width_p99_els_p4
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [395:0] data_i;
  input [3:0] sel_one_hot_i;
  output [98:0] data_o;
  wire [98:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197;
  wire [395:0] data_masked;
  assign data_masked[98] = data_i[98] & sel_one_hot_i[0];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[0];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[0];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[0];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[0];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[0];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[0];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[0];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[0];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[0];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[0];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[0];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[0];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[0];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[0];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[0];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[0];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[0];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[0];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[0];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[0];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[0];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[0];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[0];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[0];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[0];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[0];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[0];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[0];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[0];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[0];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[1];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[1];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[1];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[1];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[1];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[1];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[1];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[1];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[1];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[1];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[1];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[1];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[1];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[1];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[1];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[1];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[1];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[1];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[1];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[1];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[1];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[1];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[1];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[1];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[1];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[1];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[1];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[1];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[1];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[1];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[1];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[1];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[1];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[1];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[1];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[1];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[1];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[1];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[1];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[1];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[1];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[1];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[1];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[1];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[1];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[1];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[1];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[1];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[1];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[1];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[1];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[1];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[1];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[1];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[1];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[1];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[1];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[1];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[1];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[1];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[1];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[1];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[1];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[1];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[1];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[1];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[1];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[1];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[1];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[2];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[2];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[2];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[2];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[2];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[2];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[2];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[2];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[2];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[2];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[2];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[2];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[2];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[2];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[2];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[2];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[2];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[2];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[2];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[2];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[2];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[2];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[2];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[2];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[2];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[2];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[2];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[2];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[2];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[2];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[2];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[2];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[2];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[2];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[2];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[2];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[2];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[2];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[2];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[2];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[2];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[2];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[2];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[2];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[2];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[2];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[2];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[2];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[2];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[2];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[2];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[2];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[2];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[2];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[2];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[2];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[2];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[2];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[2];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[2];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[2];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[2];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[2];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[2];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[2];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[2];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[2];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[2];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[2];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[2];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[2];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[2];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[2];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[2];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[2];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[2];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[2];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[2];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[2];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[2];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[2];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[2];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[2];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[2];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[2];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[2];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[2];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[2];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[2];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[2];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[2];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[2];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[2];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[2];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[2];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[2];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[2];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[2];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[2];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[3];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[3];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[3];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[3];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[3];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[3];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[3];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[3];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[3];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[3];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[3];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[3];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[3];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[3];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[3];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[3];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[3];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[3];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[3];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[3];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[3];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[3];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[3];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[3];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[3];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[3];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[3];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[3];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[3];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[3];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[3];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[3];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[3];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[3];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[3];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[3];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[3];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[3];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[3];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[3];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[3];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[3];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[3];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[3];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[3];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[3];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[3];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[3];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[3];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[3];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[3];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[3];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[3];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[3];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[3];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[3];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[3];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[3];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[3];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[3];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[3];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[3];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[3];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[3];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[3];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[3];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[3];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[3];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[3];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[3];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[3];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[3];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[3];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[3];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[3];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[3];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[3];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[3];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[3];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[3];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[3];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[3];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[3];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[3];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[3];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[3];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[3];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[3];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[3];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[3];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[3];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[3];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[3];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[3];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[3];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[3];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[3];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[3];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[3];
  assign data_o[0] = N1 | data_masked[0];
  assign N1 = N0 | data_masked[99];
  assign N0 = data_masked[297] | data_masked[198];
  assign data_o[1] = N3 | data_masked[1];
  assign N3 = N2 | data_masked[100];
  assign N2 = data_masked[298] | data_masked[199];
  assign data_o[2] = N5 | data_masked[2];
  assign N5 = N4 | data_masked[101];
  assign N4 = data_masked[299] | data_masked[200];
  assign data_o[3] = N7 | data_masked[3];
  assign N7 = N6 | data_masked[102];
  assign N6 = data_masked[300] | data_masked[201];
  assign data_o[4] = N9 | data_masked[4];
  assign N9 = N8 | data_masked[103];
  assign N8 = data_masked[301] | data_masked[202];
  assign data_o[5] = N11 | data_masked[5];
  assign N11 = N10 | data_masked[104];
  assign N10 = data_masked[302] | data_masked[203];
  assign data_o[6] = N13 | data_masked[6];
  assign N13 = N12 | data_masked[105];
  assign N12 = data_masked[303] | data_masked[204];
  assign data_o[7] = N15 | data_masked[7];
  assign N15 = N14 | data_masked[106];
  assign N14 = data_masked[304] | data_masked[205];
  assign data_o[8] = N17 | data_masked[8];
  assign N17 = N16 | data_masked[107];
  assign N16 = data_masked[305] | data_masked[206];
  assign data_o[9] = N19 | data_masked[9];
  assign N19 = N18 | data_masked[108];
  assign N18 = data_masked[306] | data_masked[207];
  assign data_o[10] = N21 | data_masked[10];
  assign N21 = N20 | data_masked[109];
  assign N20 = data_masked[307] | data_masked[208];
  assign data_o[11] = N23 | data_masked[11];
  assign N23 = N22 | data_masked[110];
  assign N22 = data_masked[308] | data_masked[209];
  assign data_o[12] = N25 | data_masked[12];
  assign N25 = N24 | data_masked[111];
  assign N24 = data_masked[309] | data_masked[210];
  assign data_o[13] = N27 | data_masked[13];
  assign N27 = N26 | data_masked[112];
  assign N26 = data_masked[310] | data_masked[211];
  assign data_o[14] = N29 | data_masked[14];
  assign N29 = N28 | data_masked[113];
  assign N28 = data_masked[311] | data_masked[212];
  assign data_o[15] = N31 | data_masked[15];
  assign N31 = N30 | data_masked[114];
  assign N30 = data_masked[312] | data_masked[213];
  assign data_o[16] = N33 | data_masked[16];
  assign N33 = N32 | data_masked[115];
  assign N32 = data_masked[313] | data_masked[214];
  assign data_o[17] = N35 | data_masked[17];
  assign N35 = N34 | data_masked[116];
  assign N34 = data_masked[314] | data_masked[215];
  assign data_o[18] = N37 | data_masked[18];
  assign N37 = N36 | data_masked[117];
  assign N36 = data_masked[315] | data_masked[216];
  assign data_o[19] = N39 | data_masked[19];
  assign N39 = N38 | data_masked[118];
  assign N38 = data_masked[316] | data_masked[217];
  assign data_o[20] = N41 | data_masked[20];
  assign N41 = N40 | data_masked[119];
  assign N40 = data_masked[317] | data_masked[218];
  assign data_o[21] = N43 | data_masked[21];
  assign N43 = N42 | data_masked[120];
  assign N42 = data_masked[318] | data_masked[219];
  assign data_o[22] = N45 | data_masked[22];
  assign N45 = N44 | data_masked[121];
  assign N44 = data_masked[319] | data_masked[220];
  assign data_o[23] = N47 | data_masked[23];
  assign N47 = N46 | data_masked[122];
  assign N46 = data_masked[320] | data_masked[221];
  assign data_o[24] = N49 | data_masked[24];
  assign N49 = N48 | data_masked[123];
  assign N48 = data_masked[321] | data_masked[222];
  assign data_o[25] = N51 | data_masked[25];
  assign N51 = N50 | data_masked[124];
  assign N50 = data_masked[322] | data_masked[223];
  assign data_o[26] = N53 | data_masked[26];
  assign N53 = N52 | data_masked[125];
  assign N52 = data_masked[323] | data_masked[224];
  assign data_o[27] = N55 | data_masked[27];
  assign N55 = N54 | data_masked[126];
  assign N54 = data_masked[324] | data_masked[225];
  assign data_o[28] = N57 | data_masked[28];
  assign N57 = N56 | data_masked[127];
  assign N56 = data_masked[325] | data_masked[226];
  assign data_o[29] = N59 | data_masked[29];
  assign N59 = N58 | data_masked[128];
  assign N58 = data_masked[326] | data_masked[227];
  assign data_o[30] = N61 | data_masked[30];
  assign N61 = N60 | data_masked[129];
  assign N60 = data_masked[327] | data_masked[228];
  assign data_o[31] = N63 | data_masked[31];
  assign N63 = N62 | data_masked[130];
  assign N62 = data_masked[328] | data_masked[229];
  assign data_o[32] = N65 | data_masked[32];
  assign N65 = N64 | data_masked[131];
  assign N64 = data_masked[329] | data_masked[230];
  assign data_o[33] = N67 | data_masked[33];
  assign N67 = N66 | data_masked[132];
  assign N66 = data_masked[330] | data_masked[231];
  assign data_o[34] = N69 | data_masked[34];
  assign N69 = N68 | data_masked[133];
  assign N68 = data_masked[331] | data_masked[232];
  assign data_o[35] = N71 | data_masked[35];
  assign N71 = N70 | data_masked[134];
  assign N70 = data_masked[332] | data_masked[233];
  assign data_o[36] = N73 | data_masked[36];
  assign N73 = N72 | data_masked[135];
  assign N72 = data_masked[333] | data_masked[234];
  assign data_o[37] = N75 | data_masked[37];
  assign N75 = N74 | data_masked[136];
  assign N74 = data_masked[334] | data_masked[235];
  assign data_o[38] = N77 | data_masked[38];
  assign N77 = N76 | data_masked[137];
  assign N76 = data_masked[335] | data_masked[236];
  assign data_o[39] = N79 | data_masked[39];
  assign N79 = N78 | data_masked[138];
  assign N78 = data_masked[336] | data_masked[237];
  assign data_o[40] = N81 | data_masked[40];
  assign N81 = N80 | data_masked[139];
  assign N80 = data_masked[337] | data_masked[238];
  assign data_o[41] = N83 | data_masked[41];
  assign N83 = N82 | data_masked[140];
  assign N82 = data_masked[338] | data_masked[239];
  assign data_o[42] = N85 | data_masked[42];
  assign N85 = N84 | data_masked[141];
  assign N84 = data_masked[339] | data_masked[240];
  assign data_o[43] = N87 | data_masked[43];
  assign N87 = N86 | data_masked[142];
  assign N86 = data_masked[340] | data_masked[241];
  assign data_o[44] = N89 | data_masked[44];
  assign N89 = N88 | data_masked[143];
  assign N88 = data_masked[341] | data_masked[242];
  assign data_o[45] = N91 | data_masked[45];
  assign N91 = N90 | data_masked[144];
  assign N90 = data_masked[342] | data_masked[243];
  assign data_o[46] = N93 | data_masked[46];
  assign N93 = N92 | data_masked[145];
  assign N92 = data_masked[343] | data_masked[244];
  assign data_o[47] = N95 | data_masked[47];
  assign N95 = N94 | data_masked[146];
  assign N94 = data_masked[344] | data_masked[245];
  assign data_o[48] = N97 | data_masked[48];
  assign N97 = N96 | data_masked[147];
  assign N96 = data_masked[345] | data_masked[246];
  assign data_o[49] = N99 | data_masked[49];
  assign N99 = N98 | data_masked[148];
  assign N98 = data_masked[346] | data_masked[247];
  assign data_o[50] = N101 | data_masked[50];
  assign N101 = N100 | data_masked[149];
  assign N100 = data_masked[347] | data_masked[248];
  assign data_o[51] = N103 | data_masked[51];
  assign N103 = N102 | data_masked[150];
  assign N102 = data_masked[348] | data_masked[249];
  assign data_o[52] = N105 | data_masked[52];
  assign N105 = N104 | data_masked[151];
  assign N104 = data_masked[349] | data_masked[250];
  assign data_o[53] = N107 | data_masked[53];
  assign N107 = N106 | data_masked[152];
  assign N106 = data_masked[350] | data_masked[251];
  assign data_o[54] = N109 | data_masked[54];
  assign N109 = N108 | data_masked[153];
  assign N108 = data_masked[351] | data_masked[252];
  assign data_o[55] = N111 | data_masked[55];
  assign N111 = N110 | data_masked[154];
  assign N110 = data_masked[352] | data_masked[253];
  assign data_o[56] = N113 | data_masked[56];
  assign N113 = N112 | data_masked[155];
  assign N112 = data_masked[353] | data_masked[254];
  assign data_o[57] = N115 | data_masked[57];
  assign N115 = N114 | data_masked[156];
  assign N114 = data_masked[354] | data_masked[255];
  assign data_o[58] = N117 | data_masked[58];
  assign N117 = N116 | data_masked[157];
  assign N116 = data_masked[355] | data_masked[256];
  assign data_o[59] = N119 | data_masked[59];
  assign N119 = N118 | data_masked[158];
  assign N118 = data_masked[356] | data_masked[257];
  assign data_o[60] = N121 | data_masked[60];
  assign N121 = N120 | data_masked[159];
  assign N120 = data_masked[357] | data_masked[258];
  assign data_o[61] = N123 | data_masked[61];
  assign N123 = N122 | data_masked[160];
  assign N122 = data_masked[358] | data_masked[259];
  assign data_o[62] = N125 | data_masked[62];
  assign N125 = N124 | data_masked[161];
  assign N124 = data_masked[359] | data_masked[260];
  assign data_o[63] = N127 | data_masked[63];
  assign N127 = N126 | data_masked[162];
  assign N126 = data_masked[360] | data_masked[261];
  assign data_o[64] = N129 | data_masked[64];
  assign N129 = N128 | data_masked[163];
  assign N128 = data_masked[361] | data_masked[262];
  assign data_o[65] = N131 | data_masked[65];
  assign N131 = N130 | data_masked[164];
  assign N130 = data_masked[362] | data_masked[263];
  assign data_o[66] = N133 | data_masked[66];
  assign N133 = N132 | data_masked[165];
  assign N132 = data_masked[363] | data_masked[264];
  assign data_o[67] = N135 | data_masked[67];
  assign N135 = N134 | data_masked[166];
  assign N134 = data_masked[364] | data_masked[265];
  assign data_o[68] = N137 | data_masked[68];
  assign N137 = N136 | data_masked[167];
  assign N136 = data_masked[365] | data_masked[266];
  assign data_o[69] = N139 | data_masked[69];
  assign N139 = N138 | data_masked[168];
  assign N138 = data_masked[366] | data_masked[267];
  assign data_o[70] = N141 | data_masked[70];
  assign N141 = N140 | data_masked[169];
  assign N140 = data_masked[367] | data_masked[268];
  assign data_o[71] = N143 | data_masked[71];
  assign N143 = N142 | data_masked[170];
  assign N142 = data_masked[368] | data_masked[269];
  assign data_o[72] = N145 | data_masked[72];
  assign N145 = N144 | data_masked[171];
  assign N144 = data_masked[369] | data_masked[270];
  assign data_o[73] = N147 | data_masked[73];
  assign N147 = N146 | data_masked[172];
  assign N146 = data_masked[370] | data_masked[271];
  assign data_o[74] = N149 | data_masked[74];
  assign N149 = N148 | data_masked[173];
  assign N148 = data_masked[371] | data_masked[272];
  assign data_o[75] = N151 | data_masked[75];
  assign N151 = N150 | data_masked[174];
  assign N150 = data_masked[372] | data_masked[273];
  assign data_o[76] = N153 | data_masked[76];
  assign N153 = N152 | data_masked[175];
  assign N152 = data_masked[373] | data_masked[274];
  assign data_o[77] = N155 | data_masked[77];
  assign N155 = N154 | data_masked[176];
  assign N154 = data_masked[374] | data_masked[275];
  assign data_o[78] = N157 | data_masked[78];
  assign N157 = N156 | data_masked[177];
  assign N156 = data_masked[375] | data_masked[276];
  assign data_o[79] = N159 | data_masked[79];
  assign N159 = N158 | data_masked[178];
  assign N158 = data_masked[376] | data_masked[277];
  assign data_o[80] = N161 | data_masked[80];
  assign N161 = N160 | data_masked[179];
  assign N160 = data_masked[377] | data_masked[278];
  assign data_o[81] = N163 | data_masked[81];
  assign N163 = N162 | data_masked[180];
  assign N162 = data_masked[378] | data_masked[279];
  assign data_o[82] = N165 | data_masked[82];
  assign N165 = N164 | data_masked[181];
  assign N164 = data_masked[379] | data_masked[280];
  assign data_o[83] = N167 | data_masked[83];
  assign N167 = N166 | data_masked[182];
  assign N166 = data_masked[380] | data_masked[281];
  assign data_o[84] = N169 | data_masked[84];
  assign N169 = N168 | data_masked[183];
  assign N168 = data_masked[381] | data_masked[282];
  assign data_o[85] = N171 | data_masked[85];
  assign N171 = N170 | data_masked[184];
  assign N170 = data_masked[382] | data_masked[283];
  assign data_o[86] = N173 | data_masked[86];
  assign N173 = N172 | data_masked[185];
  assign N172 = data_masked[383] | data_masked[284];
  assign data_o[87] = N175 | data_masked[87];
  assign N175 = N174 | data_masked[186];
  assign N174 = data_masked[384] | data_masked[285];
  assign data_o[88] = N177 | data_masked[88];
  assign N177 = N176 | data_masked[187];
  assign N176 = data_masked[385] | data_masked[286];
  assign data_o[89] = N179 | data_masked[89];
  assign N179 = N178 | data_masked[188];
  assign N178 = data_masked[386] | data_masked[287];
  assign data_o[90] = N181 | data_masked[90];
  assign N181 = N180 | data_masked[189];
  assign N180 = data_masked[387] | data_masked[288];
  assign data_o[91] = N183 | data_masked[91];
  assign N183 = N182 | data_masked[190];
  assign N182 = data_masked[388] | data_masked[289];
  assign data_o[92] = N185 | data_masked[92];
  assign N185 = N184 | data_masked[191];
  assign N184 = data_masked[389] | data_masked[290];
  assign data_o[93] = N187 | data_masked[93];
  assign N187 = N186 | data_masked[192];
  assign N186 = data_masked[390] | data_masked[291];
  assign data_o[94] = N189 | data_masked[94];
  assign N189 = N188 | data_masked[193];
  assign N188 = data_masked[391] | data_masked[292];
  assign data_o[95] = N191 | data_masked[95];
  assign N191 = N190 | data_masked[194];
  assign N190 = data_masked[392] | data_masked[293];
  assign data_o[96] = N193 | data_masked[96];
  assign N193 = N192 | data_masked[195];
  assign N192 = data_masked[393] | data_masked[294];
  assign data_o[97] = N195 | data_masked[97];
  assign N195 = N194 | data_masked[196];
  assign N194 = data_masked[394] | data_masked[295];
  assign data_o[98] = N197 | data_masked[98];
  assign N197 = N196 | data_masked[197];
  assign N196 = data_masked[395] | data_masked[296];

endmodule



module bsg_mux_one_hot_width_p99_els_p2
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [197:0] data_i;
  input [1:0] sel_one_hot_i;
  output [98:0] data_o;
  wire [98:0] data_o;
  wire [197:0] data_masked;
  assign data_masked[98] = data_i[98] & sel_one_hot_i[0];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[0];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[0];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[0];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[0];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[0];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[0];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[0];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[0];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[0];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[0];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[0];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[0];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[0];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[0];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[0];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[0];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[0];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[0];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[0];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[0];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[0];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[0];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[0];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[0];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[0];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[0];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[0];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[0];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[0];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[0];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[1];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[1];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[1];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[1];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[1];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[1];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[1];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[1];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[1];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[1];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[1];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[1];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[1];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[1];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[1];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[1];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[1];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[1];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[1];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[1];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[1];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[1];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[1];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[1];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[1];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[1];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[1];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[1];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[1];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[1];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[1];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[1];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[1];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[1];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[1];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[1];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[1];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[1];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[1];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[1];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[1];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[1];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[1];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[1];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[1];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[1];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[1];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[1];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[1];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[1];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[1];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[1];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[1];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[1];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[1];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[1];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[1];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[1];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[1];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[1];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[1];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[1];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[1];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[1];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[1];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[1];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[1];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[1];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[1];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_o[0] = data_masked[99] | data_masked[0];
  assign data_o[1] = data_masked[100] | data_masked[1];
  assign data_o[2] = data_masked[101] | data_masked[2];
  assign data_o[3] = data_masked[102] | data_masked[3];
  assign data_o[4] = data_masked[103] | data_masked[4];
  assign data_o[5] = data_masked[104] | data_masked[5];
  assign data_o[6] = data_masked[105] | data_masked[6];
  assign data_o[7] = data_masked[106] | data_masked[7];
  assign data_o[8] = data_masked[107] | data_masked[8];
  assign data_o[9] = data_masked[108] | data_masked[9];
  assign data_o[10] = data_masked[109] | data_masked[10];
  assign data_o[11] = data_masked[110] | data_masked[11];
  assign data_o[12] = data_masked[111] | data_masked[12];
  assign data_o[13] = data_masked[112] | data_masked[13];
  assign data_o[14] = data_masked[113] | data_masked[14];
  assign data_o[15] = data_masked[114] | data_masked[15];
  assign data_o[16] = data_masked[115] | data_masked[16];
  assign data_o[17] = data_masked[116] | data_masked[17];
  assign data_o[18] = data_masked[117] | data_masked[18];
  assign data_o[19] = data_masked[118] | data_masked[19];
  assign data_o[20] = data_masked[119] | data_masked[20];
  assign data_o[21] = data_masked[120] | data_masked[21];
  assign data_o[22] = data_masked[121] | data_masked[22];
  assign data_o[23] = data_masked[122] | data_masked[23];
  assign data_o[24] = data_masked[123] | data_masked[24];
  assign data_o[25] = data_masked[124] | data_masked[25];
  assign data_o[26] = data_masked[125] | data_masked[26];
  assign data_o[27] = data_masked[126] | data_masked[27];
  assign data_o[28] = data_masked[127] | data_masked[28];
  assign data_o[29] = data_masked[128] | data_masked[29];
  assign data_o[30] = data_masked[129] | data_masked[30];
  assign data_o[31] = data_masked[130] | data_masked[31];
  assign data_o[32] = data_masked[131] | data_masked[32];
  assign data_o[33] = data_masked[132] | data_masked[33];
  assign data_o[34] = data_masked[133] | data_masked[34];
  assign data_o[35] = data_masked[134] | data_masked[35];
  assign data_o[36] = data_masked[135] | data_masked[36];
  assign data_o[37] = data_masked[136] | data_masked[37];
  assign data_o[38] = data_masked[137] | data_masked[38];
  assign data_o[39] = data_masked[138] | data_masked[39];
  assign data_o[40] = data_masked[139] | data_masked[40];
  assign data_o[41] = data_masked[140] | data_masked[41];
  assign data_o[42] = data_masked[141] | data_masked[42];
  assign data_o[43] = data_masked[142] | data_masked[43];
  assign data_o[44] = data_masked[143] | data_masked[44];
  assign data_o[45] = data_masked[144] | data_masked[45];
  assign data_o[46] = data_masked[145] | data_masked[46];
  assign data_o[47] = data_masked[146] | data_masked[47];
  assign data_o[48] = data_masked[147] | data_masked[48];
  assign data_o[49] = data_masked[148] | data_masked[49];
  assign data_o[50] = data_masked[149] | data_masked[50];
  assign data_o[51] = data_masked[150] | data_masked[51];
  assign data_o[52] = data_masked[151] | data_masked[52];
  assign data_o[53] = data_masked[152] | data_masked[53];
  assign data_o[54] = data_masked[153] | data_masked[54];
  assign data_o[55] = data_masked[154] | data_masked[55];
  assign data_o[56] = data_masked[155] | data_masked[56];
  assign data_o[57] = data_masked[156] | data_masked[57];
  assign data_o[58] = data_masked[157] | data_masked[58];
  assign data_o[59] = data_masked[158] | data_masked[59];
  assign data_o[60] = data_masked[159] | data_masked[60];
  assign data_o[61] = data_masked[160] | data_masked[61];
  assign data_o[62] = data_masked[161] | data_masked[62];
  assign data_o[63] = data_masked[162] | data_masked[63];
  assign data_o[64] = data_masked[163] | data_masked[64];
  assign data_o[65] = data_masked[164] | data_masked[65];
  assign data_o[66] = data_masked[165] | data_masked[66];
  assign data_o[67] = data_masked[166] | data_masked[67];
  assign data_o[68] = data_masked[167] | data_masked[68];
  assign data_o[69] = data_masked[168] | data_masked[69];
  assign data_o[70] = data_masked[169] | data_masked[70];
  assign data_o[71] = data_masked[170] | data_masked[71];
  assign data_o[72] = data_masked[171] | data_masked[72];
  assign data_o[73] = data_masked[172] | data_masked[73];
  assign data_o[74] = data_masked[173] | data_masked[74];
  assign data_o[75] = data_masked[174] | data_masked[75];
  assign data_o[76] = data_masked[175] | data_masked[76];
  assign data_o[77] = data_masked[176] | data_masked[77];
  assign data_o[78] = data_masked[177] | data_masked[78];
  assign data_o[79] = data_masked[178] | data_masked[79];
  assign data_o[80] = data_masked[179] | data_masked[80];
  assign data_o[81] = data_masked[180] | data_masked[81];
  assign data_o[82] = data_masked[181] | data_masked[82];
  assign data_o[83] = data_masked[182] | data_masked[83];
  assign data_o[84] = data_masked[183] | data_masked[84];
  assign data_o[85] = data_masked[184] | data_masked[85];
  assign data_o[86] = data_masked[185] | data_masked[86];
  assign data_o[87] = data_masked[186] | data_masked[87];
  assign data_o[88] = data_masked[187] | data_masked[88];
  assign data_o[89] = data_masked[188] | data_masked[89];
  assign data_o[90] = data_masked[189] | data_masked[90];
  assign data_o[91] = data_masked[190] | data_masked[91];
  assign data_o[92] = data_masked[191] | data_masked[92];
  assign data_o[93] = data_masked[192] | data_masked[93];
  assign data_o[94] = data_masked[193] | data_masked[94];
  assign data_o[95] = data_masked[194] | data_masked[95];
  assign data_o[96] = data_masked[195] | data_masked[96];
  assign data_o[97] = data_masked[196] | data_masked[97];
  assign data_o[98] = data_masked[197] | data_masked[98];

endmodule



module bsg_mux_one_hot_width_p99_els_p5
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [494:0] data_i;
  input [4:0] sel_one_hot_i;
  output [98:0] data_o;
  wire [98:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296;
  wire [494:0] data_masked;
  assign data_masked[98] = data_i[98] & sel_one_hot_i[0];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[0];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[0];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[0];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[0];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[0];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[0];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[0];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[0];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[0];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[0];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[0];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[0];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[0];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[0];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[0];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[0];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[0];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[0];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[0];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[0];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[0];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[0];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[0];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[0];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[0];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[0];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[0];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[0];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[0];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[0];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[1];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[1];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[1];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[1];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[1];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[1];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[1];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[1];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[1];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[1];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[1];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[1];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[1];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[1];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[1];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[1];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[1];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[1];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[1];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[1];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[1];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[1];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[1];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[1];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[1];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[1];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[1];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[1];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[1];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[1];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[1];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[1];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[1];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[1];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[1];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[1];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[1];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[1];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[1];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[1];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[1];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[1];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[1];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[1];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[1];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[1];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[1];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[1];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[1];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[1];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[1];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[1];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[1];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[1];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[1];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[1];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[1];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[1];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[1];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[1];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[1];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[1];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[1];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[1];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[1];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[1];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[1];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[1];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[1];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[1];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[1];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[1];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[1];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[2];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[2];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[2];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[2];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[2];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[2];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[2];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[2];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[2];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[2];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[2];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[2];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[2];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[2];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[2];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[2];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[2];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[2];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[2];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[2];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[2];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[2];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[2];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[2];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[2];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[2];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[2];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[2];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[2];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[2];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[2];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[2];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[2];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[2];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[2];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[2];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[2];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[2];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[2];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[2];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[2];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[2];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[2];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[2];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[2];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[2];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[2];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[2];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[2];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[2];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[2];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[2];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[2];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[2];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[2];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[2];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[2];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[2];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[2];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[2];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[2];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[2];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[2];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[2];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[2];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[2];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[2];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[2];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[2];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[2];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[2];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[2];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[2];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[2];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[2];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[2];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[2];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[2];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[2];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[2];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[2];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[2];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[2];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[2];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[2];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[2];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[2];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[2];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[2];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[2];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[2];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[2];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[2];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[2];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[2];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[2];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[2];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[2];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[2];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[3];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[3];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[3];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[3];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[3];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[3];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[3];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[3];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[3];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[3];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[3];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[3];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[3];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[3];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[3];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[3];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[3];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[3];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[3];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[3];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[3];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[3];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[3];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[3];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[3];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[3];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[3];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[3];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[3];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[3];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[3];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[3];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[3];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[3];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[3];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[3];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[3];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[3];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[3];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[3];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[3];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[3];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[3];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[3];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[3];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[3];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[3];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[3];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[3];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[3];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[3];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[3];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[3];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[3];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[3];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[3];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[3];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[3];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[3];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[3];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[3];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[3];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[3];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[3];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[3];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[3];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[3];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[3];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[3];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[3];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[3];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[3];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[3];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[3];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[3];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[3];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[3];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[3];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[3];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[3];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[3];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[3];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[3];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[3];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[3];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[3];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[3];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[3];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[3];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[3];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[3];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[3];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[3];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[3];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[3];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[3];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[3];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[3];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[3];
  assign data_masked[494] = data_i[494] & sel_one_hot_i[4];
  assign data_masked[493] = data_i[493] & sel_one_hot_i[4];
  assign data_masked[492] = data_i[492] & sel_one_hot_i[4];
  assign data_masked[491] = data_i[491] & sel_one_hot_i[4];
  assign data_masked[490] = data_i[490] & sel_one_hot_i[4];
  assign data_masked[489] = data_i[489] & sel_one_hot_i[4];
  assign data_masked[488] = data_i[488] & sel_one_hot_i[4];
  assign data_masked[487] = data_i[487] & sel_one_hot_i[4];
  assign data_masked[486] = data_i[486] & sel_one_hot_i[4];
  assign data_masked[485] = data_i[485] & sel_one_hot_i[4];
  assign data_masked[484] = data_i[484] & sel_one_hot_i[4];
  assign data_masked[483] = data_i[483] & sel_one_hot_i[4];
  assign data_masked[482] = data_i[482] & sel_one_hot_i[4];
  assign data_masked[481] = data_i[481] & sel_one_hot_i[4];
  assign data_masked[480] = data_i[480] & sel_one_hot_i[4];
  assign data_masked[479] = data_i[479] & sel_one_hot_i[4];
  assign data_masked[478] = data_i[478] & sel_one_hot_i[4];
  assign data_masked[477] = data_i[477] & sel_one_hot_i[4];
  assign data_masked[476] = data_i[476] & sel_one_hot_i[4];
  assign data_masked[475] = data_i[475] & sel_one_hot_i[4];
  assign data_masked[474] = data_i[474] & sel_one_hot_i[4];
  assign data_masked[473] = data_i[473] & sel_one_hot_i[4];
  assign data_masked[472] = data_i[472] & sel_one_hot_i[4];
  assign data_masked[471] = data_i[471] & sel_one_hot_i[4];
  assign data_masked[470] = data_i[470] & sel_one_hot_i[4];
  assign data_masked[469] = data_i[469] & sel_one_hot_i[4];
  assign data_masked[468] = data_i[468] & sel_one_hot_i[4];
  assign data_masked[467] = data_i[467] & sel_one_hot_i[4];
  assign data_masked[466] = data_i[466] & sel_one_hot_i[4];
  assign data_masked[465] = data_i[465] & sel_one_hot_i[4];
  assign data_masked[464] = data_i[464] & sel_one_hot_i[4];
  assign data_masked[463] = data_i[463] & sel_one_hot_i[4];
  assign data_masked[462] = data_i[462] & sel_one_hot_i[4];
  assign data_masked[461] = data_i[461] & sel_one_hot_i[4];
  assign data_masked[460] = data_i[460] & sel_one_hot_i[4];
  assign data_masked[459] = data_i[459] & sel_one_hot_i[4];
  assign data_masked[458] = data_i[458] & sel_one_hot_i[4];
  assign data_masked[457] = data_i[457] & sel_one_hot_i[4];
  assign data_masked[456] = data_i[456] & sel_one_hot_i[4];
  assign data_masked[455] = data_i[455] & sel_one_hot_i[4];
  assign data_masked[454] = data_i[454] & sel_one_hot_i[4];
  assign data_masked[453] = data_i[453] & sel_one_hot_i[4];
  assign data_masked[452] = data_i[452] & sel_one_hot_i[4];
  assign data_masked[451] = data_i[451] & sel_one_hot_i[4];
  assign data_masked[450] = data_i[450] & sel_one_hot_i[4];
  assign data_masked[449] = data_i[449] & sel_one_hot_i[4];
  assign data_masked[448] = data_i[448] & sel_one_hot_i[4];
  assign data_masked[447] = data_i[447] & sel_one_hot_i[4];
  assign data_masked[446] = data_i[446] & sel_one_hot_i[4];
  assign data_masked[445] = data_i[445] & sel_one_hot_i[4];
  assign data_masked[444] = data_i[444] & sel_one_hot_i[4];
  assign data_masked[443] = data_i[443] & sel_one_hot_i[4];
  assign data_masked[442] = data_i[442] & sel_one_hot_i[4];
  assign data_masked[441] = data_i[441] & sel_one_hot_i[4];
  assign data_masked[440] = data_i[440] & sel_one_hot_i[4];
  assign data_masked[439] = data_i[439] & sel_one_hot_i[4];
  assign data_masked[438] = data_i[438] & sel_one_hot_i[4];
  assign data_masked[437] = data_i[437] & sel_one_hot_i[4];
  assign data_masked[436] = data_i[436] & sel_one_hot_i[4];
  assign data_masked[435] = data_i[435] & sel_one_hot_i[4];
  assign data_masked[434] = data_i[434] & sel_one_hot_i[4];
  assign data_masked[433] = data_i[433] & sel_one_hot_i[4];
  assign data_masked[432] = data_i[432] & sel_one_hot_i[4];
  assign data_masked[431] = data_i[431] & sel_one_hot_i[4];
  assign data_masked[430] = data_i[430] & sel_one_hot_i[4];
  assign data_masked[429] = data_i[429] & sel_one_hot_i[4];
  assign data_masked[428] = data_i[428] & sel_one_hot_i[4];
  assign data_masked[427] = data_i[427] & sel_one_hot_i[4];
  assign data_masked[426] = data_i[426] & sel_one_hot_i[4];
  assign data_masked[425] = data_i[425] & sel_one_hot_i[4];
  assign data_masked[424] = data_i[424] & sel_one_hot_i[4];
  assign data_masked[423] = data_i[423] & sel_one_hot_i[4];
  assign data_masked[422] = data_i[422] & sel_one_hot_i[4];
  assign data_masked[421] = data_i[421] & sel_one_hot_i[4];
  assign data_masked[420] = data_i[420] & sel_one_hot_i[4];
  assign data_masked[419] = data_i[419] & sel_one_hot_i[4];
  assign data_masked[418] = data_i[418] & sel_one_hot_i[4];
  assign data_masked[417] = data_i[417] & sel_one_hot_i[4];
  assign data_masked[416] = data_i[416] & sel_one_hot_i[4];
  assign data_masked[415] = data_i[415] & sel_one_hot_i[4];
  assign data_masked[414] = data_i[414] & sel_one_hot_i[4];
  assign data_masked[413] = data_i[413] & sel_one_hot_i[4];
  assign data_masked[412] = data_i[412] & sel_one_hot_i[4];
  assign data_masked[411] = data_i[411] & sel_one_hot_i[4];
  assign data_masked[410] = data_i[410] & sel_one_hot_i[4];
  assign data_masked[409] = data_i[409] & sel_one_hot_i[4];
  assign data_masked[408] = data_i[408] & sel_one_hot_i[4];
  assign data_masked[407] = data_i[407] & sel_one_hot_i[4];
  assign data_masked[406] = data_i[406] & sel_one_hot_i[4];
  assign data_masked[405] = data_i[405] & sel_one_hot_i[4];
  assign data_masked[404] = data_i[404] & sel_one_hot_i[4];
  assign data_masked[403] = data_i[403] & sel_one_hot_i[4];
  assign data_masked[402] = data_i[402] & sel_one_hot_i[4];
  assign data_masked[401] = data_i[401] & sel_one_hot_i[4];
  assign data_masked[400] = data_i[400] & sel_one_hot_i[4];
  assign data_masked[399] = data_i[399] & sel_one_hot_i[4];
  assign data_masked[398] = data_i[398] & sel_one_hot_i[4];
  assign data_masked[397] = data_i[397] & sel_one_hot_i[4];
  assign data_masked[396] = data_i[396] & sel_one_hot_i[4];
  assign data_o[0] = N2 | data_masked[0];
  assign N2 = N1 | data_masked[99];
  assign N1 = N0 | data_masked[198];
  assign N0 = data_masked[396] | data_masked[297];
  assign data_o[1] = N5 | data_masked[1];
  assign N5 = N4 | data_masked[100];
  assign N4 = N3 | data_masked[199];
  assign N3 = data_masked[397] | data_masked[298];
  assign data_o[2] = N8 | data_masked[2];
  assign N8 = N7 | data_masked[101];
  assign N7 = N6 | data_masked[200];
  assign N6 = data_masked[398] | data_masked[299];
  assign data_o[3] = N11 | data_masked[3];
  assign N11 = N10 | data_masked[102];
  assign N10 = N9 | data_masked[201];
  assign N9 = data_masked[399] | data_masked[300];
  assign data_o[4] = N14 | data_masked[4];
  assign N14 = N13 | data_masked[103];
  assign N13 = N12 | data_masked[202];
  assign N12 = data_masked[400] | data_masked[301];
  assign data_o[5] = N17 | data_masked[5];
  assign N17 = N16 | data_masked[104];
  assign N16 = N15 | data_masked[203];
  assign N15 = data_masked[401] | data_masked[302];
  assign data_o[6] = N20 | data_masked[6];
  assign N20 = N19 | data_masked[105];
  assign N19 = N18 | data_masked[204];
  assign N18 = data_masked[402] | data_masked[303];
  assign data_o[7] = N23 | data_masked[7];
  assign N23 = N22 | data_masked[106];
  assign N22 = N21 | data_masked[205];
  assign N21 = data_masked[403] | data_masked[304];
  assign data_o[8] = N26 | data_masked[8];
  assign N26 = N25 | data_masked[107];
  assign N25 = N24 | data_masked[206];
  assign N24 = data_masked[404] | data_masked[305];
  assign data_o[9] = N29 | data_masked[9];
  assign N29 = N28 | data_masked[108];
  assign N28 = N27 | data_masked[207];
  assign N27 = data_masked[405] | data_masked[306];
  assign data_o[10] = N32 | data_masked[10];
  assign N32 = N31 | data_masked[109];
  assign N31 = N30 | data_masked[208];
  assign N30 = data_masked[406] | data_masked[307];
  assign data_o[11] = N35 | data_masked[11];
  assign N35 = N34 | data_masked[110];
  assign N34 = N33 | data_masked[209];
  assign N33 = data_masked[407] | data_masked[308];
  assign data_o[12] = N38 | data_masked[12];
  assign N38 = N37 | data_masked[111];
  assign N37 = N36 | data_masked[210];
  assign N36 = data_masked[408] | data_masked[309];
  assign data_o[13] = N41 | data_masked[13];
  assign N41 = N40 | data_masked[112];
  assign N40 = N39 | data_masked[211];
  assign N39 = data_masked[409] | data_masked[310];
  assign data_o[14] = N44 | data_masked[14];
  assign N44 = N43 | data_masked[113];
  assign N43 = N42 | data_masked[212];
  assign N42 = data_masked[410] | data_masked[311];
  assign data_o[15] = N47 | data_masked[15];
  assign N47 = N46 | data_masked[114];
  assign N46 = N45 | data_masked[213];
  assign N45 = data_masked[411] | data_masked[312];
  assign data_o[16] = N50 | data_masked[16];
  assign N50 = N49 | data_masked[115];
  assign N49 = N48 | data_masked[214];
  assign N48 = data_masked[412] | data_masked[313];
  assign data_o[17] = N53 | data_masked[17];
  assign N53 = N52 | data_masked[116];
  assign N52 = N51 | data_masked[215];
  assign N51 = data_masked[413] | data_masked[314];
  assign data_o[18] = N56 | data_masked[18];
  assign N56 = N55 | data_masked[117];
  assign N55 = N54 | data_masked[216];
  assign N54 = data_masked[414] | data_masked[315];
  assign data_o[19] = N59 | data_masked[19];
  assign N59 = N58 | data_masked[118];
  assign N58 = N57 | data_masked[217];
  assign N57 = data_masked[415] | data_masked[316];
  assign data_o[20] = N62 | data_masked[20];
  assign N62 = N61 | data_masked[119];
  assign N61 = N60 | data_masked[218];
  assign N60 = data_masked[416] | data_masked[317];
  assign data_o[21] = N65 | data_masked[21];
  assign N65 = N64 | data_masked[120];
  assign N64 = N63 | data_masked[219];
  assign N63 = data_masked[417] | data_masked[318];
  assign data_o[22] = N68 | data_masked[22];
  assign N68 = N67 | data_masked[121];
  assign N67 = N66 | data_masked[220];
  assign N66 = data_masked[418] | data_masked[319];
  assign data_o[23] = N71 | data_masked[23];
  assign N71 = N70 | data_masked[122];
  assign N70 = N69 | data_masked[221];
  assign N69 = data_masked[419] | data_masked[320];
  assign data_o[24] = N74 | data_masked[24];
  assign N74 = N73 | data_masked[123];
  assign N73 = N72 | data_masked[222];
  assign N72 = data_masked[420] | data_masked[321];
  assign data_o[25] = N77 | data_masked[25];
  assign N77 = N76 | data_masked[124];
  assign N76 = N75 | data_masked[223];
  assign N75 = data_masked[421] | data_masked[322];
  assign data_o[26] = N80 | data_masked[26];
  assign N80 = N79 | data_masked[125];
  assign N79 = N78 | data_masked[224];
  assign N78 = data_masked[422] | data_masked[323];
  assign data_o[27] = N83 | data_masked[27];
  assign N83 = N82 | data_masked[126];
  assign N82 = N81 | data_masked[225];
  assign N81 = data_masked[423] | data_masked[324];
  assign data_o[28] = N86 | data_masked[28];
  assign N86 = N85 | data_masked[127];
  assign N85 = N84 | data_masked[226];
  assign N84 = data_masked[424] | data_masked[325];
  assign data_o[29] = N89 | data_masked[29];
  assign N89 = N88 | data_masked[128];
  assign N88 = N87 | data_masked[227];
  assign N87 = data_masked[425] | data_masked[326];
  assign data_o[30] = N92 | data_masked[30];
  assign N92 = N91 | data_masked[129];
  assign N91 = N90 | data_masked[228];
  assign N90 = data_masked[426] | data_masked[327];
  assign data_o[31] = N95 | data_masked[31];
  assign N95 = N94 | data_masked[130];
  assign N94 = N93 | data_masked[229];
  assign N93 = data_masked[427] | data_masked[328];
  assign data_o[32] = N98 | data_masked[32];
  assign N98 = N97 | data_masked[131];
  assign N97 = N96 | data_masked[230];
  assign N96 = data_masked[428] | data_masked[329];
  assign data_o[33] = N101 | data_masked[33];
  assign N101 = N100 | data_masked[132];
  assign N100 = N99 | data_masked[231];
  assign N99 = data_masked[429] | data_masked[330];
  assign data_o[34] = N104 | data_masked[34];
  assign N104 = N103 | data_masked[133];
  assign N103 = N102 | data_masked[232];
  assign N102 = data_masked[430] | data_masked[331];
  assign data_o[35] = N107 | data_masked[35];
  assign N107 = N106 | data_masked[134];
  assign N106 = N105 | data_masked[233];
  assign N105 = data_masked[431] | data_masked[332];
  assign data_o[36] = N110 | data_masked[36];
  assign N110 = N109 | data_masked[135];
  assign N109 = N108 | data_masked[234];
  assign N108 = data_masked[432] | data_masked[333];
  assign data_o[37] = N113 | data_masked[37];
  assign N113 = N112 | data_masked[136];
  assign N112 = N111 | data_masked[235];
  assign N111 = data_masked[433] | data_masked[334];
  assign data_o[38] = N116 | data_masked[38];
  assign N116 = N115 | data_masked[137];
  assign N115 = N114 | data_masked[236];
  assign N114 = data_masked[434] | data_masked[335];
  assign data_o[39] = N119 | data_masked[39];
  assign N119 = N118 | data_masked[138];
  assign N118 = N117 | data_masked[237];
  assign N117 = data_masked[435] | data_masked[336];
  assign data_o[40] = N122 | data_masked[40];
  assign N122 = N121 | data_masked[139];
  assign N121 = N120 | data_masked[238];
  assign N120 = data_masked[436] | data_masked[337];
  assign data_o[41] = N125 | data_masked[41];
  assign N125 = N124 | data_masked[140];
  assign N124 = N123 | data_masked[239];
  assign N123 = data_masked[437] | data_masked[338];
  assign data_o[42] = N128 | data_masked[42];
  assign N128 = N127 | data_masked[141];
  assign N127 = N126 | data_masked[240];
  assign N126 = data_masked[438] | data_masked[339];
  assign data_o[43] = N131 | data_masked[43];
  assign N131 = N130 | data_masked[142];
  assign N130 = N129 | data_masked[241];
  assign N129 = data_masked[439] | data_masked[340];
  assign data_o[44] = N134 | data_masked[44];
  assign N134 = N133 | data_masked[143];
  assign N133 = N132 | data_masked[242];
  assign N132 = data_masked[440] | data_masked[341];
  assign data_o[45] = N137 | data_masked[45];
  assign N137 = N136 | data_masked[144];
  assign N136 = N135 | data_masked[243];
  assign N135 = data_masked[441] | data_masked[342];
  assign data_o[46] = N140 | data_masked[46];
  assign N140 = N139 | data_masked[145];
  assign N139 = N138 | data_masked[244];
  assign N138 = data_masked[442] | data_masked[343];
  assign data_o[47] = N143 | data_masked[47];
  assign N143 = N142 | data_masked[146];
  assign N142 = N141 | data_masked[245];
  assign N141 = data_masked[443] | data_masked[344];
  assign data_o[48] = N146 | data_masked[48];
  assign N146 = N145 | data_masked[147];
  assign N145 = N144 | data_masked[246];
  assign N144 = data_masked[444] | data_masked[345];
  assign data_o[49] = N149 | data_masked[49];
  assign N149 = N148 | data_masked[148];
  assign N148 = N147 | data_masked[247];
  assign N147 = data_masked[445] | data_masked[346];
  assign data_o[50] = N152 | data_masked[50];
  assign N152 = N151 | data_masked[149];
  assign N151 = N150 | data_masked[248];
  assign N150 = data_masked[446] | data_masked[347];
  assign data_o[51] = N155 | data_masked[51];
  assign N155 = N154 | data_masked[150];
  assign N154 = N153 | data_masked[249];
  assign N153 = data_masked[447] | data_masked[348];
  assign data_o[52] = N158 | data_masked[52];
  assign N158 = N157 | data_masked[151];
  assign N157 = N156 | data_masked[250];
  assign N156 = data_masked[448] | data_masked[349];
  assign data_o[53] = N161 | data_masked[53];
  assign N161 = N160 | data_masked[152];
  assign N160 = N159 | data_masked[251];
  assign N159 = data_masked[449] | data_masked[350];
  assign data_o[54] = N164 | data_masked[54];
  assign N164 = N163 | data_masked[153];
  assign N163 = N162 | data_masked[252];
  assign N162 = data_masked[450] | data_masked[351];
  assign data_o[55] = N167 | data_masked[55];
  assign N167 = N166 | data_masked[154];
  assign N166 = N165 | data_masked[253];
  assign N165 = data_masked[451] | data_masked[352];
  assign data_o[56] = N170 | data_masked[56];
  assign N170 = N169 | data_masked[155];
  assign N169 = N168 | data_masked[254];
  assign N168 = data_masked[452] | data_masked[353];
  assign data_o[57] = N173 | data_masked[57];
  assign N173 = N172 | data_masked[156];
  assign N172 = N171 | data_masked[255];
  assign N171 = data_masked[453] | data_masked[354];
  assign data_o[58] = N176 | data_masked[58];
  assign N176 = N175 | data_masked[157];
  assign N175 = N174 | data_masked[256];
  assign N174 = data_masked[454] | data_masked[355];
  assign data_o[59] = N179 | data_masked[59];
  assign N179 = N178 | data_masked[158];
  assign N178 = N177 | data_masked[257];
  assign N177 = data_masked[455] | data_masked[356];
  assign data_o[60] = N182 | data_masked[60];
  assign N182 = N181 | data_masked[159];
  assign N181 = N180 | data_masked[258];
  assign N180 = data_masked[456] | data_masked[357];
  assign data_o[61] = N185 | data_masked[61];
  assign N185 = N184 | data_masked[160];
  assign N184 = N183 | data_masked[259];
  assign N183 = data_masked[457] | data_masked[358];
  assign data_o[62] = N188 | data_masked[62];
  assign N188 = N187 | data_masked[161];
  assign N187 = N186 | data_masked[260];
  assign N186 = data_masked[458] | data_masked[359];
  assign data_o[63] = N191 | data_masked[63];
  assign N191 = N190 | data_masked[162];
  assign N190 = N189 | data_masked[261];
  assign N189 = data_masked[459] | data_masked[360];
  assign data_o[64] = N194 | data_masked[64];
  assign N194 = N193 | data_masked[163];
  assign N193 = N192 | data_masked[262];
  assign N192 = data_masked[460] | data_masked[361];
  assign data_o[65] = N197 | data_masked[65];
  assign N197 = N196 | data_masked[164];
  assign N196 = N195 | data_masked[263];
  assign N195 = data_masked[461] | data_masked[362];
  assign data_o[66] = N200 | data_masked[66];
  assign N200 = N199 | data_masked[165];
  assign N199 = N198 | data_masked[264];
  assign N198 = data_masked[462] | data_masked[363];
  assign data_o[67] = N203 | data_masked[67];
  assign N203 = N202 | data_masked[166];
  assign N202 = N201 | data_masked[265];
  assign N201 = data_masked[463] | data_masked[364];
  assign data_o[68] = N206 | data_masked[68];
  assign N206 = N205 | data_masked[167];
  assign N205 = N204 | data_masked[266];
  assign N204 = data_masked[464] | data_masked[365];
  assign data_o[69] = N209 | data_masked[69];
  assign N209 = N208 | data_masked[168];
  assign N208 = N207 | data_masked[267];
  assign N207 = data_masked[465] | data_masked[366];
  assign data_o[70] = N212 | data_masked[70];
  assign N212 = N211 | data_masked[169];
  assign N211 = N210 | data_masked[268];
  assign N210 = data_masked[466] | data_masked[367];
  assign data_o[71] = N215 | data_masked[71];
  assign N215 = N214 | data_masked[170];
  assign N214 = N213 | data_masked[269];
  assign N213 = data_masked[467] | data_masked[368];
  assign data_o[72] = N218 | data_masked[72];
  assign N218 = N217 | data_masked[171];
  assign N217 = N216 | data_masked[270];
  assign N216 = data_masked[468] | data_masked[369];
  assign data_o[73] = N221 | data_masked[73];
  assign N221 = N220 | data_masked[172];
  assign N220 = N219 | data_masked[271];
  assign N219 = data_masked[469] | data_masked[370];
  assign data_o[74] = N224 | data_masked[74];
  assign N224 = N223 | data_masked[173];
  assign N223 = N222 | data_masked[272];
  assign N222 = data_masked[470] | data_masked[371];
  assign data_o[75] = N227 | data_masked[75];
  assign N227 = N226 | data_masked[174];
  assign N226 = N225 | data_masked[273];
  assign N225 = data_masked[471] | data_masked[372];
  assign data_o[76] = N230 | data_masked[76];
  assign N230 = N229 | data_masked[175];
  assign N229 = N228 | data_masked[274];
  assign N228 = data_masked[472] | data_masked[373];
  assign data_o[77] = N233 | data_masked[77];
  assign N233 = N232 | data_masked[176];
  assign N232 = N231 | data_masked[275];
  assign N231 = data_masked[473] | data_masked[374];
  assign data_o[78] = N236 | data_masked[78];
  assign N236 = N235 | data_masked[177];
  assign N235 = N234 | data_masked[276];
  assign N234 = data_masked[474] | data_masked[375];
  assign data_o[79] = N239 | data_masked[79];
  assign N239 = N238 | data_masked[178];
  assign N238 = N237 | data_masked[277];
  assign N237 = data_masked[475] | data_masked[376];
  assign data_o[80] = N242 | data_masked[80];
  assign N242 = N241 | data_masked[179];
  assign N241 = N240 | data_masked[278];
  assign N240 = data_masked[476] | data_masked[377];
  assign data_o[81] = N245 | data_masked[81];
  assign N245 = N244 | data_masked[180];
  assign N244 = N243 | data_masked[279];
  assign N243 = data_masked[477] | data_masked[378];
  assign data_o[82] = N248 | data_masked[82];
  assign N248 = N247 | data_masked[181];
  assign N247 = N246 | data_masked[280];
  assign N246 = data_masked[478] | data_masked[379];
  assign data_o[83] = N251 | data_masked[83];
  assign N251 = N250 | data_masked[182];
  assign N250 = N249 | data_masked[281];
  assign N249 = data_masked[479] | data_masked[380];
  assign data_o[84] = N254 | data_masked[84];
  assign N254 = N253 | data_masked[183];
  assign N253 = N252 | data_masked[282];
  assign N252 = data_masked[480] | data_masked[381];
  assign data_o[85] = N257 | data_masked[85];
  assign N257 = N256 | data_masked[184];
  assign N256 = N255 | data_masked[283];
  assign N255 = data_masked[481] | data_masked[382];
  assign data_o[86] = N260 | data_masked[86];
  assign N260 = N259 | data_masked[185];
  assign N259 = N258 | data_masked[284];
  assign N258 = data_masked[482] | data_masked[383];
  assign data_o[87] = N263 | data_masked[87];
  assign N263 = N262 | data_masked[186];
  assign N262 = N261 | data_masked[285];
  assign N261 = data_masked[483] | data_masked[384];
  assign data_o[88] = N266 | data_masked[88];
  assign N266 = N265 | data_masked[187];
  assign N265 = N264 | data_masked[286];
  assign N264 = data_masked[484] | data_masked[385];
  assign data_o[89] = N269 | data_masked[89];
  assign N269 = N268 | data_masked[188];
  assign N268 = N267 | data_masked[287];
  assign N267 = data_masked[485] | data_masked[386];
  assign data_o[90] = N272 | data_masked[90];
  assign N272 = N271 | data_masked[189];
  assign N271 = N270 | data_masked[288];
  assign N270 = data_masked[486] | data_masked[387];
  assign data_o[91] = N275 | data_masked[91];
  assign N275 = N274 | data_masked[190];
  assign N274 = N273 | data_masked[289];
  assign N273 = data_masked[487] | data_masked[388];
  assign data_o[92] = N278 | data_masked[92];
  assign N278 = N277 | data_masked[191];
  assign N277 = N276 | data_masked[290];
  assign N276 = data_masked[488] | data_masked[389];
  assign data_o[93] = N281 | data_masked[93];
  assign N281 = N280 | data_masked[192];
  assign N280 = N279 | data_masked[291];
  assign N279 = data_masked[489] | data_masked[390];
  assign data_o[94] = N284 | data_masked[94];
  assign N284 = N283 | data_masked[193];
  assign N283 = N282 | data_masked[292];
  assign N282 = data_masked[490] | data_masked[391];
  assign data_o[95] = N287 | data_masked[95];
  assign N287 = N286 | data_masked[194];
  assign N286 = N285 | data_masked[293];
  assign N285 = data_masked[491] | data_masked[392];
  assign data_o[96] = N290 | data_masked[96];
  assign N290 = N289 | data_masked[195];
  assign N289 = N288 | data_masked[294];
  assign N288 = data_masked[492] | data_masked[393];
  assign data_o[97] = N293 | data_masked[97];
  assign N293 = N292 | data_masked[196];
  assign N292 = N291 | data_masked[295];
  assign N291 = data_masked[493] | data_masked[394];
  assign data_o[98] = N296 | data_masked[98];
  assign N296 = N295 | data_masked[197];
  assign N295 = N294 | data_masked[296];
  assign N294 = data_masked[494] | data_masked[395];

endmodule



module bsg_mesh_router_99_1_1_0_0a_0
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  yumi_o,
  ready_i,
  data_o,
  v_o,
  my_x_i,
  my_y_i
);

  input [494:0] data_i;
  input [4:0] v_i;
  output [4:0] yumi_o;
  input [4:0] ready_i;
  output [494:0] data_o;
  output [4:0] v_o;
  input [0:0] my_x_i;
  input [0:0] my_y_i;
  input clk_i;
  input reset_i;
  wire [4:0] yumi_o,v_o;
  wire [494:0] data_o;
  wire n_3_net_,W_sel_e,W_sel_p,W_sel_n,W_sel_s,W_gnt_e,W_gnt_p,W_gnt_n,W_gnt_s,
  n_9_net_,E_sel_w,E_sel_p,E_sel_n,E_sel_s,E_gnt_w,E_gnt_p,E_gnt_n,E_gnt_s,n_15_net_,
  N_sel_s,N_sel_p,N_gnt_s,N_gnt_p,n_21_net_,S_sel_n,S_sel_p,S_gnt_n,S_gnt_p,n_27_net_,
  P_sel_s,P_sel_n,P_sel_e,P_sel_w,P_sel_p,P_gnt_s,P_gnt_n,P_gnt_e,P_gnt_w,P_gnt_p,
  N0,N1,N2,N3,N4,N5,N6,SV2V_UNCONNECTED_1,SV2V_UNCONNECTED_2,
  SV2V_UNCONNECTED_3,SV2V_UNCONNECTED_4,SV2V_UNCONNECTED_5,SV2V_UNCONNECTED_6,
  SV2V_UNCONNECTED_7,SV2V_UNCONNECTED_8,SV2V_UNCONNECTED_9;
  wire [24:0] req;

  bsg_mesh_router_dor_decoder_x_cord_width_p1_y_cord_width_p1_dirs_lp5_XY_order_p0
  dor_decoder
  (
    .clk_i(clk_i),
    .v_i({ v_i[4:4], 1'b0, v_i[2:2], 1'b0, v_i[0:0] }),
    .x_dirs_i({ data_i[396:396], data_i[297:297], data_i[198:198], data_i[99:99], data_i[0:0] }),
    .y_dirs_i({ data_i[397:397], data_i[298:298], data_i[199:199], data_i[100:100], data_i[1:1] }),
    .my_x_i(my_x_i[0]),
    .my_y_i(my_y_i[0]),
    .req_o(req)
  );


  bsg_round_robin_arb_inputs_p4
  genblk2_west_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ req[11:11], req[1:1], req[16:16], req[21:21] }),
    .grants_o({ W_gnt_e, W_gnt_p, W_gnt_n, W_gnt_s }),
    .sel_one_hot_o({ W_sel_e, W_sel_p, W_sel_n, W_sel_s }),
    .v_o(v_o[1]),
    .tag_o({ SV2V_UNCONNECTED_1, SV2V_UNCONNECTED_2 }),
    .yumi_i(n_3_net_)
  );


  bsg_mux_one_hot_width_p99_els_p4
  genblk2_mux_data_west
  (
    .data_i({ data_i[98:0], data_i[296:198], data_i[395:297], data_i[494:396] }),
    .sel_one_hot_i({ W_sel_p, W_sel_e, W_sel_n, W_sel_s }),
    .data_o(data_o[197:99])
  );


  bsg_round_robin_arb_inputs_p4
  genblk3_east_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[2]),
    .reqs_i({ req[7:7], req[2:2], req[17:17], req[22:22] }),
    .grants_o({ E_gnt_w, E_gnt_p, E_gnt_n, E_gnt_s }),
    .sel_one_hot_o({ E_sel_w, E_sel_p, E_sel_n, E_sel_s }),
    .v_o(v_o[2]),
    .tag_o({ SV2V_UNCONNECTED_3, SV2V_UNCONNECTED_4 }),
    .yumi_i(n_9_net_)
  );


  bsg_mux_one_hot_width_p99_els_p4
  genblk3_mux_data_east
  (
    .data_i({ data_i[98:0], data_i[197:99], data_i[395:297], data_i[494:396] }),
    .sel_one_hot_i({ E_sel_p, E_sel_w, E_sel_n, E_sel_s }),
    .data_o(data_o[296:198])
  );


  bsg_round_robin_arb_inputs_p2
  genblk4_north_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ req[23:23], req[3:3] }),
    .grants_o({ N_gnt_s, N_gnt_p }),
    .sel_one_hot_o({ N_sel_s, N_sel_p }),
    .v_o(v_o[3]),
    .tag_o(SV2V_UNCONNECTED_5),
    .yumi_i(n_15_net_)
  );


  bsg_mux_one_hot_width_p99_els_p2
  genblk4_mux_data_north
  (
    .data_i({ data_i[98:0], data_i[494:396] }),
    .sel_one_hot_i({ N_sel_p, N_sel_s }),
    .data_o(data_o[395:297])
  );


  bsg_round_robin_arb_inputs_p2
  genblk5_south_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[4]),
    .reqs_i({ req[19:19], req[4:4] }),
    .grants_o({ S_gnt_n, S_gnt_p }),
    .sel_one_hot_o({ S_sel_n, S_sel_p }),
    .v_o(v_o[4]),
    .tag_o(SV2V_UNCONNECTED_6),
    .yumi_i(n_21_net_)
  );


  bsg_mux_one_hot_width_p99_els_p2
  genblk5_mux_data_south
  (
    .data_i({ data_i[98:0], data_i[395:297] }),
    .sel_one_hot_i({ S_sel_p, S_sel_n }),
    .data_o(data_o[494:396])
  );


  bsg_round_robin_arb_inputs_p5
  proc_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[0]),
    .reqs_i({ req[20:20], req[15:15], req[10:10], req[5:5], req[0:0] }),
    .grants_o({ P_gnt_s, P_gnt_n, P_gnt_e, P_gnt_w, P_gnt_p }),
    .sel_one_hot_o({ P_sel_s, P_sel_n, P_sel_e, P_sel_w, P_sel_p }),
    .v_o(v_o[0]),
    .tag_o({ SV2V_UNCONNECTED_7, SV2V_UNCONNECTED_8, SV2V_UNCONNECTED_9 }),
    .yumi_i(n_27_net_)
  );


  bsg_mux_one_hot_width_p99_els_p5
  mux_data_proc
  (
    .data_i({ data_i[98:0], data_i[296:198], data_i[494:396], data_i[197:99], data_i[395:297] }),
    .sel_one_hot_i({ P_sel_p, P_sel_e, P_sel_s, P_sel_w, P_sel_n }),
    .data_o(data_o[98:0])
  );

  assign n_3_net_ = v_o[1] & 1'b1;
  assign n_9_net_ = v_o[2] & ready_i[2];
  assign n_15_net_ = v_o[3] & 1'b1;
  assign n_21_net_ = v_o[4] & ready_i[4];
  assign n_27_net_ = v_o[0] & ready_i[0];
  assign yumi_o[0] = N2 | W_gnt_p;
  assign N2 = N1 | P_gnt_p;
  assign N1 = N0 | S_gnt_p;
  assign N0 = E_gnt_p | N_gnt_p;
  assign yumi_o[1] = E_gnt_w | P_gnt_w;
  assign yumi_o[2] = W_gnt_e | P_gnt_e;
  assign yumi_o[3] = N4 | P_gnt_n;
  assign N4 = N3 | E_gnt_n;
  assign N3 = S_gnt_n | W_gnt_n;
  assign yumi_o[4] = N6 | P_gnt_s;
  assign N6 = N5 | E_gnt_s;
  assign N5 = N_gnt_s | W_gnt_s;

endmodule



module bsg_mesh_router_buffered_99_1_1_0_5_0a_0_101_00
(
  clk_i,
  reset_i,
  link_i,
  link_o,
  my_x_i,
  my_y_i
);

  input [504:0] link_i;
  output [504:0] link_o;
  input [0:0] my_x_i;
  input [0:0] my_y_i;
  input clk_i;
  input reset_i;
  wire [504:0] link_o;
  wire fifo_valid_2,fifo_valid_0,fifo_data_4__98_,fifo_data_4__97_,fifo_data_4__96_,
  fifo_data_4__95_,fifo_data_4__94_,fifo_data_4__93_,fifo_data_4__92_,
  fifo_data_4__91_,fifo_data_4__90_,fifo_data_4__89_,fifo_data_4__88_,fifo_data_4__87_,
  fifo_data_4__86_,fifo_data_4__85_,fifo_data_4__84_,fifo_data_4__83_,fifo_data_4__82_,
  fifo_data_4__81_,fifo_data_4__80_,fifo_data_4__79_,fifo_data_4__78_,fifo_data_4__77_,
  fifo_data_4__76_,fifo_data_4__75_,fifo_data_4__74_,fifo_data_4__73_,
  fifo_data_4__72_,fifo_data_4__71_,fifo_data_4__70_,fifo_data_4__69_,fifo_data_4__68_,
  fifo_data_4__67_,fifo_data_4__66_,fifo_data_4__65_,fifo_data_4__64_,fifo_data_4__63_,
  fifo_data_4__62_,fifo_data_4__61_,fifo_data_4__60_,fifo_data_4__59_,
  fifo_data_4__58_,fifo_data_4__57_,fifo_data_4__56_,fifo_data_4__55_,fifo_data_4__54_,
  fifo_data_4__53_,fifo_data_4__52_,fifo_data_4__51_,fifo_data_4__50_,fifo_data_4__49_,
  fifo_data_4__48_,fifo_data_4__47_,fifo_data_4__46_,fifo_data_4__45_,
  fifo_data_4__44_,fifo_data_4__43_,fifo_data_4__42_,fifo_data_4__41_,fifo_data_4__40_,
  fifo_data_4__39_,fifo_data_4__38_,fifo_data_4__37_,fifo_data_4__36_,fifo_data_4__35_,
  fifo_data_4__34_,fifo_data_4__33_,fifo_data_4__32_,fifo_data_4__31_,fifo_data_4__30_,
  fifo_data_4__29_,fifo_data_4__28_,fifo_data_4__27_,fifo_data_4__26_,
  fifo_data_4__25_,fifo_data_4__24_,fifo_data_4__23_,fifo_data_4__22_,fifo_data_4__21_,
  fifo_data_4__20_,fifo_data_4__19_,fifo_data_4__18_,fifo_data_4__17_,fifo_data_4__16_,
  fifo_data_4__15_,fifo_data_4__14_,fifo_data_4__13_,fifo_data_4__12_,
  fifo_data_4__11_,fifo_data_4__10_,fifo_data_4__9_,fifo_data_4__8_,fifo_data_4__7_,
  fifo_data_4__6_,fifo_data_4__5_,fifo_data_4__4_,fifo_data_4__3_,fifo_data_4__2_,
  fifo_data_4__1_,fifo_data_4__0_,fifo_data_2__98_,fifo_data_2__97_,fifo_data_2__96_,
  fifo_data_2__95_,fifo_data_2__94_,fifo_data_2__93_,fifo_data_2__92_,fifo_data_2__91_,
  fifo_data_2__90_,fifo_data_2__89_,fifo_data_2__88_,fifo_data_2__87_,fifo_data_2__86_,
  fifo_data_2__85_,fifo_data_2__84_,fifo_data_2__83_,fifo_data_2__82_,
  fifo_data_2__81_,fifo_data_2__80_,fifo_data_2__79_,fifo_data_2__78_,fifo_data_2__77_,
  fifo_data_2__76_,fifo_data_2__75_,fifo_data_2__74_,fifo_data_2__73_,fifo_data_2__72_,
  fifo_data_2__71_,fifo_data_2__70_,fifo_data_2__69_,fifo_data_2__68_,
  fifo_data_2__67_,fifo_data_2__66_,fifo_data_2__65_,fifo_data_2__64_,fifo_data_2__63_,
  fifo_data_2__62_,fifo_data_2__61_,fifo_data_2__60_,fifo_data_2__59_,fifo_data_2__58_,
  fifo_data_2__57_,fifo_data_2__56_,fifo_data_2__55_,fifo_data_2__54_,
  fifo_data_2__53_,fifo_data_2__52_,fifo_data_2__51_,fifo_data_2__50_,fifo_data_2__49_,
  fifo_data_2__48_,fifo_data_2__47_,fifo_data_2__46_,fifo_data_2__45_,fifo_data_2__44_,
  fifo_data_2__43_,fifo_data_2__42_,fifo_data_2__41_,fifo_data_2__40_,fifo_data_2__39_,
  fifo_data_2__38_,fifo_data_2__37_,fifo_data_2__36_,fifo_data_2__35_,
  fifo_data_2__34_,fifo_data_2__33_,fifo_data_2__32_,fifo_data_2__31_,fifo_data_2__30_,
  fifo_data_2__29_,fifo_data_2__28_,fifo_data_2__27_,fifo_data_2__26_,fifo_data_2__25_,
  fifo_data_2__24_,fifo_data_2__23_,fifo_data_2__22_,fifo_data_2__21_,
  fifo_data_2__20_,fifo_data_2__19_,fifo_data_2__18_,fifo_data_2__17_,fifo_data_2__16_,
  fifo_data_2__15_,fifo_data_2__14_,fifo_data_2__13_,fifo_data_2__12_,fifo_data_2__11_,
  fifo_data_2__10_,fifo_data_2__9_,fifo_data_2__8_,fifo_data_2__7_,fifo_data_2__6_,
  fifo_data_2__5_,fifo_data_2__4_,fifo_data_2__3_,fifo_data_2__2_,fifo_data_2__1_,
  fifo_data_2__0_,fifo_data_0__98_,fifo_data_0__97_,fifo_data_0__96_,fifo_data_0__95_,
  fifo_data_0__94_,fifo_data_0__93_,fifo_data_0__92_,fifo_data_0__91_,
  fifo_data_0__90_,fifo_data_0__89_,fifo_data_0__88_,fifo_data_0__87_,fifo_data_0__86_,
  fifo_data_0__85_,fifo_data_0__84_,fifo_data_0__83_,fifo_data_0__82_,fifo_data_0__81_,
  fifo_data_0__80_,fifo_data_0__79_,fifo_data_0__78_,fifo_data_0__77_,
  fifo_data_0__76_,fifo_data_0__75_,fifo_data_0__74_,fifo_data_0__73_,fifo_data_0__72_,
  fifo_data_0__71_,fifo_data_0__70_,fifo_data_0__69_,fifo_data_0__68_,fifo_data_0__67_,
  fifo_data_0__66_,fifo_data_0__65_,fifo_data_0__64_,fifo_data_0__63_,
  fifo_data_0__62_,fifo_data_0__61_,fifo_data_0__60_,fifo_data_0__59_,fifo_data_0__58_,
  fifo_data_0__57_,fifo_data_0__56_,fifo_data_0__55_,fifo_data_0__54_,fifo_data_0__53_,
  fifo_data_0__52_,fifo_data_0__51_,fifo_data_0__50_,fifo_data_0__49_,fifo_data_0__48_,
  fifo_data_0__47_,fifo_data_0__46_,fifo_data_0__45_,fifo_data_0__44_,
  fifo_data_0__43_,fifo_data_0__42_,fifo_data_0__41_,fifo_data_0__40_,fifo_data_0__39_,
  fifo_data_0__38_,fifo_data_0__37_,fifo_data_0__36_,fifo_data_0__35_,fifo_data_0__34_,
  fifo_data_0__33_,fifo_data_0__32_,fifo_data_0__31_,fifo_data_0__30_,
  fifo_data_0__29_,fifo_data_0__28_,fifo_data_0__27_,fifo_data_0__26_,fifo_data_0__25_,
  fifo_data_0__24_,fifo_data_0__23_,fifo_data_0__22_,fifo_data_0__21_,fifo_data_0__20_,
  fifo_data_0__19_,fifo_data_0__18_,fifo_data_0__17_,fifo_data_0__16_,fifo_data_0__15_,
  fifo_data_0__14_,fifo_data_0__13_,fifo_data_0__12_,fifo_data_0__11_,
  fifo_data_0__10_,fifo_data_0__9_,fifo_data_0__8_,fifo_data_0__7_,fifo_data_0__6_,
  fifo_data_0__5_,fifo_data_0__4_,fifo_data_0__3_,fifo_data_0__2_,fifo_data_0__1_,
  fifo_data_0__0_;
  wire [4:4] fifo_valid;
  wire [4:0] fifo_yumi;
  assign link_o[200] = 1'b0;
  assign link_o[402] = 1'b0;

  bsg_two_fifo_width_p99
  rof_0__fi_twofer
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(link_o[99]),
    .data_i(link_i[98:0]),
    .v_i(link_i[100]),
    .v_o(fifo_valid_0),
    .data_o({ fifo_data_0__98_, fifo_data_0__97_, fifo_data_0__96_, fifo_data_0__95_, fifo_data_0__94_, fifo_data_0__93_, fifo_data_0__92_, fifo_data_0__91_, fifo_data_0__90_, fifo_data_0__89_, fifo_data_0__88_, fifo_data_0__87_, fifo_data_0__86_, fifo_data_0__85_, fifo_data_0__84_, fifo_data_0__83_, fifo_data_0__82_, fifo_data_0__81_, fifo_data_0__80_, fifo_data_0__79_, fifo_data_0__78_, fifo_data_0__77_, fifo_data_0__76_, fifo_data_0__75_, fifo_data_0__74_, fifo_data_0__73_, fifo_data_0__72_, fifo_data_0__71_, fifo_data_0__70_, fifo_data_0__69_, fifo_data_0__68_, fifo_data_0__67_, fifo_data_0__66_, fifo_data_0__65_, fifo_data_0__64_, fifo_data_0__63_, fifo_data_0__62_, fifo_data_0__61_, fifo_data_0__60_, fifo_data_0__59_, fifo_data_0__58_, fifo_data_0__57_, fifo_data_0__56_, fifo_data_0__55_, fifo_data_0__54_, fifo_data_0__53_, fifo_data_0__52_, fifo_data_0__51_, fifo_data_0__50_, fifo_data_0__49_, fifo_data_0__48_, fifo_data_0__47_, fifo_data_0__46_, fifo_data_0__45_, fifo_data_0__44_, fifo_data_0__43_, fifo_data_0__42_, fifo_data_0__41_, fifo_data_0__40_, fifo_data_0__39_, fifo_data_0__38_, fifo_data_0__37_, fifo_data_0__36_, fifo_data_0__35_, fifo_data_0__34_, fifo_data_0__33_, fifo_data_0__32_, fifo_data_0__31_, fifo_data_0__30_, fifo_data_0__29_, fifo_data_0__28_, fifo_data_0__27_, fifo_data_0__26_, fifo_data_0__25_, fifo_data_0__24_, fifo_data_0__23_, fifo_data_0__22_, fifo_data_0__21_, fifo_data_0__20_, fifo_data_0__19_, fifo_data_0__18_, fifo_data_0__17_, fifo_data_0__16_, fifo_data_0__15_, fifo_data_0__14_, fifo_data_0__13_, fifo_data_0__12_, fifo_data_0__11_, fifo_data_0__10_, fifo_data_0__9_, fifo_data_0__8_, fifo_data_0__7_, fifo_data_0__6_, fifo_data_0__5_, fifo_data_0__4_, fifo_data_0__3_, fifo_data_0__2_, fifo_data_0__1_, fifo_data_0__0_ }),
    .yumi_i(fifo_yumi[0])
  );


  bsg_two_fifo_width_p99
  rof_2__fi_twofer
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(link_o[301]),
    .data_i(link_i[300:202]),
    .v_i(link_i[302]),
    .v_o(fifo_valid_2),
    .data_o({ fifo_data_2__98_, fifo_data_2__97_, fifo_data_2__96_, fifo_data_2__95_, fifo_data_2__94_, fifo_data_2__93_, fifo_data_2__92_, fifo_data_2__91_, fifo_data_2__90_, fifo_data_2__89_, fifo_data_2__88_, fifo_data_2__87_, fifo_data_2__86_, fifo_data_2__85_, fifo_data_2__84_, fifo_data_2__83_, fifo_data_2__82_, fifo_data_2__81_, fifo_data_2__80_, fifo_data_2__79_, fifo_data_2__78_, fifo_data_2__77_, fifo_data_2__76_, fifo_data_2__75_, fifo_data_2__74_, fifo_data_2__73_, fifo_data_2__72_, fifo_data_2__71_, fifo_data_2__70_, fifo_data_2__69_, fifo_data_2__68_, fifo_data_2__67_, fifo_data_2__66_, fifo_data_2__65_, fifo_data_2__64_, fifo_data_2__63_, fifo_data_2__62_, fifo_data_2__61_, fifo_data_2__60_, fifo_data_2__59_, fifo_data_2__58_, fifo_data_2__57_, fifo_data_2__56_, fifo_data_2__55_, fifo_data_2__54_, fifo_data_2__53_, fifo_data_2__52_, fifo_data_2__51_, fifo_data_2__50_, fifo_data_2__49_, fifo_data_2__48_, fifo_data_2__47_, fifo_data_2__46_, fifo_data_2__45_, fifo_data_2__44_, fifo_data_2__43_, fifo_data_2__42_, fifo_data_2__41_, fifo_data_2__40_, fifo_data_2__39_, fifo_data_2__38_, fifo_data_2__37_, fifo_data_2__36_, fifo_data_2__35_, fifo_data_2__34_, fifo_data_2__33_, fifo_data_2__32_, fifo_data_2__31_, fifo_data_2__30_, fifo_data_2__29_, fifo_data_2__28_, fifo_data_2__27_, fifo_data_2__26_, fifo_data_2__25_, fifo_data_2__24_, fifo_data_2__23_, fifo_data_2__22_, fifo_data_2__21_, fifo_data_2__20_, fifo_data_2__19_, fifo_data_2__18_, fifo_data_2__17_, fifo_data_2__16_, fifo_data_2__15_, fifo_data_2__14_, fifo_data_2__13_, fifo_data_2__12_, fifo_data_2__11_, fifo_data_2__10_, fifo_data_2__9_, fifo_data_2__8_, fifo_data_2__7_, fifo_data_2__6_, fifo_data_2__5_, fifo_data_2__4_, fifo_data_2__3_, fifo_data_2__2_, fifo_data_2__1_, fifo_data_2__0_ }),
    .yumi_i(fifo_yumi[2])
  );


  bsg_two_fifo_width_p99
  rof_4__fi_twofer
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(link_o[503]),
    .data_i(link_i[502:404]),
    .v_i(link_i[504]),
    .v_o(fifo_valid[4]),
    .data_o({ fifo_data_4__98_, fifo_data_4__97_, fifo_data_4__96_, fifo_data_4__95_, fifo_data_4__94_, fifo_data_4__93_, fifo_data_4__92_, fifo_data_4__91_, fifo_data_4__90_, fifo_data_4__89_, fifo_data_4__88_, fifo_data_4__87_, fifo_data_4__86_, fifo_data_4__85_, fifo_data_4__84_, fifo_data_4__83_, fifo_data_4__82_, fifo_data_4__81_, fifo_data_4__80_, fifo_data_4__79_, fifo_data_4__78_, fifo_data_4__77_, fifo_data_4__76_, fifo_data_4__75_, fifo_data_4__74_, fifo_data_4__73_, fifo_data_4__72_, fifo_data_4__71_, fifo_data_4__70_, fifo_data_4__69_, fifo_data_4__68_, fifo_data_4__67_, fifo_data_4__66_, fifo_data_4__65_, fifo_data_4__64_, fifo_data_4__63_, fifo_data_4__62_, fifo_data_4__61_, fifo_data_4__60_, fifo_data_4__59_, fifo_data_4__58_, fifo_data_4__57_, fifo_data_4__56_, fifo_data_4__55_, fifo_data_4__54_, fifo_data_4__53_, fifo_data_4__52_, fifo_data_4__51_, fifo_data_4__50_, fifo_data_4__49_, fifo_data_4__48_, fifo_data_4__47_, fifo_data_4__46_, fifo_data_4__45_, fifo_data_4__44_, fifo_data_4__43_, fifo_data_4__42_, fifo_data_4__41_, fifo_data_4__40_, fifo_data_4__39_, fifo_data_4__38_, fifo_data_4__37_, fifo_data_4__36_, fifo_data_4__35_, fifo_data_4__34_, fifo_data_4__33_, fifo_data_4__32_, fifo_data_4__31_, fifo_data_4__30_, fifo_data_4__29_, fifo_data_4__28_, fifo_data_4__27_, fifo_data_4__26_, fifo_data_4__25_, fifo_data_4__24_, fifo_data_4__23_, fifo_data_4__22_, fifo_data_4__21_, fifo_data_4__20_, fifo_data_4__19_, fifo_data_4__18_, fifo_data_4__17_, fifo_data_4__16_, fifo_data_4__15_, fifo_data_4__14_, fifo_data_4__13_, fifo_data_4__12_, fifo_data_4__11_, fifo_data_4__10_, fifo_data_4__9_, fifo_data_4__8_, fifo_data_4__7_, fifo_data_4__6_, fifo_data_4__5_, fifo_data_4__4_, fifo_data_4__3_, fifo_data_4__2_, fifo_data_4__1_, fifo_data_4__0_ }),
    .yumi_i(fifo_yumi[4])
  );


  bsg_mesh_router_99_1_1_0_0a_0
  bmr
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ fifo_data_4__98_, fifo_data_4__97_, fifo_data_4__96_, fifo_data_4__95_, fifo_data_4__94_, fifo_data_4__93_, fifo_data_4__92_, fifo_data_4__91_, fifo_data_4__90_, fifo_data_4__89_, fifo_data_4__88_, fifo_data_4__87_, fifo_data_4__86_, fifo_data_4__85_, fifo_data_4__84_, fifo_data_4__83_, fifo_data_4__82_, fifo_data_4__81_, fifo_data_4__80_, fifo_data_4__79_, fifo_data_4__78_, fifo_data_4__77_, fifo_data_4__76_, fifo_data_4__75_, fifo_data_4__74_, fifo_data_4__73_, fifo_data_4__72_, fifo_data_4__71_, fifo_data_4__70_, fifo_data_4__69_, fifo_data_4__68_, fifo_data_4__67_, fifo_data_4__66_, fifo_data_4__65_, fifo_data_4__64_, fifo_data_4__63_, fifo_data_4__62_, fifo_data_4__61_, fifo_data_4__60_, fifo_data_4__59_, fifo_data_4__58_, fifo_data_4__57_, fifo_data_4__56_, fifo_data_4__55_, fifo_data_4__54_, fifo_data_4__53_, fifo_data_4__52_, fifo_data_4__51_, fifo_data_4__50_, fifo_data_4__49_, fifo_data_4__48_, fifo_data_4__47_, fifo_data_4__46_, fifo_data_4__45_, fifo_data_4__44_, fifo_data_4__43_, fifo_data_4__42_, fifo_data_4__41_, fifo_data_4__40_, fifo_data_4__39_, fifo_data_4__38_, fifo_data_4__37_, fifo_data_4__36_, fifo_data_4__35_, fifo_data_4__34_, fifo_data_4__33_, fifo_data_4__32_, fifo_data_4__31_, fifo_data_4__30_, fifo_data_4__29_, fifo_data_4__28_, fifo_data_4__27_, fifo_data_4__26_, fifo_data_4__25_, fifo_data_4__24_, fifo_data_4__23_, fifo_data_4__22_, fifo_data_4__21_, fifo_data_4__20_, fifo_data_4__19_, fifo_data_4__18_, fifo_data_4__17_, fifo_data_4__16_, fifo_data_4__15_, fifo_data_4__14_, fifo_data_4__13_, fifo_data_4__12_, fifo_data_4__11_, fifo_data_4__10_, fifo_data_4__9_, fifo_data_4__8_, fifo_data_4__7_, fifo_data_4__6_, fifo_data_4__5_, fifo_data_4__4_, fifo_data_4__3_, fifo_data_4__2_, fifo_data_4__1_, fifo_data_4__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_2__98_, fifo_data_2__97_, fifo_data_2__96_, fifo_data_2__95_, fifo_data_2__94_, fifo_data_2__93_, fifo_data_2__92_, fifo_data_2__91_, fifo_data_2__90_, fifo_data_2__89_, fifo_data_2__88_, fifo_data_2__87_, fifo_data_2__86_, fifo_data_2__85_, fifo_data_2__84_, fifo_data_2__83_, fifo_data_2__82_, fifo_data_2__81_, fifo_data_2__80_, fifo_data_2__79_, fifo_data_2__78_, fifo_data_2__77_, fifo_data_2__76_, fifo_data_2__75_, fifo_data_2__74_, fifo_data_2__73_, fifo_data_2__72_, fifo_data_2__71_, fifo_data_2__70_, fifo_data_2__69_, fifo_data_2__68_, fifo_data_2__67_, fifo_data_2__66_, fifo_data_2__65_, fifo_data_2__64_, fifo_data_2__63_, fifo_data_2__62_, fifo_data_2__61_, fifo_data_2__60_, fifo_data_2__59_, fifo_data_2__58_, fifo_data_2__57_, fifo_data_2__56_, fifo_data_2__55_, fifo_data_2__54_, fifo_data_2__53_, fifo_data_2__52_, fifo_data_2__51_, fifo_data_2__50_, fifo_data_2__49_, fifo_data_2__48_, fifo_data_2__47_, fifo_data_2__46_, fifo_data_2__45_, fifo_data_2__44_, fifo_data_2__43_, fifo_data_2__42_, fifo_data_2__41_, fifo_data_2__40_, fifo_data_2__39_, fifo_data_2__38_, fifo_data_2__37_, fifo_data_2__36_, fifo_data_2__35_, fifo_data_2__34_, fifo_data_2__33_, fifo_data_2__32_, fifo_data_2__31_, fifo_data_2__30_, fifo_data_2__29_, fifo_data_2__28_, fifo_data_2__27_, fifo_data_2__26_, fifo_data_2__25_, fifo_data_2__24_, fifo_data_2__23_, fifo_data_2__22_, fifo_data_2__21_, fifo_data_2__20_, fifo_data_2__19_, fifo_data_2__18_, fifo_data_2__17_, fifo_data_2__16_, fifo_data_2__15_, fifo_data_2__14_, fifo_data_2__13_, fifo_data_2__12_, fifo_data_2__11_, fifo_data_2__10_, fifo_data_2__9_, fifo_data_2__8_, fifo_data_2__7_, fifo_data_2__6_, fifo_data_2__5_, fifo_data_2__4_, fifo_data_2__3_, fifo_data_2__2_, fifo_data_2__1_, fifo_data_2__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_0__98_, fifo_data_0__97_, fifo_data_0__96_, fifo_data_0__95_, fifo_data_0__94_, fifo_data_0__93_, fifo_data_0__92_, fifo_data_0__91_, fifo_data_0__90_, fifo_data_0__89_, fifo_data_0__88_, fifo_data_0__87_, fifo_data_0__86_, fifo_data_0__85_, fifo_data_0__84_, fifo_data_0__83_, fifo_data_0__82_, fifo_data_0__81_, fifo_data_0__80_, fifo_data_0__79_, fifo_data_0__78_, fifo_data_0__77_, fifo_data_0__76_, fifo_data_0__75_, fifo_data_0__74_, fifo_data_0__73_, fifo_data_0__72_, fifo_data_0__71_, fifo_data_0__70_, fifo_data_0__69_, fifo_data_0__68_, fifo_data_0__67_, fifo_data_0__66_, fifo_data_0__65_, fifo_data_0__64_, fifo_data_0__63_, fifo_data_0__62_, fifo_data_0__61_, fifo_data_0__60_, fifo_data_0__59_, fifo_data_0__58_, fifo_data_0__57_, fifo_data_0__56_, fifo_data_0__55_, fifo_data_0__54_, fifo_data_0__53_, fifo_data_0__52_, fifo_data_0__51_, fifo_data_0__50_, fifo_data_0__49_, fifo_data_0__48_, fifo_data_0__47_, fifo_data_0__46_, fifo_data_0__45_, fifo_data_0__44_, fifo_data_0__43_, fifo_data_0__42_, fifo_data_0__41_, fifo_data_0__40_, fifo_data_0__39_, fifo_data_0__38_, fifo_data_0__37_, fifo_data_0__36_, fifo_data_0__35_, fifo_data_0__34_, fifo_data_0__33_, fifo_data_0__32_, fifo_data_0__31_, fifo_data_0__30_, fifo_data_0__29_, fifo_data_0__28_, fifo_data_0__27_, fifo_data_0__26_, fifo_data_0__25_, fifo_data_0__24_, fifo_data_0__23_, fifo_data_0__22_, fifo_data_0__21_, fifo_data_0__20_, fifo_data_0__19_, fifo_data_0__18_, fifo_data_0__17_, fifo_data_0__16_, fifo_data_0__15_, fifo_data_0__14_, fifo_data_0__13_, fifo_data_0__12_, fifo_data_0__11_, fifo_data_0__10_, fifo_data_0__9_, fifo_data_0__8_, fifo_data_0__7_, fifo_data_0__6_, fifo_data_0__5_, fifo_data_0__4_, fifo_data_0__3_, fifo_data_0__2_, fifo_data_0__1_, fifo_data_0__0_ }),
    .v_i({ fifo_valid[4:4], 1'b0, fifo_valid_2, 1'b0, fifo_valid_0 }),
    .yumi_o(fifo_yumi),
    .ready_i({ link_i[503:503], link_i[402:402], link_i[301:301], link_i[200:200], link_i[99:99] }),
    .data_o({ link_o[502:404], link_o[401:303], link_o[300:202], link_o[199:101], link_o[98:0] }),
    .v_o({ link_o[504:504], link_o[403:403], link_o[302:302], link_o[201:201], link_o[100:100] }),
    .my_x_i(my_x_i[0]),
    .my_y_i(my_y_i[0])
  );


endmodule



module bsg_mesh_router_99_1_1_0_0d_0
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  yumi_o,
  ready_i,
  data_o,
  v_o,
  my_x_i,
  my_y_i
);

  input [494:0] data_i;
  input [4:0] v_i;
  output [4:0] yumi_o;
  input [4:0] ready_i;
  output [494:0] data_o;
  output [4:0] v_o;
  input [0:0] my_x_i;
  input [0:0] my_y_i;
  input clk_i;
  input reset_i;
  wire [4:0] yumi_o,v_o;
  wire [494:0] data_o;
  wire n_3_net_,W_sel_e,W_sel_p,W_sel_n,W_sel_s,W_gnt_e,W_gnt_p,W_gnt_n,W_gnt_s,
  n_9_net_,E_sel_w,E_sel_p,E_sel_n,E_sel_s,E_gnt_w,E_gnt_p,E_gnt_n,E_gnt_s,n_15_net_,
  N_sel_s,N_sel_p,N_gnt_s,N_gnt_p,n_21_net_,S_sel_n,S_sel_p,S_gnt_n,S_gnt_p,n_27_net_,
  P_sel_s,P_sel_n,P_sel_e,P_sel_w,P_sel_p,P_gnt_s,P_gnt_n,P_gnt_e,P_gnt_w,P_gnt_p,
  N0,N1,N2,N3,N4,N5,N6,SV2V_UNCONNECTED_1,SV2V_UNCONNECTED_2,
  SV2V_UNCONNECTED_3,SV2V_UNCONNECTED_4,SV2V_UNCONNECTED_5,SV2V_UNCONNECTED_6,
  SV2V_UNCONNECTED_7,SV2V_UNCONNECTED_8,SV2V_UNCONNECTED_9;
  wire [24:0] req;

  bsg_mesh_router_dor_decoder_x_cord_width_p1_y_cord_width_p1_dirs_lp5_XY_order_p0
  dor_decoder
  (
    .clk_i(clk_i),
    .v_i({ v_i[4:4], 1'b0, 1'b0, v_i[1:1], 1'b0 }),
    .x_dirs_i({ data_i[396:396], data_i[297:297], data_i[198:198], data_i[99:99], data_i[0:0] }),
    .y_dirs_i({ data_i[397:397], data_i[298:298], data_i[199:199], data_i[100:100], data_i[1:1] }),
    .my_x_i(my_x_i[0]),
    .my_y_i(my_y_i[0]),
    .req_o(req)
  );


  bsg_round_robin_arb_inputs_p4
  genblk2_west_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[1]),
    .reqs_i({ req[11:11], req[1:1], req[16:16], req[21:21] }),
    .grants_o({ W_gnt_e, W_gnt_p, W_gnt_n, W_gnt_s }),
    .sel_one_hot_o({ W_sel_e, W_sel_p, W_sel_n, W_sel_s }),
    .v_o(v_o[1]),
    .tag_o({ SV2V_UNCONNECTED_1, SV2V_UNCONNECTED_2 }),
    .yumi_i(n_3_net_)
  );


  bsg_mux_one_hot_width_p99_els_p4
  genblk2_mux_data_west
  (
    .data_i({ data_i[98:0], data_i[296:198], data_i[395:297], data_i[494:396] }),
    .sel_one_hot_i({ W_sel_p, W_sel_e, W_sel_n, W_sel_s }),
    .data_o(data_o[197:99])
  );


  bsg_round_robin_arb_inputs_p4
  genblk3_east_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ req[7:7], req[2:2], req[17:17], req[22:22] }),
    .grants_o({ E_gnt_w, E_gnt_p, E_gnt_n, E_gnt_s }),
    .sel_one_hot_o({ E_sel_w, E_sel_p, E_sel_n, E_sel_s }),
    .v_o(v_o[2]),
    .tag_o({ SV2V_UNCONNECTED_3, SV2V_UNCONNECTED_4 }),
    .yumi_i(n_9_net_)
  );


  bsg_mux_one_hot_width_p99_els_p4
  genblk3_mux_data_east
  (
    .data_i({ data_i[98:0], data_i[197:99], data_i[395:297], data_i[494:396] }),
    .sel_one_hot_i({ E_sel_p, E_sel_w, E_sel_n, E_sel_s }),
    .data_o(data_o[296:198])
  );


  bsg_round_robin_arb_inputs_p2
  genblk4_north_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ req[23:23], req[3:3] }),
    .grants_o({ N_gnt_s, N_gnt_p }),
    .sel_one_hot_o({ N_sel_s, N_sel_p }),
    .v_o(v_o[3]),
    .tag_o(SV2V_UNCONNECTED_5),
    .yumi_i(n_15_net_)
  );


  bsg_mux_one_hot_width_p99_els_p2
  genblk4_mux_data_north
  (
    .data_i({ data_i[98:0], data_i[494:396] }),
    .sel_one_hot_i({ N_sel_p, N_sel_s }),
    .data_o(data_o[395:297])
  );


  bsg_round_robin_arb_inputs_p2
  genblk5_south_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[4]),
    .reqs_i({ req[19:19], req[4:4] }),
    .grants_o({ S_gnt_n, S_gnt_p }),
    .sel_one_hot_o({ S_sel_n, S_sel_p }),
    .v_o(v_o[4]),
    .tag_o(SV2V_UNCONNECTED_6),
    .yumi_i(n_21_net_)
  );


  bsg_mux_one_hot_width_p99_els_p2
  genblk5_mux_data_south
  (
    .data_i({ data_i[98:0], data_i[395:297] }),
    .sel_one_hot_i({ S_sel_p, S_sel_n }),
    .data_o(data_o[494:396])
  );


  bsg_round_robin_arb_inputs_p5
  proc_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ req[20:20], req[15:15], req[10:10], req[5:5], req[0:0] }),
    .grants_o({ P_gnt_s, P_gnt_n, P_gnt_e, P_gnt_w, P_gnt_p }),
    .sel_one_hot_o({ P_sel_s, P_sel_n, P_sel_e, P_sel_w, P_sel_p }),
    .v_o(v_o[0]),
    .tag_o({ SV2V_UNCONNECTED_7, SV2V_UNCONNECTED_8, SV2V_UNCONNECTED_9 }),
    .yumi_i(n_27_net_)
  );


  bsg_mux_one_hot_width_p99_els_p5
  mux_data_proc
  (
    .data_i({ data_i[98:0], data_i[296:198], data_i[494:396], data_i[197:99], data_i[395:297] }),
    .sel_one_hot_i({ P_sel_p, P_sel_e, P_sel_s, P_sel_w, P_sel_n }),
    .data_o(data_o[98:0])
  );

  assign n_3_net_ = v_o[1] & ready_i[1];
  assign n_9_net_ = v_o[2] & 1'b1;
  assign n_15_net_ = v_o[3] & 1'b1;
  assign n_21_net_ = v_o[4] & ready_i[4];
  assign n_27_net_ = v_o[0] & 1'b1;
  assign yumi_o[0] = N2 | W_gnt_p;
  assign N2 = N1 | P_gnt_p;
  assign N1 = N0 | S_gnt_p;
  assign N0 = E_gnt_p | N_gnt_p;
  assign yumi_o[1] = E_gnt_w | P_gnt_w;
  assign yumi_o[2] = W_gnt_e | P_gnt_e;
  assign yumi_o[3] = N4 | P_gnt_n;
  assign N4 = N3 | E_gnt_n;
  assign N3 = S_gnt_n | W_gnt_n;
  assign yumi_o[4] = N6 | P_gnt_s;
  assign N6 = N5 | E_gnt_s;
  assign N5 = N_gnt_s | W_gnt_s;

endmodule



module bsg_mesh_router_buffered_99_1_1_0_5_0d_0_101_00
(
  clk_i,
  reset_i,
  link_i,
  link_o,
  my_x_i,
  my_y_i
);

  input [504:0] link_i;
  output [504:0] link_o;
  input [0:0] my_x_i;
  input [0:0] my_y_i;
  input clk_i;
  input reset_i;
  wire [504:0] link_o;
  wire fifo_data_4__98_,fifo_data_4__97_,fifo_data_4__96_,fifo_data_4__95_,
  fifo_data_4__94_,fifo_data_4__93_,fifo_data_4__92_,fifo_data_4__91_,fifo_data_4__90_,
  fifo_data_4__89_,fifo_data_4__88_,fifo_data_4__87_,fifo_data_4__86_,fifo_data_4__85_,
  fifo_data_4__84_,fifo_data_4__83_,fifo_data_4__82_,fifo_data_4__81_,
  fifo_data_4__80_,fifo_data_4__79_,fifo_data_4__78_,fifo_data_4__77_,fifo_data_4__76_,
  fifo_data_4__75_,fifo_data_4__74_,fifo_data_4__73_,fifo_data_4__72_,fifo_data_4__71_,
  fifo_data_4__70_,fifo_data_4__69_,fifo_data_4__68_,fifo_data_4__67_,
  fifo_data_4__66_,fifo_data_4__65_,fifo_data_4__64_,fifo_data_4__63_,fifo_data_4__62_,
  fifo_data_4__61_,fifo_data_4__60_,fifo_data_4__59_,fifo_data_4__58_,fifo_data_4__57_,
  fifo_data_4__56_,fifo_data_4__55_,fifo_data_4__54_,fifo_data_4__53_,fifo_data_4__52_,
  fifo_data_4__51_,fifo_data_4__50_,fifo_data_4__49_,fifo_data_4__48_,
  fifo_data_4__47_,fifo_data_4__46_,fifo_data_4__45_,fifo_data_4__44_,fifo_data_4__43_,
  fifo_data_4__42_,fifo_data_4__41_,fifo_data_4__40_,fifo_data_4__39_,fifo_data_4__38_,
  fifo_data_4__37_,fifo_data_4__36_,fifo_data_4__35_,fifo_data_4__34_,
  fifo_data_4__33_,fifo_data_4__32_,fifo_data_4__31_,fifo_data_4__30_,fifo_data_4__29_,
  fifo_data_4__28_,fifo_data_4__27_,fifo_data_4__26_,fifo_data_4__25_,fifo_data_4__24_,
  fifo_data_4__23_,fifo_data_4__22_,fifo_data_4__21_,fifo_data_4__20_,fifo_data_4__19_,
  fifo_data_4__18_,fifo_data_4__17_,fifo_data_4__16_,fifo_data_4__15_,
  fifo_data_4__14_,fifo_data_4__13_,fifo_data_4__12_,fifo_data_4__11_,fifo_data_4__10_,
  fifo_data_4__9_,fifo_data_4__8_,fifo_data_4__7_,fifo_data_4__6_,fifo_data_4__5_,
  fifo_data_4__4_,fifo_data_4__3_,fifo_data_4__2_,fifo_data_4__1_,fifo_data_4__0_,
  fifo_data_1__98_,fifo_data_1__97_,fifo_data_1__96_,fifo_data_1__95_,fifo_data_1__94_,
  fifo_data_1__93_,fifo_data_1__92_,fifo_data_1__91_,fifo_data_1__90_,
  fifo_data_1__89_,fifo_data_1__88_,fifo_data_1__87_,fifo_data_1__86_,fifo_data_1__85_,
  fifo_data_1__84_,fifo_data_1__83_,fifo_data_1__82_,fifo_data_1__81_,fifo_data_1__80_,
  fifo_data_1__79_,fifo_data_1__78_,fifo_data_1__77_,fifo_data_1__76_,
  fifo_data_1__75_,fifo_data_1__74_,fifo_data_1__73_,fifo_data_1__72_,fifo_data_1__71_,
  fifo_data_1__70_,fifo_data_1__69_,fifo_data_1__68_,fifo_data_1__67_,fifo_data_1__66_,
  fifo_data_1__65_,fifo_data_1__64_,fifo_data_1__63_,fifo_data_1__62_,fifo_data_1__61_,
  fifo_data_1__60_,fifo_data_1__59_,fifo_data_1__58_,fifo_data_1__57_,
  fifo_data_1__56_,fifo_data_1__55_,fifo_data_1__54_,fifo_data_1__53_,fifo_data_1__52_,
  fifo_data_1__51_,fifo_data_1__50_,fifo_data_1__49_,fifo_data_1__48_,fifo_data_1__47_,
  fifo_data_1__46_,fifo_data_1__45_,fifo_data_1__44_,fifo_data_1__43_,
  fifo_data_1__42_,fifo_data_1__41_,fifo_data_1__40_,fifo_data_1__39_,fifo_data_1__38_,
  fifo_data_1__37_,fifo_data_1__36_,fifo_data_1__35_,fifo_data_1__34_,fifo_data_1__33_,
  fifo_data_1__32_,fifo_data_1__31_,fifo_data_1__30_,fifo_data_1__29_,fifo_data_1__28_,
  fifo_data_1__27_,fifo_data_1__26_,fifo_data_1__25_,fifo_data_1__24_,
  fifo_data_1__23_,fifo_data_1__22_,fifo_data_1__21_,fifo_data_1__20_,fifo_data_1__19_,
  fifo_data_1__18_,fifo_data_1__17_,fifo_data_1__16_,fifo_data_1__15_,fifo_data_1__14_,
  fifo_data_1__13_,fifo_data_1__12_,fifo_data_1__11_,fifo_data_1__10_,
  fifo_data_1__9_,fifo_data_1__8_,fifo_data_1__7_,fifo_data_1__6_,fifo_data_1__5_,
  fifo_data_1__4_,fifo_data_1__3_,fifo_data_1__2_,fifo_data_1__1_,fifo_data_1__0_,fifo_valid_1;
  wire [4:4] fifo_valid;
  wire [4:0] fifo_yumi;
  assign link_o[99] = 1'b0;
  assign link_o[301] = 1'b0;
  assign link_o[402] = 1'b0;

  bsg_two_fifo_width_p99
  rof_1__fi_twofer
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(link_o[200]),
    .data_i(link_i[199:101]),
    .v_i(link_i[201]),
    .v_o(fifo_valid_1),
    .data_o({ fifo_data_1__98_, fifo_data_1__97_, fifo_data_1__96_, fifo_data_1__95_, fifo_data_1__94_, fifo_data_1__93_, fifo_data_1__92_, fifo_data_1__91_, fifo_data_1__90_, fifo_data_1__89_, fifo_data_1__88_, fifo_data_1__87_, fifo_data_1__86_, fifo_data_1__85_, fifo_data_1__84_, fifo_data_1__83_, fifo_data_1__82_, fifo_data_1__81_, fifo_data_1__80_, fifo_data_1__79_, fifo_data_1__78_, fifo_data_1__77_, fifo_data_1__76_, fifo_data_1__75_, fifo_data_1__74_, fifo_data_1__73_, fifo_data_1__72_, fifo_data_1__71_, fifo_data_1__70_, fifo_data_1__69_, fifo_data_1__68_, fifo_data_1__67_, fifo_data_1__66_, fifo_data_1__65_, fifo_data_1__64_, fifo_data_1__63_, fifo_data_1__62_, fifo_data_1__61_, fifo_data_1__60_, fifo_data_1__59_, fifo_data_1__58_, fifo_data_1__57_, fifo_data_1__56_, fifo_data_1__55_, fifo_data_1__54_, fifo_data_1__53_, fifo_data_1__52_, fifo_data_1__51_, fifo_data_1__50_, fifo_data_1__49_, fifo_data_1__48_, fifo_data_1__47_, fifo_data_1__46_, fifo_data_1__45_, fifo_data_1__44_, fifo_data_1__43_, fifo_data_1__42_, fifo_data_1__41_, fifo_data_1__40_, fifo_data_1__39_, fifo_data_1__38_, fifo_data_1__37_, fifo_data_1__36_, fifo_data_1__35_, fifo_data_1__34_, fifo_data_1__33_, fifo_data_1__32_, fifo_data_1__31_, fifo_data_1__30_, fifo_data_1__29_, fifo_data_1__28_, fifo_data_1__27_, fifo_data_1__26_, fifo_data_1__25_, fifo_data_1__24_, fifo_data_1__23_, fifo_data_1__22_, fifo_data_1__21_, fifo_data_1__20_, fifo_data_1__19_, fifo_data_1__18_, fifo_data_1__17_, fifo_data_1__16_, fifo_data_1__15_, fifo_data_1__14_, fifo_data_1__13_, fifo_data_1__12_, fifo_data_1__11_, fifo_data_1__10_, fifo_data_1__9_, fifo_data_1__8_, fifo_data_1__7_, fifo_data_1__6_, fifo_data_1__5_, fifo_data_1__4_, fifo_data_1__3_, fifo_data_1__2_, fifo_data_1__1_, fifo_data_1__0_ }),
    .yumi_i(fifo_yumi[1])
  );


  bsg_two_fifo_width_p99
  rof_4__fi_twofer
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(link_o[503]),
    .data_i(link_i[502:404]),
    .v_i(link_i[504]),
    .v_o(fifo_valid[4]),
    .data_o({ fifo_data_4__98_, fifo_data_4__97_, fifo_data_4__96_, fifo_data_4__95_, fifo_data_4__94_, fifo_data_4__93_, fifo_data_4__92_, fifo_data_4__91_, fifo_data_4__90_, fifo_data_4__89_, fifo_data_4__88_, fifo_data_4__87_, fifo_data_4__86_, fifo_data_4__85_, fifo_data_4__84_, fifo_data_4__83_, fifo_data_4__82_, fifo_data_4__81_, fifo_data_4__80_, fifo_data_4__79_, fifo_data_4__78_, fifo_data_4__77_, fifo_data_4__76_, fifo_data_4__75_, fifo_data_4__74_, fifo_data_4__73_, fifo_data_4__72_, fifo_data_4__71_, fifo_data_4__70_, fifo_data_4__69_, fifo_data_4__68_, fifo_data_4__67_, fifo_data_4__66_, fifo_data_4__65_, fifo_data_4__64_, fifo_data_4__63_, fifo_data_4__62_, fifo_data_4__61_, fifo_data_4__60_, fifo_data_4__59_, fifo_data_4__58_, fifo_data_4__57_, fifo_data_4__56_, fifo_data_4__55_, fifo_data_4__54_, fifo_data_4__53_, fifo_data_4__52_, fifo_data_4__51_, fifo_data_4__50_, fifo_data_4__49_, fifo_data_4__48_, fifo_data_4__47_, fifo_data_4__46_, fifo_data_4__45_, fifo_data_4__44_, fifo_data_4__43_, fifo_data_4__42_, fifo_data_4__41_, fifo_data_4__40_, fifo_data_4__39_, fifo_data_4__38_, fifo_data_4__37_, fifo_data_4__36_, fifo_data_4__35_, fifo_data_4__34_, fifo_data_4__33_, fifo_data_4__32_, fifo_data_4__31_, fifo_data_4__30_, fifo_data_4__29_, fifo_data_4__28_, fifo_data_4__27_, fifo_data_4__26_, fifo_data_4__25_, fifo_data_4__24_, fifo_data_4__23_, fifo_data_4__22_, fifo_data_4__21_, fifo_data_4__20_, fifo_data_4__19_, fifo_data_4__18_, fifo_data_4__17_, fifo_data_4__16_, fifo_data_4__15_, fifo_data_4__14_, fifo_data_4__13_, fifo_data_4__12_, fifo_data_4__11_, fifo_data_4__10_, fifo_data_4__9_, fifo_data_4__8_, fifo_data_4__7_, fifo_data_4__6_, fifo_data_4__5_, fifo_data_4__4_, fifo_data_4__3_, fifo_data_4__2_, fifo_data_4__1_, fifo_data_4__0_ }),
    .yumi_i(fifo_yumi[4])
  );


  bsg_mesh_router_99_1_1_0_0d_0
  bmr
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ fifo_data_4__98_, fifo_data_4__97_, fifo_data_4__96_, fifo_data_4__95_, fifo_data_4__94_, fifo_data_4__93_, fifo_data_4__92_, fifo_data_4__91_, fifo_data_4__90_, fifo_data_4__89_, fifo_data_4__88_, fifo_data_4__87_, fifo_data_4__86_, fifo_data_4__85_, fifo_data_4__84_, fifo_data_4__83_, fifo_data_4__82_, fifo_data_4__81_, fifo_data_4__80_, fifo_data_4__79_, fifo_data_4__78_, fifo_data_4__77_, fifo_data_4__76_, fifo_data_4__75_, fifo_data_4__74_, fifo_data_4__73_, fifo_data_4__72_, fifo_data_4__71_, fifo_data_4__70_, fifo_data_4__69_, fifo_data_4__68_, fifo_data_4__67_, fifo_data_4__66_, fifo_data_4__65_, fifo_data_4__64_, fifo_data_4__63_, fifo_data_4__62_, fifo_data_4__61_, fifo_data_4__60_, fifo_data_4__59_, fifo_data_4__58_, fifo_data_4__57_, fifo_data_4__56_, fifo_data_4__55_, fifo_data_4__54_, fifo_data_4__53_, fifo_data_4__52_, fifo_data_4__51_, fifo_data_4__50_, fifo_data_4__49_, fifo_data_4__48_, fifo_data_4__47_, fifo_data_4__46_, fifo_data_4__45_, fifo_data_4__44_, fifo_data_4__43_, fifo_data_4__42_, fifo_data_4__41_, fifo_data_4__40_, fifo_data_4__39_, fifo_data_4__38_, fifo_data_4__37_, fifo_data_4__36_, fifo_data_4__35_, fifo_data_4__34_, fifo_data_4__33_, fifo_data_4__32_, fifo_data_4__31_, fifo_data_4__30_, fifo_data_4__29_, fifo_data_4__28_, fifo_data_4__27_, fifo_data_4__26_, fifo_data_4__25_, fifo_data_4__24_, fifo_data_4__23_, fifo_data_4__22_, fifo_data_4__21_, fifo_data_4__20_, fifo_data_4__19_, fifo_data_4__18_, fifo_data_4__17_, fifo_data_4__16_, fifo_data_4__15_, fifo_data_4__14_, fifo_data_4__13_, fifo_data_4__12_, fifo_data_4__11_, fifo_data_4__10_, fifo_data_4__9_, fifo_data_4__8_, fifo_data_4__7_, fifo_data_4__6_, fifo_data_4__5_, fifo_data_4__4_, fifo_data_4__3_, fifo_data_4__2_, fifo_data_4__1_, fifo_data_4__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_1__98_, fifo_data_1__97_, fifo_data_1__96_, fifo_data_1__95_, fifo_data_1__94_, fifo_data_1__93_, fifo_data_1__92_, fifo_data_1__91_, fifo_data_1__90_, fifo_data_1__89_, fifo_data_1__88_, fifo_data_1__87_, fifo_data_1__86_, fifo_data_1__85_, fifo_data_1__84_, fifo_data_1__83_, fifo_data_1__82_, fifo_data_1__81_, fifo_data_1__80_, fifo_data_1__79_, fifo_data_1__78_, fifo_data_1__77_, fifo_data_1__76_, fifo_data_1__75_, fifo_data_1__74_, fifo_data_1__73_, fifo_data_1__72_, fifo_data_1__71_, fifo_data_1__70_, fifo_data_1__69_, fifo_data_1__68_, fifo_data_1__67_, fifo_data_1__66_, fifo_data_1__65_, fifo_data_1__64_, fifo_data_1__63_, fifo_data_1__62_, fifo_data_1__61_, fifo_data_1__60_, fifo_data_1__59_, fifo_data_1__58_, fifo_data_1__57_, fifo_data_1__56_, fifo_data_1__55_, fifo_data_1__54_, fifo_data_1__53_, fifo_data_1__52_, fifo_data_1__51_, fifo_data_1__50_, fifo_data_1__49_, fifo_data_1__48_, fifo_data_1__47_, fifo_data_1__46_, fifo_data_1__45_, fifo_data_1__44_, fifo_data_1__43_, fifo_data_1__42_, fifo_data_1__41_, fifo_data_1__40_, fifo_data_1__39_, fifo_data_1__38_, fifo_data_1__37_, fifo_data_1__36_, fifo_data_1__35_, fifo_data_1__34_, fifo_data_1__33_, fifo_data_1__32_, fifo_data_1__31_, fifo_data_1__30_, fifo_data_1__29_, fifo_data_1__28_, fifo_data_1__27_, fifo_data_1__26_, fifo_data_1__25_, fifo_data_1__24_, fifo_data_1__23_, fifo_data_1__22_, fifo_data_1__21_, fifo_data_1__20_, fifo_data_1__19_, fifo_data_1__18_, fifo_data_1__17_, fifo_data_1__16_, fifo_data_1__15_, fifo_data_1__14_, fifo_data_1__13_, fifo_data_1__12_, fifo_data_1__11_, fifo_data_1__10_, fifo_data_1__9_, fifo_data_1__8_, fifo_data_1__7_, fifo_data_1__6_, fifo_data_1__5_, fifo_data_1__4_, fifo_data_1__3_, fifo_data_1__2_, fifo_data_1__1_, fifo_data_1__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .v_i({ fifo_valid[4:4], 1'b0, 1'b0, fifo_valid_1, 1'b0 }),
    .yumi_o(fifo_yumi),
    .ready_i({ link_i[503:503], link_i[402:402], link_i[301:301], link_i[200:200], link_i[99:99] }),
    .data_o({ link_o[502:404], link_o[401:303], link_o[300:202], link_o[199:101], link_o[98:0] }),
    .v_o({ link_o[504:504], link_o[403:403], link_o[302:302], link_o[201:201], link_o[100:100] }),
    .my_x_i(my_x_i[0]),
    .my_y_i(my_y_i[0])
  );


endmodule



module bp_me_network_channel_mesh_packet_width_p97_num_src_p2_num_dst_p1_debug_p0
(
  clk_i,
  reset_i,
  src_data_i,
  src_v_i,
  src_ready_o,
  dst_data_o,
  dst_v_o,
  dst_ready_i
);

  input [193:0] src_data_i;
  input [1:0] src_v_i;
  output [1:0] src_ready_o;
  output [96:0] dst_data_o;
  output [0:0] dst_v_o;
  input [0:0] dst_ready_i;
  input clk_i;
  input reset_i;
  wire [1:0] src_ready_o;
  wire [96:0] dst_data_o;
  wire [0:0] dst_v_o;
  wire link_i_stitch_0__2__v_,link_i_stitch_0__2__ready_then_rev_,
  link_i_stitch_0__2__data__98_,link_i_stitch_0__2__data__97_,link_i_stitch_0__2__data__96_,
  link_i_stitch_0__2__data__95_,link_i_stitch_0__2__data__94_,link_i_stitch_0__2__data__93_,
  link_i_stitch_0__2__data__92_,link_i_stitch_0__2__data__91_,
  link_i_stitch_0__2__data__90_,link_i_stitch_0__2__data__89_,link_i_stitch_0__2__data__88_,
  link_i_stitch_0__2__data__87_,link_i_stitch_0__2__data__86_,link_i_stitch_0__2__data__85_,
  link_i_stitch_0__2__data__84_,link_i_stitch_0__2__data__83_,
  link_i_stitch_0__2__data__82_,link_i_stitch_0__2__data__81_,link_i_stitch_0__2__data__80_,
  link_i_stitch_0__2__data__79_,link_i_stitch_0__2__data__78_,link_i_stitch_0__2__data__77_,
  link_i_stitch_0__2__data__76_,link_i_stitch_0__2__data__75_,
  link_i_stitch_0__2__data__74_,link_i_stitch_0__2__data__73_,link_i_stitch_0__2__data__72_,
  link_i_stitch_0__2__data__71_,link_i_stitch_0__2__data__70_,link_i_stitch_0__2__data__69_,
  link_i_stitch_0__2__data__68_,link_i_stitch_0__2__data__67_,
  link_i_stitch_0__2__data__66_,link_i_stitch_0__2__data__65_,link_i_stitch_0__2__data__64_,
  link_i_stitch_0__2__data__63_,link_i_stitch_0__2__data__62_,link_i_stitch_0__2__data__61_,
  link_i_stitch_0__2__data__60_,link_i_stitch_0__2__data__59_,
  link_i_stitch_0__2__data__58_,link_i_stitch_0__2__data__57_,link_i_stitch_0__2__data__56_,
  link_i_stitch_0__2__data__55_,link_i_stitch_0__2__data__54_,link_i_stitch_0__2__data__53_,
  link_i_stitch_0__2__data__52_,link_i_stitch_0__2__data__51_,
  link_i_stitch_0__2__data__50_,link_i_stitch_0__2__data__49_,link_i_stitch_0__2__data__48_,
  link_i_stitch_0__2__data__47_,link_i_stitch_0__2__data__46_,link_i_stitch_0__2__data__45_,
  link_i_stitch_0__2__data__44_,link_i_stitch_0__2__data__43_,
  link_i_stitch_0__2__data__42_,link_i_stitch_0__2__data__41_,link_i_stitch_0__2__data__40_,
  link_i_stitch_0__2__data__39_,link_i_stitch_0__2__data__38_,link_i_stitch_0__2__data__37_,
  link_i_stitch_0__2__data__36_,link_i_stitch_0__2__data__35_,
  link_i_stitch_0__2__data__34_,link_i_stitch_0__2__data__33_,link_i_stitch_0__2__data__32_,
  link_i_stitch_0__2__data__31_,link_i_stitch_0__2__data__30_,link_i_stitch_0__2__data__29_,
  link_i_stitch_0__2__data__28_,link_i_stitch_0__2__data__27_,
  link_i_stitch_0__2__data__26_,link_i_stitch_0__2__data__25_,link_i_stitch_0__2__data__24_,
  link_i_stitch_0__2__data__23_,link_i_stitch_0__2__data__22_,link_i_stitch_0__2__data__21_,
  link_i_stitch_0__2__data__20_,link_i_stitch_0__2__data__19_,
  link_i_stitch_0__2__data__18_,link_i_stitch_0__2__data__17_,link_i_stitch_0__2__data__16_,
  link_i_stitch_0__2__data__15_,link_i_stitch_0__2__data__14_,link_i_stitch_0__2__data__13_,
  link_i_stitch_0__2__data__12_,link_i_stitch_0__2__data__11_,
  link_i_stitch_0__2__data__10_,link_i_stitch_0__2__data__9_,link_i_stitch_0__2__data__8_,
  link_i_stitch_0__2__data__7_,link_i_stitch_0__2__data__6_,link_i_stitch_0__2__data__5_,
  link_i_stitch_0__2__data__4_,link_i_stitch_0__2__data__3_,
  link_i_stitch_0__2__data__2_,link_i_stitch_0__2__data__1_,link_i_stitch_0__2__data__0_,
  link_o_stitch_1__4__v_,link_o_stitch_1__4__data__98_,link_o_stitch_1__4__data__97_,
  link_o_stitch_1__4__data__96_,link_o_stitch_1__4__data__95_,link_o_stitch_1__4__data__94_,
  link_o_stitch_1__4__data__93_,link_o_stitch_1__4__data__92_,
  link_o_stitch_1__4__data__91_,link_o_stitch_1__4__data__90_,link_o_stitch_1__4__data__89_,
  link_o_stitch_1__4__data__88_,link_o_stitch_1__4__data__87_,link_o_stitch_1__4__data__86_,
  link_o_stitch_1__4__data__85_,link_o_stitch_1__4__data__84_,
  link_o_stitch_1__4__data__83_,link_o_stitch_1__4__data__82_,link_o_stitch_1__4__data__81_,
  link_o_stitch_1__4__data__80_,link_o_stitch_1__4__data__79_,link_o_stitch_1__4__data__78_,
  link_o_stitch_1__4__data__77_,link_o_stitch_1__4__data__76_,
  link_o_stitch_1__4__data__75_,link_o_stitch_1__4__data__74_,link_o_stitch_1__4__data__73_,
  link_o_stitch_1__4__data__72_,link_o_stitch_1__4__data__71_,link_o_stitch_1__4__data__70_,
  link_o_stitch_1__4__data__69_,link_o_stitch_1__4__data__68_,
  link_o_stitch_1__4__data__67_,link_o_stitch_1__4__data__66_,link_o_stitch_1__4__data__65_,
  link_o_stitch_1__4__data__64_,link_o_stitch_1__4__data__63_,link_o_stitch_1__4__data__62_,
  link_o_stitch_1__4__data__61_,link_o_stitch_1__4__data__60_,
  link_o_stitch_1__4__data__59_,link_o_stitch_1__4__data__58_,link_o_stitch_1__4__data__57_,
  link_o_stitch_1__4__data__56_,link_o_stitch_1__4__data__55_,link_o_stitch_1__4__data__54_,
  link_o_stitch_1__4__data__53_,link_o_stitch_1__4__data__52_,
  link_o_stitch_1__4__data__51_,link_o_stitch_1__4__data__50_,link_o_stitch_1__4__data__49_,
  link_o_stitch_1__4__data__48_,link_o_stitch_1__4__data__47_,link_o_stitch_1__4__data__46_,
  link_o_stitch_1__4__data__45_,link_o_stitch_1__4__data__44_,
  link_o_stitch_1__4__data__43_,link_o_stitch_1__4__data__42_,link_o_stitch_1__4__data__41_,
  link_o_stitch_1__4__data__40_,link_o_stitch_1__4__data__39_,link_o_stitch_1__4__data__38_,
  link_o_stitch_1__4__data__37_,link_o_stitch_1__4__data__36_,
  link_o_stitch_1__4__data__35_,link_o_stitch_1__4__data__34_,link_o_stitch_1__4__data__33_,
  link_o_stitch_1__4__data__32_,link_o_stitch_1__4__data__31_,link_o_stitch_1__4__data__30_,
  link_o_stitch_1__4__data__29_,link_o_stitch_1__4__data__28_,
  link_o_stitch_1__4__data__27_,link_o_stitch_1__4__data__26_,link_o_stitch_1__4__data__25_,
  link_o_stitch_1__4__data__24_,link_o_stitch_1__4__data__23_,link_o_stitch_1__4__data__22_,
  link_o_stitch_1__4__data__21_,link_o_stitch_1__4__data__20_,
  link_o_stitch_1__4__data__19_,link_o_stitch_1__4__data__18_,link_o_stitch_1__4__data__17_,
  link_o_stitch_1__4__data__16_,link_o_stitch_1__4__data__15_,link_o_stitch_1__4__data__14_,
  link_o_stitch_1__4__data__13_,link_o_stitch_1__4__data__12_,
  link_o_stitch_1__4__data__11_,link_o_stitch_1__4__data__10_,link_o_stitch_1__4__data__9_,
  link_o_stitch_1__4__data__8_,link_o_stitch_1__4__data__7_,link_o_stitch_1__4__data__6_,
  link_o_stitch_1__4__data__5_,link_o_stitch_1__4__data__4_,link_o_stitch_1__4__data__3_,
  link_o_stitch_1__4__data__2_,link_o_stitch_1__4__data__1_,
  link_o_stitch_1__4__data__0_,link_o_stitch_1__3__v_,link_o_stitch_1__3__ready_then_rev_,
  link_o_stitch_1__3__data__98_,link_o_stitch_1__3__data__97_,link_o_stitch_1__3__data__96_,
  link_o_stitch_1__3__data__95_,link_o_stitch_1__3__data__94_,
  link_o_stitch_1__3__data__93_,link_o_stitch_1__3__data__92_,link_o_stitch_1__3__data__91_,
  link_o_stitch_1__3__data__90_,link_o_stitch_1__3__data__89_,link_o_stitch_1__3__data__88_,
  link_o_stitch_1__3__data__87_,link_o_stitch_1__3__data__86_,
  link_o_stitch_1__3__data__85_,link_o_stitch_1__3__data__84_,link_o_stitch_1__3__data__83_,
  link_o_stitch_1__3__data__82_,link_o_stitch_1__3__data__81_,link_o_stitch_1__3__data__80_,
  link_o_stitch_1__3__data__79_,link_o_stitch_1__3__data__78_,
  link_o_stitch_1__3__data__77_,link_o_stitch_1__3__data__76_,link_o_stitch_1__3__data__75_,
  link_o_stitch_1__3__data__74_,link_o_stitch_1__3__data__73_,link_o_stitch_1__3__data__72_,
  link_o_stitch_1__3__data__71_,link_o_stitch_1__3__data__70_,
  link_o_stitch_1__3__data__69_,link_o_stitch_1__3__data__68_,link_o_stitch_1__3__data__67_,
  link_o_stitch_1__3__data__66_,link_o_stitch_1__3__data__65_,link_o_stitch_1__3__data__64_,
  link_o_stitch_1__3__data__63_,link_o_stitch_1__3__data__62_,
  link_o_stitch_1__3__data__61_,link_o_stitch_1__3__data__60_,link_o_stitch_1__3__data__59_,
  link_o_stitch_1__3__data__58_,link_o_stitch_1__3__data__57_,link_o_stitch_1__3__data__56_,
  link_o_stitch_1__3__data__55_,link_o_stitch_1__3__data__54_,
  link_o_stitch_1__3__data__53_,link_o_stitch_1__3__data__52_,link_o_stitch_1__3__data__51_,
  link_o_stitch_1__3__data__50_,link_o_stitch_1__3__data__49_,link_o_stitch_1__3__data__48_,
  link_o_stitch_1__3__data__47_,link_o_stitch_1__3__data__46_,
  link_o_stitch_1__3__data__45_,link_o_stitch_1__3__data__44_,link_o_stitch_1__3__data__43_,
  link_o_stitch_1__3__data__42_,link_o_stitch_1__3__data__41_,link_o_stitch_1__3__data__40_,
  link_o_stitch_1__3__data__39_,link_o_stitch_1__3__data__38_,
  link_o_stitch_1__3__data__37_,link_o_stitch_1__3__data__36_,link_o_stitch_1__3__data__35_,
  link_o_stitch_1__3__data__34_,link_o_stitch_1__3__data__33_,link_o_stitch_1__3__data__32_,
  link_o_stitch_1__3__data__31_,link_o_stitch_1__3__data__30_,
  link_o_stitch_1__3__data__29_,link_o_stitch_1__3__data__28_,link_o_stitch_1__3__data__27_,
  link_o_stitch_1__3__data__26_,link_o_stitch_1__3__data__25_,link_o_stitch_1__3__data__24_,
  link_o_stitch_1__3__data__23_,link_o_stitch_1__3__data__22_,
  link_o_stitch_1__3__data__21_,link_o_stitch_1__3__data__20_,link_o_stitch_1__3__data__19_,
  link_o_stitch_1__3__data__18_,link_o_stitch_1__3__data__17_,link_o_stitch_1__3__data__16_,
  link_o_stitch_1__3__data__15_,link_o_stitch_1__3__data__14_,
  link_o_stitch_1__3__data__13_,link_o_stitch_1__3__data__12_,link_o_stitch_1__3__data__11_,
  link_o_stitch_1__3__data__10_,link_o_stitch_1__3__data__9_,link_o_stitch_1__3__data__8_,
  link_o_stitch_1__3__data__7_,link_o_stitch_1__3__data__6_,link_o_stitch_1__3__data__5_,
  link_o_stitch_1__3__data__4_,link_o_stitch_1__3__data__3_,
  link_o_stitch_1__3__data__2_,link_o_stitch_1__3__data__1_,link_o_stitch_1__3__data__0_,
  link_o_stitch_1__2__v_,link_o_stitch_1__2__ready_then_rev_,link_o_stitch_1__2__data__98_,
  link_o_stitch_1__2__data__97_,link_o_stitch_1__2__data__96_,link_o_stitch_1__2__data__95_,
  link_o_stitch_1__2__data__94_,link_o_stitch_1__2__data__93_,
  link_o_stitch_1__2__data__92_,link_o_stitch_1__2__data__91_,link_o_stitch_1__2__data__90_,
  link_o_stitch_1__2__data__89_,link_o_stitch_1__2__data__88_,link_o_stitch_1__2__data__87_,
  link_o_stitch_1__2__data__86_,link_o_stitch_1__2__data__85_,
  link_o_stitch_1__2__data__84_,link_o_stitch_1__2__data__83_,link_o_stitch_1__2__data__82_,
  link_o_stitch_1__2__data__81_,link_o_stitch_1__2__data__80_,link_o_stitch_1__2__data__79_,
  link_o_stitch_1__2__data__78_,link_o_stitch_1__2__data__77_,
  link_o_stitch_1__2__data__76_,link_o_stitch_1__2__data__75_,link_o_stitch_1__2__data__74_,
  link_o_stitch_1__2__data__73_,link_o_stitch_1__2__data__72_,link_o_stitch_1__2__data__71_,
  link_o_stitch_1__2__data__70_,link_o_stitch_1__2__data__69_,
  link_o_stitch_1__2__data__68_,link_o_stitch_1__2__data__67_,link_o_stitch_1__2__data__66_,
  link_o_stitch_1__2__data__65_,link_o_stitch_1__2__data__64_,link_o_stitch_1__2__data__63_,
  link_o_stitch_1__2__data__62_,link_o_stitch_1__2__data__61_,
  link_o_stitch_1__2__data__60_,link_o_stitch_1__2__data__59_,link_o_stitch_1__2__data__58_,
  link_o_stitch_1__2__data__57_,link_o_stitch_1__2__data__56_,link_o_stitch_1__2__data__55_,
  link_o_stitch_1__2__data__54_,link_o_stitch_1__2__data__53_,
  link_o_stitch_1__2__data__52_,link_o_stitch_1__2__data__51_,link_o_stitch_1__2__data__50_,
  link_o_stitch_1__2__data__49_,link_o_stitch_1__2__data__48_,link_o_stitch_1__2__data__47_,
  link_o_stitch_1__2__data__46_,link_o_stitch_1__2__data__45_,
  link_o_stitch_1__2__data__44_,link_o_stitch_1__2__data__43_,link_o_stitch_1__2__data__42_,
  link_o_stitch_1__2__data__41_,link_o_stitch_1__2__data__40_,link_o_stitch_1__2__data__39_,
  link_o_stitch_1__2__data__38_,link_o_stitch_1__2__data__37_,
  link_o_stitch_1__2__data__36_,link_o_stitch_1__2__data__35_,link_o_stitch_1__2__data__34_,
  link_o_stitch_1__2__data__33_,link_o_stitch_1__2__data__32_,link_o_stitch_1__2__data__31_,
  link_o_stitch_1__2__data__30_,link_o_stitch_1__2__data__29_,
  link_o_stitch_1__2__data__28_,link_o_stitch_1__2__data__27_,link_o_stitch_1__2__data__26_,
  link_o_stitch_1__2__data__25_,link_o_stitch_1__2__data__24_,link_o_stitch_1__2__data__23_,
  link_o_stitch_1__2__data__22_,link_o_stitch_1__2__data__21_,
  link_o_stitch_1__2__data__20_,link_o_stitch_1__2__data__19_,link_o_stitch_1__2__data__18_,
  link_o_stitch_1__2__data__17_,link_o_stitch_1__2__data__16_,link_o_stitch_1__2__data__15_,
  link_o_stitch_1__2__data__14_,link_o_stitch_1__2__data__13_,
  link_o_stitch_1__2__data__12_,link_o_stitch_1__2__data__11_,link_o_stitch_1__2__data__10_,
  link_o_stitch_1__2__data__9_,link_o_stitch_1__2__data__8_,link_o_stitch_1__2__data__7_,
  link_o_stitch_1__2__data__6_,link_o_stitch_1__2__data__5_,
  link_o_stitch_1__2__data__4_,link_o_stitch_1__2__data__3_,link_o_stitch_1__2__data__2_,
  link_o_stitch_1__2__data__1_,link_o_stitch_1__2__data__0_,link_o_stitch_1__0__v_,
  link_o_stitch_1__0__ready_then_rev_,link_o_stitch_1__0__data__98_,link_o_stitch_1__0__data__97_,
  link_o_stitch_1__0__data__96_,link_o_stitch_1__0__data__95_,
  link_o_stitch_1__0__data__94_,link_o_stitch_1__0__data__93_,link_o_stitch_1__0__data__92_,
  link_o_stitch_1__0__data__91_,link_o_stitch_1__0__data__90_,link_o_stitch_1__0__data__89_,
  link_o_stitch_1__0__data__88_,link_o_stitch_1__0__data__87_,
  link_o_stitch_1__0__data__86_,link_o_stitch_1__0__data__85_,link_o_stitch_1__0__data__84_,
  link_o_stitch_1__0__data__83_,link_o_stitch_1__0__data__82_,link_o_stitch_1__0__data__81_,
  link_o_stitch_1__0__data__80_,link_o_stitch_1__0__data__79_,
  link_o_stitch_1__0__data__78_,link_o_stitch_1__0__data__77_,link_o_stitch_1__0__data__76_,
  link_o_stitch_1__0__data__75_,link_o_stitch_1__0__data__74_,link_o_stitch_1__0__data__73_,
  link_o_stitch_1__0__data__72_,link_o_stitch_1__0__data__71_,
  link_o_stitch_1__0__data__70_,link_o_stitch_1__0__data__69_,link_o_stitch_1__0__data__68_,
  link_o_stitch_1__0__data__67_,link_o_stitch_1__0__data__66_,link_o_stitch_1__0__data__65_,
  link_o_stitch_1__0__data__64_,link_o_stitch_1__0__data__63_,
  link_o_stitch_1__0__data__62_,link_o_stitch_1__0__data__61_,link_o_stitch_1__0__data__60_,
  link_o_stitch_1__0__data__59_,link_o_stitch_1__0__data__58_,link_o_stitch_1__0__data__57_,
  link_o_stitch_1__0__data__56_,link_o_stitch_1__0__data__55_,
  link_o_stitch_1__0__data__54_,link_o_stitch_1__0__data__53_,link_o_stitch_1__0__data__52_,
  link_o_stitch_1__0__data__51_,link_o_stitch_1__0__data__50_,link_o_stitch_1__0__data__49_,
  link_o_stitch_1__0__data__48_,link_o_stitch_1__0__data__47_,
  link_o_stitch_1__0__data__46_,link_o_stitch_1__0__data__45_,link_o_stitch_1__0__data__44_,
  link_o_stitch_1__0__data__43_,link_o_stitch_1__0__data__42_,link_o_stitch_1__0__data__41_,
  link_o_stitch_1__0__data__40_,link_o_stitch_1__0__data__39_,
  link_o_stitch_1__0__data__38_,link_o_stitch_1__0__data__37_,link_o_stitch_1__0__data__36_,
  link_o_stitch_1__0__data__35_,link_o_stitch_1__0__data__34_,link_o_stitch_1__0__data__33_,
  link_o_stitch_1__0__data__32_,link_o_stitch_1__0__data__31_,
  link_o_stitch_1__0__data__30_,link_o_stitch_1__0__data__29_,link_o_stitch_1__0__data__28_,
  link_o_stitch_1__0__data__27_,link_o_stitch_1__0__data__26_,link_o_stitch_1__0__data__25_,
  link_o_stitch_1__0__data__24_,link_o_stitch_1__0__data__23_,
  link_o_stitch_1__0__data__22_,link_o_stitch_1__0__data__21_,link_o_stitch_1__0__data__20_,
  link_o_stitch_1__0__data__19_,link_o_stitch_1__0__data__18_,link_o_stitch_1__0__data__17_,
  link_o_stitch_1__0__data__16_,link_o_stitch_1__0__data__15_,
  link_o_stitch_1__0__data__14_,link_o_stitch_1__0__data__13_,link_o_stitch_1__0__data__12_,
  link_o_stitch_1__0__data__11_,link_o_stitch_1__0__data__10_,link_o_stitch_1__0__data__9_,
  link_o_stitch_1__0__data__8_,link_o_stitch_1__0__data__7_,
  link_o_stitch_1__0__data__6_,link_o_stitch_1__0__data__5_,link_o_stitch_1__0__data__4_,
  link_o_stitch_1__0__data__3_,link_o_stitch_1__0__data__2_,link_o_stitch_1__0__data__1_,
  link_o_stitch_1__0__data__0_,link_o_stitch_0__4__v_,link_o_stitch_0__4__data__98_,
  link_o_stitch_0__4__data__97_,link_o_stitch_0__4__data__96_,
  link_o_stitch_0__4__data__95_,link_o_stitch_0__4__data__94_,link_o_stitch_0__4__data__93_,
  link_o_stitch_0__4__data__92_,link_o_stitch_0__4__data__91_,link_o_stitch_0__4__data__90_,
  link_o_stitch_0__4__data__89_,link_o_stitch_0__4__data__88_,
  link_o_stitch_0__4__data__87_,link_o_stitch_0__4__data__86_,link_o_stitch_0__4__data__85_,
  link_o_stitch_0__4__data__84_,link_o_stitch_0__4__data__83_,link_o_stitch_0__4__data__82_,
  link_o_stitch_0__4__data__81_,link_o_stitch_0__4__data__80_,
  link_o_stitch_0__4__data__79_,link_o_stitch_0__4__data__78_,link_o_stitch_0__4__data__77_,
  link_o_stitch_0__4__data__76_,link_o_stitch_0__4__data__75_,link_o_stitch_0__4__data__74_,
  link_o_stitch_0__4__data__73_,link_o_stitch_0__4__data__72_,
  link_o_stitch_0__4__data__71_,link_o_stitch_0__4__data__70_,link_o_stitch_0__4__data__69_,
  link_o_stitch_0__4__data__68_,link_o_stitch_0__4__data__67_,link_o_stitch_0__4__data__66_,
  link_o_stitch_0__4__data__65_,link_o_stitch_0__4__data__64_,
  link_o_stitch_0__4__data__63_,link_o_stitch_0__4__data__62_,link_o_stitch_0__4__data__61_,
  link_o_stitch_0__4__data__60_,link_o_stitch_0__4__data__59_,link_o_stitch_0__4__data__58_,
  link_o_stitch_0__4__data__57_,link_o_stitch_0__4__data__56_,
  link_o_stitch_0__4__data__55_,link_o_stitch_0__4__data__54_,link_o_stitch_0__4__data__53_,
  link_o_stitch_0__4__data__52_,link_o_stitch_0__4__data__51_,link_o_stitch_0__4__data__50_,
  link_o_stitch_0__4__data__49_,link_o_stitch_0__4__data__48_,
  link_o_stitch_0__4__data__47_,link_o_stitch_0__4__data__46_,link_o_stitch_0__4__data__45_,
  link_o_stitch_0__4__data__44_,link_o_stitch_0__4__data__43_,link_o_stitch_0__4__data__42_,
  link_o_stitch_0__4__data__41_,link_o_stitch_0__4__data__40_,
  link_o_stitch_0__4__data__39_,link_o_stitch_0__4__data__38_,link_o_stitch_0__4__data__37_,
  link_o_stitch_0__4__data__36_,link_o_stitch_0__4__data__35_,link_o_stitch_0__4__data__34_,
  link_o_stitch_0__4__data__33_,link_o_stitch_0__4__data__32_,
  link_o_stitch_0__4__data__31_,link_o_stitch_0__4__data__30_,link_o_stitch_0__4__data__29_,
  link_o_stitch_0__4__data__28_,link_o_stitch_0__4__data__27_,link_o_stitch_0__4__data__26_,
  link_o_stitch_0__4__data__25_,link_o_stitch_0__4__data__24_,
  link_o_stitch_0__4__data__23_,link_o_stitch_0__4__data__22_,link_o_stitch_0__4__data__21_,
  link_o_stitch_0__4__data__20_,link_o_stitch_0__4__data__19_,link_o_stitch_0__4__data__18_,
  link_o_stitch_0__4__data__17_,link_o_stitch_0__4__data__16_,
  link_o_stitch_0__4__data__15_,link_o_stitch_0__4__data__14_,link_o_stitch_0__4__data__13_,
  link_o_stitch_0__4__data__12_,link_o_stitch_0__4__data__11_,link_o_stitch_0__4__data__10_,
  link_o_stitch_0__4__data__9_,link_o_stitch_0__4__data__8_,link_o_stitch_0__4__data__7_,
  link_o_stitch_0__4__data__6_,link_o_stitch_0__4__data__5_,
  link_o_stitch_0__4__data__4_,link_o_stitch_0__4__data__3_,link_o_stitch_0__4__data__2_,
  link_o_stitch_0__4__data__1_,link_o_stitch_0__4__data__0_,link_o_stitch_0__3__v_,
  link_o_stitch_0__3__ready_then_rev_,link_o_stitch_0__3__data__98_,
  link_o_stitch_0__3__data__97_,link_o_stitch_0__3__data__96_,link_o_stitch_0__3__data__95_,
  link_o_stitch_0__3__data__94_,link_o_stitch_0__3__data__93_,link_o_stitch_0__3__data__92_,
  link_o_stitch_0__3__data__91_,link_o_stitch_0__3__data__90_,
  link_o_stitch_0__3__data__89_,link_o_stitch_0__3__data__88_,link_o_stitch_0__3__data__87_,
  link_o_stitch_0__3__data__86_,link_o_stitch_0__3__data__85_,link_o_stitch_0__3__data__84_,
  link_o_stitch_0__3__data__83_,link_o_stitch_0__3__data__82_,
  link_o_stitch_0__3__data__81_,link_o_stitch_0__3__data__80_,link_o_stitch_0__3__data__79_,
  link_o_stitch_0__3__data__78_,link_o_stitch_0__3__data__77_,link_o_stitch_0__3__data__76_,
  link_o_stitch_0__3__data__75_,link_o_stitch_0__3__data__74_,
  link_o_stitch_0__3__data__73_,link_o_stitch_0__3__data__72_,link_o_stitch_0__3__data__71_,
  link_o_stitch_0__3__data__70_,link_o_stitch_0__3__data__69_,link_o_stitch_0__3__data__68_,
  link_o_stitch_0__3__data__67_,link_o_stitch_0__3__data__66_,
  link_o_stitch_0__3__data__65_,link_o_stitch_0__3__data__64_,link_o_stitch_0__3__data__63_,
  link_o_stitch_0__3__data__62_,link_o_stitch_0__3__data__61_,link_o_stitch_0__3__data__60_,
  link_o_stitch_0__3__data__59_,link_o_stitch_0__3__data__58_,
  link_o_stitch_0__3__data__57_,link_o_stitch_0__3__data__56_,link_o_stitch_0__3__data__55_,
  link_o_stitch_0__3__data__54_,link_o_stitch_0__3__data__53_,link_o_stitch_0__3__data__52_,
  link_o_stitch_0__3__data__51_,link_o_stitch_0__3__data__50_,
  link_o_stitch_0__3__data__49_,link_o_stitch_0__3__data__48_,link_o_stitch_0__3__data__47_,
  link_o_stitch_0__3__data__46_,link_o_stitch_0__3__data__45_,link_o_stitch_0__3__data__44_,
  link_o_stitch_0__3__data__43_,link_o_stitch_0__3__data__42_,
  link_o_stitch_0__3__data__41_,link_o_stitch_0__3__data__40_,link_o_stitch_0__3__data__39_,
  link_o_stitch_0__3__data__38_,link_o_stitch_0__3__data__37_,link_o_stitch_0__3__data__36_,
  link_o_stitch_0__3__data__35_,link_o_stitch_0__3__data__34_,
  link_o_stitch_0__3__data__33_,link_o_stitch_0__3__data__32_,link_o_stitch_0__3__data__31_,
  link_o_stitch_0__3__data__30_,link_o_stitch_0__3__data__29_,link_o_stitch_0__3__data__28_,
  link_o_stitch_0__3__data__27_,link_o_stitch_0__3__data__26_,
  link_o_stitch_0__3__data__25_,link_o_stitch_0__3__data__24_,link_o_stitch_0__3__data__23_,
  link_o_stitch_0__3__data__22_,link_o_stitch_0__3__data__21_,link_o_stitch_0__3__data__20_,
  link_o_stitch_0__3__data__19_,link_o_stitch_0__3__data__18_,
  link_o_stitch_0__3__data__17_,link_o_stitch_0__3__data__16_,link_o_stitch_0__3__data__15_,
  link_o_stitch_0__3__data__14_,link_o_stitch_0__3__data__13_,link_o_stitch_0__3__data__12_,
  link_o_stitch_0__3__data__11_,link_o_stitch_0__3__data__10_,link_o_stitch_0__3__data__9_,
  link_o_stitch_0__3__data__8_,link_o_stitch_0__3__data__7_,
  link_o_stitch_0__3__data__6_,link_o_stitch_0__3__data__5_,link_o_stitch_0__3__data__4_,
  link_o_stitch_0__3__data__3_,link_o_stitch_0__3__data__2_,link_o_stitch_0__3__data__1_,
  link_o_stitch_0__3__data__0_,link_o_stitch_0__2__v_,link_o_stitch_0__2__ready_then_rev_,
  link_o_stitch_0__2__data__98_,link_o_stitch_0__2__data__97_,
  link_o_stitch_0__2__data__96_,link_o_stitch_0__2__data__95_,link_o_stitch_0__2__data__94_,
  link_o_stitch_0__2__data__93_,link_o_stitch_0__2__data__92_,link_o_stitch_0__2__data__91_,
  link_o_stitch_0__2__data__90_,link_o_stitch_0__2__data__89_,
  link_o_stitch_0__2__data__88_,link_o_stitch_0__2__data__87_,link_o_stitch_0__2__data__86_,
  link_o_stitch_0__2__data__85_,link_o_stitch_0__2__data__84_,link_o_stitch_0__2__data__83_,
  link_o_stitch_0__2__data__82_,link_o_stitch_0__2__data__81_,
  link_o_stitch_0__2__data__80_,link_o_stitch_0__2__data__79_,link_o_stitch_0__2__data__78_,
  link_o_stitch_0__2__data__77_,link_o_stitch_0__2__data__76_,link_o_stitch_0__2__data__75_,
  link_o_stitch_0__2__data__74_,link_o_stitch_0__2__data__73_,
  link_o_stitch_0__2__data__72_,link_o_stitch_0__2__data__71_,link_o_stitch_0__2__data__70_,
  link_o_stitch_0__2__data__69_,link_o_stitch_0__2__data__68_,link_o_stitch_0__2__data__67_,
  link_o_stitch_0__2__data__66_,link_o_stitch_0__2__data__65_,
  link_o_stitch_0__2__data__64_,link_o_stitch_0__2__data__63_,link_o_stitch_0__2__data__62_,
  link_o_stitch_0__2__data__61_,link_o_stitch_0__2__data__60_,link_o_stitch_0__2__data__59_,
  link_o_stitch_0__2__data__58_,link_o_stitch_0__2__data__57_,
  link_o_stitch_0__2__data__56_,link_o_stitch_0__2__data__55_,link_o_stitch_0__2__data__54_,
  link_o_stitch_0__2__data__53_,link_o_stitch_0__2__data__52_,link_o_stitch_0__2__data__51_,
  link_o_stitch_0__2__data__50_,link_o_stitch_0__2__data__49_,
  link_o_stitch_0__2__data__48_,link_o_stitch_0__2__data__47_,link_o_stitch_0__2__data__46_,
  link_o_stitch_0__2__data__45_,link_o_stitch_0__2__data__44_,link_o_stitch_0__2__data__43_,
  link_o_stitch_0__2__data__42_,link_o_stitch_0__2__data__41_,
  link_o_stitch_0__2__data__40_,link_o_stitch_0__2__data__39_,link_o_stitch_0__2__data__38_,
  link_o_stitch_0__2__data__37_,link_o_stitch_0__2__data__36_,link_o_stitch_0__2__data__35_,
  link_o_stitch_0__2__data__34_,link_o_stitch_0__2__data__33_,
  link_o_stitch_0__2__data__32_,link_o_stitch_0__2__data__31_,link_o_stitch_0__2__data__30_,
  link_o_stitch_0__2__data__29_,link_o_stitch_0__2__data__28_,link_o_stitch_0__2__data__27_,
  link_o_stitch_0__2__data__26_,link_o_stitch_0__2__data__25_,
  link_o_stitch_0__2__data__24_,link_o_stitch_0__2__data__23_,link_o_stitch_0__2__data__22_,
  link_o_stitch_0__2__data__21_,link_o_stitch_0__2__data__20_,link_o_stitch_0__2__data__19_,
  link_o_stitch_0__2__data__18_,link_o_stitch_0__2__data__17_,
  link_o_stitch_0__2__data__16_,link_o_stitch_0__2__data__15_,link_o_stitch_0__2__data__14_,
  link_o_stitch_0__2__data__13_,link_o_stitch_0__2__data__12_,link_o_stitch_0__2__data__11_,
  link_o_stitch_0__2__data__10_,link_o_stitch_0__2__data__9_,
  link_o_stitch_0__2__data__8_,link_o_stitch_0__2__data__7_,link_o_stitch_0__2__data__6_,
  link_o_stitch_0__2__data__5_,link_o_stitch_0__2__data__4_,link_o_stitch_0__2__data__3_,
  link_o_stitch_0__2__data__2_,link_o_stitch_0__2__data__1_,link_o_stitch_0__2__data__0_,
  link_o_stitch_0__1__v_,link_o_stitch_0__1__ready_then_rev_,
  link_o_stitch_0__1__data__98_,link_o_stitch_0__1__data__97_,link_o_stitch_0__1__data__96_,
  link_o_stitch_0__1__data__95_,link_o_stitch_0__1__data__94_,link_o_stitch_0__1__data__93_,
  link_o_stitch_0__1__data__92_,link_o_stitch_0__1__data__91_,
  link_o_stitch_0__1__data__90_,link_o_stitch_0__1__data__89_,link_o_stitch_0__1__data__88_,
  link_o_stitch_0__1__data__87_,link_o_stitch_0__1__data__86_,link_o_stitch_0__1__data__85_,
  link_o_stitch_0__1__data__84_,link_o_stitch_0__1__data__83_,
  link_o_stitch_0__1__data__82_,link_o_stitch_0__1__data__81_,link_o_stitch_0__1__data__80_,
  link_o_stitch_0__1__data__79_,link_o_stitch_0__1__data__78_,link_o_stitch_0__1__data__77_,
  link_o_stitch_0__1__data__76_,link_o_stitch_0__1__data__75_,
  link_o_stitch_0__1__data__74_,link_o_stitch_0__1__data__73_,link_o_stitch_0__1__data__72_,
  link_o_stitch_0__1__data__71_,link_o_stitch_0__1__data__70_,link_o_stitch_0__1__data__69_,
  link_o_stitch_0__1__data__68_,link_o_stitch_0__1__data__67_,
  link_o_stitch_0__1__data__66_,link_o_stitch_0__1__data__65_,link_o_stitch_0__1__data__64_,
  link_o_stitch_0__1__data__63_,link_o_stitch_0__1__data__62_,link_o_stitch_0__1__data__61_,
  link_o_stitch_0__1__data__60_,link_o_stitch_0__1__data__59_,
  link_o_stitch_0__1__data__58_,link_o_stitch_0__1__data__57_,link_o_stitch_0__1__data__56_,
  link_o_stitch_0__1__data__55_,link_o_stitch_0__1__data__54_,link_o_stitch_0__1__data__53_,
  link_o_stitch_0__1__data__52_,link_o_stitch_0__1__data__51_,
  link_o_stitch_0__1__data__50_,link_o_stitch_0__1__data__49_,link_o_stitch_0__1__data__48_,
  link_o_stitch_0__1__data__47_,link_o_stitch_0__1__data__46_,link_o_stitch_0__1__data__45_,
  link_o_stitch_0__1__data__44_,link_o_stitch_0__1__data__43_,
  link_o_stitch_0__1__data__42_,link_o_stitch_0__1__data__41_,link_o_stitch_0__1__data__40_,
  link_o_stitch_0__1__data__39_,link_o_stitch_0__1__data__38_,link_o_stitch_0__1__data__37_,
  link_o_stitch_0__1__data__36_,link_o_stitch_0__1__data__35_,
  link_o_stitch_0__1__data__34_,link_o_stitch_0__1__data__33_,link_o_stitch_0__1__data__32_,
  link_o_stitch_0__1__data__31_,link_o_stitch_0__1__data__30_,link_o_stitch_0__1__data__29_,
  link_o_stitch_0__1__data__28_,link_o_stitch_0__1__data__27_,
  link_o_stitch_0__1__data__26_,link_o_stitch_0__1__data__25_,link_o_stitch_0__1__data__24_,
  link_o_stitch_0__1__data__23_,link_o_stitch_0__1__data__22_,link_o_stitch_0__1__data__21_,
  link_o_stitch_0__1__data__20_,link_o_stitch_0__1__data__19_,
  link_o_stitch_0__1__data__18_,link_o_stitch_0__1__data__17_,link_o_stitch_0__1__data__16_,
  link_o_stitch_0__1__data__15_,link_o_stitch_0__1__data__14_,link_o_stitch_0__1__data__13_,
  link_o_stitch_0__1__data__12_,link_o_stitch_0__1__data__11_,
  link_o_stitch_0__1__data__10_,link_o_stitch_0__1__data__9_,link_o_stitch_0__1__data__8_,
  link_o_stitch_0__1__data__7_,link_o_stitch_0__1__data__6_,link_o_stitch_0__1__data__5_,
  link_o_stitch_0__1__data__4_,link_o_stitch_0__1__data__3_,
  link_o_stitch_0__1__data__2_,link_o_stitch_0__1__data__1_,link_o_stitch_0__1__data__0_,
  link_o_stitch_0__0__ready_then_rev_,link_o_stitch_0__0__data__1_,link_o_stitch_0__0__data__0_;

  bsg_mesh_router_buffered_99_1_1_0_5_0a_0_101_00
  rof_0__fi2_efi3_coherence_network_channel_node
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .link_i({ src_v_i[0:0], 1'b0, src_data_i[96:0], 1'b1, src_data_i[96:96], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, link_i_stitch_0__2__v_, link_i_stitch_0__2__ready_then_rev_, link_i_stitch_0__2__data__98_, link_i_stitch_0__2__data__97_, link_i_stitch_0__2__data__96_, link_i_stitch_0__2__data__95_, link_i_stitch_0__2__data__94_, link_i_stitch_0__2__data__93_, link_i_stitch_0__2__data__92_, link_i_stitch_0__2__data__91_, link_i_stitch_0__2__data__90_, link_i_stitch_0__2__data__89_, link_i_stitch_0__2__data__88_, link_i_stitch_0__2__data__87_, link_i_stitch_0__2__data__86_, link_i_stitch_0__2__data__85_, link_i_stitch_0__2__data__84_, link_i_stitch_0__2__data__83_, link_i_stitch_0__2__data__82_, link_i_stitch_0__2__data__81_, link_i_stitch_0__2__data__80_, link_i_stitch_0__2__data__79_, link_i_stitch_0__2__data__78_, link_i_stitch_0__2__data__77_, link_i_stitch_0__2__data__76_, link_i_stitch_0__2__data__75_, link_i_stitch_0__2__data__74_, link_i_stitch_0__2__data__73_, link_i_stitch_0__2__data__72_, link_i_stitch_0__2__data__71_, link_i_stitch_0__2__data__70_, link_i_stitch_0__2__data__69_, link_i_stitch_0__2__data__68_, link_i_stitch_0__2__data__67_, link_i_stitch_0__2__data__66_, link_i_stitch_0__2__data__65_, link_i_stitch_0__2__data__64_, link_i_stitch_0__2__data__63_, link_i_stitch_0__2__data__62_, link_i_stitch_0__2__data__61_, link_i_stitch_0__2__data__60_, link_i_stitch_0__2__data__59_, link_i_stitch_0__2__data__58_, link_i_stitch_0__2__data__57_, link_i_stitch_0__2__data__56_, link_i_stitch_0__2__data__55_, link_i_stitch_0__2__data__54_, link_i_stitch_0__2__data__53_, link_i_stitch_0__2__data__52_, link_i_stitch_0__2__data__51_, link_i_stitch_0__2__data__50_, link_i_stitch_0__2__data__49_, link_i_stitch_0__2__data__48_, link_i_stitch_0__2__data__47_, link_i_stitch_0__2__data__46_, link_i_stitch_0__2__data__45_, link_i_stitch_0__2__data__44_, link_i_stitch_0__2__data__43_, link_i_stitch_0__2__data__42_, link_i_stitch_0__2__data__41_, link_i_stitch_0__2__data__40_, link_i_stitch_0__2__data__39_, link_i_stitch_0__2__data__38_, link_i_stitch_0__2__data__37_, link_i_stitch_0__2__data__36_, link_i_stitch_0__2__data__35_, link_i_stitch_0__2__data__34_, link_i_stitch_0__2__data__33_, link_i_stitch_0__2__data__32_, link_i_stitch_0__2__data__31_, link_i_stitch_0__2__data__30_, link_i_stitch_0__2__data__29_, link_i_stitch_0__2__data__28_, link_i_stitch_0__2__data__27_, link_i_stitch_0__2__data__26_, link_i_stitch_0__2__data__25_, link_i_stitch_0__2__data__24_, link_i_stitch_0__2__data__23_, link_i_stitch_0__2__data__22_, link_i_stitch_0__2__data__21_, link_i_stitch_0__2__data__20_, link_i_stitch_0__2__data__19_, link_i_stitch_0__2__data__18_, link_i_stitch_0__2__data__17_, link_i_stitch_0__2__data__16_, link_i_stitch_0__2__data__15_, link_i_stitch_0__2__data__14_, link_i_stitch_0__2__data__13_, link_i_stitch_0__2__data__12_, link_i_stitch_0__2__data__11_, link_i_stitch_0__2__data__10_, link_i_stitch_0__2__data__9_, link_i_stitch_0__2__data__8_, link_i_stitch_0__2__data__7_, link_i_stitch_0__2__data__6_, link_i_stitch_0__2__data__5_, link_i_stitch_0__2__data__4_, link_i_stitch_0__2__data__3_, link_i_stitch_0__2__data__2_, link_i_stitch_0__2__data__1_, link_i_stitch_0__2__data__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, dst_ready_i[0:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .link_o({ link_o_stitch_0__4__v_, src_ready_o[0:0], link_o_stitch_0__4__data__98_, link_o_stitch_0__4__data__97_, link_o_stitch_0__4__data__96_, link_o_stitch_0__4__data__95_, link_o_stitch_0__4__data__94_, link_o_stitch_0__4__data__93_, link_o_stitch_0__4__data__92_, link_o_stitch_0__4__data__91_, link_o_stitch_0__4__data__90_, link_o_stitch_0__4__data__89_, link_o_stitch_0__4__data__88_, link_o_stitch_0__4__data__87_, link_o_stitch_0__4__data__86_, link_o_stitch_0__4__data__85_, link_o_stitch_0__4__data__84_, link_o_stitch_0__4__data__83_, link_o_stitch_0__4__data__82_, link_o_stitch_0__4__data__81_, link_o_stitch_0__4__data__80_, link_o_stitch_0__4__data__79_, link_o_stitch_0__4__data__78_, link_o_stitch_0__4__data__77_, link_o_stitch_0__4__data__76_, link_o_stitch_0__4__data__75_, link_o_stitch_0__4__data__74_, link_o_stitch_0__4__data__73_, link_o_stitch_0__4__data__72_, link_o_stitch_0__4__data__71_, link_o_stitch_0__4__data__70_, link_o_stitch_0__4__data__69_, link_o_stitch_0__4__data__68_, link_o_stitch_0__4__data__67_, link_o_stitch_0__4__data__66_, link_o_stitch_0__4__data__65_, link_o_stitch_0__4__data__64_, link_o_stitch_0__4__data__63_, link_o_stitch_0__4__data__62_, link_o_stitch_0__4__data__61_, link_o_stitch_0__4__data__60_, link_o_stitch_0__4__data__59_, link_o_stitch_0__4__data__58_, link_o_stitch_0__4__data__57_, link_o_stitch_0__4__data__56_, link_o_stitch_0__4__data__55_, link_o_stitch_0__4__data__54_, link_o_stitch_0__4__data__53_, link_o_stitch_0__4__data__52_, link_o_stitch_0__4__data__51_, link_o_stitch_0__4__data__50_, link_o_stitch_0__4__data__49_, link_o_stitch_0__4__data__48_, link_o_stitch_0__4__data__47_, link_o_stitch_0__4__data__46_, link_o_stitch_0__4__data__45_, link_o_stitch_0__4__data__44_, link_o_stitch_0__4__data__43_, link_o_stitch_0__4__data__42_, link_o_stitch_0__4__data__41_, link_o_stitch_0__4__data__40_, link_o_stitch_0__4__data__39_, link_o_stitch_0__4__data__38_, link_o_stitch_0__4__data__37_, link_o_stitch_0__4__data__36_, link_o_stitch_0__4__data__35_, link_o_stitch_0__4__data__34_, link_o_stitch_0__4__data__33_, link_o_stitch_0__4__data__32_, link_o_stitch_0__4__data__31_, link_o_stitch_0__4__data__30_, link_o_stitch_0__4__data__29_, link_o_stitch_0__4__data__28_, link_o_stitch_0__4__data__27_, link_o_stitch_0__4__data__26_, link_o_stitch_0__4__data__25_, link_o_stitch_0__4__data__24_, link_o_stitch_0__4__data__23_, link_o_stitch_0__4__data__22_, link_o_stitch_0__4__data__21_, link_o_stitch_0__4__data__20_, link_o_stitch_0__4__data__19_, link_o_stitch_0__4__data__18_, link_o_stitch_0__4__data__17_, link_o_stitch_0__4__data__16_, link_o_stitch_0__4__data__15_, link_o_stitch_0__4__data__14_, link_o_stitch_0__4__data__13_, link_o_stitch_0__4__data__12_, link_o_stitch_0__4__data__11_, link_o_stitch_0__4__data__10_, link_o_stitch_0__4__data__9_, link_o_stitch_0__4__data__8_, link_o_stitch_0__4__data__7_, link_o_stitch_0__4__data__6_, link_o_stitch_0__4__data__5_, link_o_stitch_0__4__data__4_, link_o_stitch_0__4__data__3_, link_o_stitch_0__4__data__2_, link_o_stitch_0__4__data__1_, link_o_stitch_0__4__data__0_, link_o_stitch_0__3__v_, link_o_stitch_0__3__ready_then_rev_, link_o_stitch_0__3__data__98_, link_o_stitch_0__3__data__97_, link_o_stitch_0__3__data__96_, link_o_stitch_0__3__data__95_, link_o_stitch_0__3__data__94_, link_o_stitch_0__3__data__93_, link_o_stitch_0__3__data__92_, link_o_stitch_0__3__data__91_, link_o_stitch_0__3__data__90_, link_o_stitch_0__3__data__89_, link_o_stitch_0__3__data__88_, link_o_stitch_0__3__data__87_, link_o_stitch_0__3__data__86_, link_o_stitch_0__3__data__85_, link_o_stitch_0__3__data__84_, link_o_stitch_0__3__data__83_, link_o_stitch_0__3__data__82_, link_o_stitch_0__3__data__81_, link_o_stitch_0__3__data__80_, link_o_stitch_0__3__data__79_, link_o_stitch_0__3__data__78_, link_o_stitch_0__3__data__77_, link_o_stitch_0__3__data__76_, link_o_stitch_0__3__data__75_, link_o_stitch_0__3__data__74_, link_o_stitch_0__3__data__73_, link_o_stitch_0__3__data__72_, link_o_stitch_0__3__data__71_, link_o_stitch_0__3__data__70_, link_o_stitch_0__3__data__69_, link_o_stitch_0__3__data__68_, link_o_stitch_0__3__data__67_, link_o_stitch_0__3__data__66_, link_o_stitch_0__3__data__65_, link_o_stitch_0__3__data__64_, link_o_stitch_0__3__data__63_, link_o_stitch_0__3__data__62_, link_o_stitch_0__3__data__61_, link_o_stitch_0__3__data__60_, link_o_stitch_0__3__data__59_, link_o_stitch_0__3__data__58_, link_o_stitch_0__3__data__57_, link_o_stitch_0__3__data__56_, link_o_stitch_0__3__data__55_, link_o_stitch_0__3__data__54_, link_o_stitch_0__3__data__53_, link_o_stitch_0__3__data__52_, link_o_stitch_0__3__data__51_, link_o_stitch_0__3__data__50_, link_o_stitch_0__3__data__49_, link_o_stitch_0__3__data__48_, link_o_stitch_0__3__data__47_, link_o_stitch_0__3__data__46_, link_o_stitch_0__3__data__45_, link_o_stitch_0__3__data__44_, link_o_stitch_0__3__data__43_, link_o_stitch_0__3__data__42_, link_o_stitch_0__3__data__41_, link_o_stitch_0__3__data__40_, link_o_stitch_0__3__data__39_, link_o_stitch_0__3__data__38_, link_o_stitch_0__3__data__37_, link_o_stitch_0__3__data__36_, link_o_stitch_0__3__data__35_, link_o_stitch_0__3__data__34_, link_o_stitch_0__3__data__33_, link_o_stitch_0__3__data__32_, link_o_stitch_0__3__data__31_, link_o_stitch_0__3__data__30_, link_o_stitch_0__3__data__29_, link_o_stitch_0__3__data__28_, link_o_stitch_0__3__data__27_, link_o_stitch_0__3__data__26_, link_o_stitch_0__3__data__25_, link_o_stitch_0__3__data__24_, link_o_stitch_0__3__data__23_, link_o_stitch_0__3__data__22_, link_o_stitch_0__3__data__21_, link_o_stitch_0__3__data__20_, link_o_stitch_0__3__data__19_, link_o_stitch_0__3__data__18_, link_o_stitch_0__3__data__17_, link_o_stitch_0__3__data__16_, link_o_stitch_0__3__data__15_, link_o_stitch_0__3__data__14_, link_o_stitch_0__3__data__13_, link_o_stitch_0__3__data__12_, link_o_stitch_0__3__data__11_, link_o_stitch_0__3__data__10_, link_o_stitch_0__3__data__9_, link_o_stitch_0__3__data__8_, link_o_stitch_0__3__data__7_, link_o_stitch_0__3__data__6_, link_o_stitch_0__3__data__5_, link_o_stitch_0__3__data__4_, link_o_stitch_0__3__data__3_, link_o_stitch_0__3__data__2_, link_o_stitch_0__3__data__1_, link_o_stitch_0__3__data__0_, link_o_stitch_0__2__v_, link_o_stitch_0__2__ready_then_rev_, link_o_stitch_0__2__data__98_, link_o_stitch_0__2__data__97_, link_o_stitch_0__2__data__96_, link_o_stitch_0__2__data__95_, link_o_stitch_0__2__data__94_, link_o_stitch_0__2__data__93_, link_o_stitch_0__2__data__92_, link_o_stitch_0__2__data__91_, link_o_stitch_0__2__data__90_, link_o_stitch_0__2__data__89_, link_o_stitch_0__2__data__88_, link_o_stitch_0__2__data__87_, link_o_stitch_0__2__data__86_, link_o_stitch_0__2__data__85_, link_o_stitch_0__2__data__84_, link_o_stitch_0__2__data__83_, link_o_stitch_0__2__data__82_, link_o_stitch_0__2__data__81_, link_o_stitch_0__2__data__80_, link_o_stitch_0__2__data__79_, link_o_stitch_0__2__data__78_, link_o_stitch_0__2__data__77_, link_o_stitch_0__2__data__76_, link_o_stitch_0__2__data__75_, link_o_stitch_0__2__data__74_, link_o_stitch_0__2__data__73_, link_o_stitch_0__2__data__72_, link_o_stitch_0__2__data__71_, link_o_stitch_0__2__data__70_, link_o_stitch_0__2__data__69_, link_o_stitch_0__2__data__68_, link_o_stitch_0__2__data__67_, link_o_stitch_0__2__data__66_, link_o_stitch_0__2__data__65_, link_o_stitch_0__2__data__64_, link_o_stitch_0__2__data__63_, link_o_stitch_0__2__data__62_, link_o_stitch_0__2__data__61_, link_o_stitch_0__2__data__60_, link_o_stitch_0__2__data__59_, link_o_stitch_0__2__data__58_, link_o_stitch_0__2__data__57_, link_o_stitch_0__2__data__56_, link_o_stitch_0__2__data__55_, link_o_stitch_0__2__data__54_, link_o_stitch_0__2__data__53_, link_o_stitch_0__2__data__52_, link_o_stitch_0__2__data__51_, link_o_stitch_0__2__data__50_, link_o_stitch_0__2__data__49_, link_o_stitch_0__2__data__48_, link_o_stitch_0__2__data__47_, link_o_stitch_0__2__data__46_, link_o_stitch_0__2__data__45_, link_o_stitch_0__2__data__44_, link_o_stitch_0__2__data__43_, link_o_stitch_0__2__data__42_, link_o_stitch_0__2__data__41_, link_o_stitch_0__2__data__40_, link_o_stitch_0__2__data__39_, link_o_stitch_0__2__data__38_, link_o_stitch_0__2__data__37_, link_o_stitch_0__2__data__36_, link_o_stitch_0__2__data__35_, link_o_stitch_0__2__data__34_, link_o_stitch_0__2__data__33_, link_o_stitch_0__2__data__32_, link_o_stitch_0__2__data__31_, link_o_stitch_0__2__data__30_, link_o_stitch_0__2__data__29_, link_o_stitch_0__2__data__28_, link_o_stitch_0__2__data__27_, link_o_stitch_0__2__data__26_, link_o_stitch_0__2__data__25_, link_o_stitch_0__2__data__24_, link_o_stitch_0__2__data__23_, link_o_stitch_0__2__data__22_, link_o_stitch_0__2__data__21_, link_o_stitch_0__2__data__20_, link_o_stitch_0__2__data__19_, link_o_stitch_0__2__data__18_, link_o_stitch_0__2__data__17_, link_o_stitch_0__2__data__16_, link_o_stitch_0__2__data__15_, link_o_stitch_0__2__data__14_, link_o_stitch_0__2__data__13_, link_o_stitch_0__2__data__12_, link_o_stitch_0__2__data__11_, link_o_stitch_0__2__data__10_, link_o_stitch_0__2__data__9_, link_o_stitch_0__2__data__8_, link_o_stitch_0__2__data__7_, link_o_stitch_0__2__data__6_, link_o_stitch_0__2__data__5_, link_o_stitch_0__2__data__4_, link_o_stitch_0__2__data__3_, link_o_stitch_0__2__data__2_, link_o_stitch_0__2__data__1_, link_o_stitch_0__2__data__0_, link_o_stitch_0__1__v_, link_o_stitch_0__1__ready_then_rev_, link_o_stitch_0__1__data__98_, link_o_stitch_0__1__data__97_, link_o_stitch_0__1__data__96_, link_o_stitch_0__1__data__95_, link_o_stitch_0__1__data__94_, link_o_stitch_0__1__data__93_, link_o_stitch_0__1__data__92_, link_o_stitch_0__1__data__91_, link_o_stitch_0__1__data__90_, link_o_stitch_0__1__data__89_, link_o_stitch_0__1__data__88_, link_o_stitch_0__1__data__87_, link_o_stitch_0__1__data__86_, link_o_stitch_0__1__data__85_, link_o_stitch_0__1__data__84_, link_o_stitch_0__1__data__83_, link_o_stitch_0__1__data__82_, link_o_stitch_0__1__data__81_, link_o_stitch_0__1__data__80_, link_o_stitch_0__1__data__79_, link_o_stitch_0__1__data__78_, link_o_stitch_0__1__data__77_, link_o_stitch_0__1__data__76_, link_o_stitch_0__1__data__75_, link_o_stitch_0__1__data__74_, link_o_stitch_0__1__data__73_, link_o_stitch_0__1__data__72_, link_o_stitch_0__1__data__71_, link_o_stitch_0__1__data__70_, link_o_stitch_0__1__data__69_, link_o_stitch_0__1__data__68_, link_o_stitch_0__1__data__67_, link_o_stitch_0__1__data__66_, link_o_stitch_0__1__data__65_, link_o_stitch_0__1__data__64_, link_o_stitch_0__1__data__63_, link_o_stitch_0__1__data__62_, link_o_stitch_0__1__data__61_, link_o_stitch_0__1__data__60_, link_o_stitch_0__1__data__59_, link_o_stitch_0__1__data__58_, link_o_stitch_0__1__data__57_, link_o_stitch_0__1__data__56_, link_o_stitch_0__1__data__55_, link_o_stitch_0__1__data__54_, link_o_stitch_0__1__data__53_, link_o_stitch_0__1__data__52_, link_o_stitch_0__1__data__51_, link_o_stitch_0__1__data__50_, link_o_stitch_0__1__data__49_, link_o_stitch_0__1__data__48_, link_o_stitch_0__1__data__47_, link_o_stitch_0__1__data__46_, link_o_stitch_0__1__data__45_, link_o_stitch_0__1__data__44_, link_o_stitch_0__1__data__43_, link_o_stitch_0__1__data__42_, link_o_stitch_0__1__data__41_, link_o_stitch_0__1__data__40_, link_o_stitch_0__1__data__39_, link_o_stitch_0__1__data__38_, link_o_stitch_0__1__data__37_, link_o_stitch_0__1__data__36_, link_o_stitch_0__1__data__35_, link_o_stitch_0__1__data__34_, link_o_stitch_0__1__data__33_, link_o_stitch_0__1__data__32_, link_o_stitch_0__1__data__31_, link_o_stitch_0__1__data__30_, link_o_stitch_0__1__data__29_, link_o_stitch_0__1__data__28_, link_o_stitch_0__1__data__27_, link_o_stitch_0__1__data__26_, link_o_stitch_0__1__data__25_, link_o_stitch_0__1__data__24_, link_o_stitch_0__1__data__23_, link_o_stitch_0__1__data__22_, link_o_stitch_0__1__data__21_, link_o_stitch_0__1__data__20_, link_o_stitch_0__1__data__19_, link_o_stitch_0__1__data__18_, link_o_stitch_0__1__data__17_, link_o_stitch_0__1__data__16_, link_o_stitch_0__1__data__15_, link_o_stitch_0__1__data__14_, link_o_stitch_0__1__data__13_, link_o_stitch_0__1__data__12_, link_o_stitch_0__1__data__11_, link_o_stitch_0__1__data__10_, link_o_stitch_0__1__data__9_, link_o_stitch_0__1__data__8_, link_o_stitch_0__1__data__7_, link_o_stitch_0__1__data__6_, link_o_stitch_0__1__data__5_, link_o_stitch_0__1__data__4_, link_o_stitch_0__1__data__3_, link_o_stitch_0__1__data__2_, link_o_stitch_0__1__data__1_, link_o_stitch_0__1__data__0_, dst_v_o[0:0], link_o_stitch_0__0__ready_then_rev_, dst_data_o, link_o_stitch_0__0__data__1_, link_o_stitch_0__0__data__0_ }),
    .my_x_i(1'b0),
    .my_y_i(1'b1)
  );


  bsg_mesh_router_buffered_99_1_1_0_5_0d_0_101_00
  rof_1__efi2_fi7_coherence_network_channel_node
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .link_i({ src_v_i[1:1], 1'b0, src_data_i[193:97], 1'b1, src_data_i[193:193], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, link_o_stitch_0__2__v_, link_o_stitch_0__2__ready_then_rev_, link_o_stitch_0__2__data__98_, link_o_stitch_0__2__data__97_, link_o_stitch_0__2__data__96_, link_o_stitch_0__2__data__95_, link_o_stitch_0__2__data__94_, link_o_stitch_0__2__data__93_, link_o_stitch_0__2__data__92_, link_o_stitch_0__2__data__91_, link_o_stitch_0__2__data__90_, link_o_stitch_0__2__data__89_, link_o_stitch_0__2__data__88_, link_o_stitch_0__2__data__87_, link_o_stitch_0__2__data__86_, link_o_stitch_0__2__data__85_, link_o_stitch_0__2__data__84_, link_o_stitch_0__2__data__83_, link_o_stitch_0__2__data__82_, link_o_stitch_0__2__data__81_, link_o_stitch_0__2__data__80_, link_o_stitch_0__2__data__79_, link_o_stitch_0__2__data__78_, link_o_stitch_0__2__data__77_, link_o_stitch_0__2__data__76_, link_o_stitch_0__2__data__75_, link_o_stitch_0__2__data__74_, link_o_stitch_0__2__data__73_, link_o_stitch_0__2__data__72_, link_o_stitch_0__2__data__71_, link_o_stitch_0__2__data__70_, link_o_stitch_0__2__data__69_, link_o_stitch_0__2__data__68_, link_o_stitch_0__2__data__67_, link_o_stitch_0__2__data__66_, link_o_stitch_0__2__data__65_, link_o_stitch_0__2__data__64_, link_o_stitch_0__2__data__63_, link_o_stitch_0__2__data__62_, link_o_stitch_0__2__data__61_, link_o_stitch_0__2__data__60_, link_o_stitch_0__2__data__59_, link_o_stitch_0__2__data__58_, link_o_stitch_0__2__data__57_, link_o_stitch_0__2__data__56_, link_o_stitch_0__2__data__55_, link_o_stitch_0__2__data__54_, link_o_stitch_0__2__data__53_, link_o_stitch_0__2__data__52_, link_o_stitch_0__2__data__51_, link_o_stitch_0__2__data__50_, link_o_stitch_0__2__data__49_, link_o_stitch_0__2__data__48_, link_o_stitch_0__2__data__47_, link_o_stitch_0__2__data__46_, link_o_stitch_0__2__data__45_, link_o_stitch_0__2__data__44_, link_o_stitch_0__2__data__43_, link_o_stitch_0__2__data__42_, link_o_stitch_0__2__data__41_, link_o_stitch_0__2__data__40_, link_o_stitch_0__2__data__39_, link_o_stitch_0__2__data__38_, link_o_stitch_0__2__data__37_, link_o_stitch_0__2__data__36_, link_o_stitch_0__2__data__35_, link_o_stitch_0__2__data__34_, link_o_stitch_0__2__data__33_, link_o_stitch_0__2__data__32_, link_o_stitch_0__2__data__31_, link_o_stitch_0__2__data__30_, link_o_stitch_0__2__data__29_, link_o_stitch_0__2__data__28_, link_o_stitch_0__2__data__27_, link_o_stitch_0__2__data__26_, link_o_stitch_0__2__data__25_, link_o_stitch_0__2__data__24_, link_o_stitch_0__2__data__23_, link_o_stitch_0__2__data__22_, link_o_stitch_0__2__data__21_, link_o_stitch_0__2__data__20_, link_o_stitch_0__2__data__19_, link_o_stitch_0__2__data__18_, link_o_stitch_0__2__data__17_, link_o_stitch_0__2__data__16_, link_o_stitch_0__2__data__15_, link_o_stitch_0__2__data__14_, link_o_stitch_0__2__data__13_, link_o_stitch_0__2__data__12_, link_o_stitch_0__2__data__11_, link_o_stitch_0__2__data__10_, link_o_stitch_0__2__data__9_, link_o_stitch_0__2__data__8_, link_o_stitch_0__2__data__7_, link_o_stitch_0__2__data__6_, link_o_stitch_0__2__data__5_, link_o_stitch_0__2__data__4_, link_o_stitch_0__2__data__3_, link_o_stitch_0__2__data__2_, link_o_stitch_0__2__data__1_, link_o_stitch_0__2__data__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .link_o({ link_o_stitch_1__4__v_, src_ready_o[1:1], link_o_stitch_1__4__data__98_, link_o_stitch_1__4__data__97_, link_o_stitch_1__4__data__96_, link_o_stitch_1__4__data__95_, link_o_stitch_1__4__data__94_, link_o_stitch_1__4__data__93_, link_o_stitch_1__4__data__92_, link_o_stitch_1__4__data__91_, link_o_stitch_1__4__data__90_, link_o_stitch_1__4__data__89_, link_o_stitch_1__4__data__88_, link_o_stitch_1__4__data__87_, link_o_stitch_1__4__data__86_, link_o_stitch_1__4__data__85_, link_o_stitch_1__4__data__84_, link_o_stitch_1__4__data__83_, link_o_stitch_1__4__data__82_, link_o_stitch_1__4__data__81_, link_o_stitch_1__4__data__80_, link_o_stitch_1__4__data__79_, link_o_stitch_1__4__data__78_, link_o_stitch_1__4__data__77_, link_o_stitch_1__4__data__76_, link_o_stitch_1__4__data__75_, link_o_stitch_1__4__data__74_, link_o_stitch_1__4__data__73_, link_o_stitch_1__4__data__72_, link_o_stitch_1__4__data__71_, link_o_stitch_1__4__data__70_, link_o_stitch_1__4__data__69_, link_o_stitch_1__4__data__68_, link_o_stitch_1__4__data__67_, link_o_stitch_1__4__data__66_, link_o_stitch_1__4__data__65_, link_o_stitch_1__4__data__64_, link_o_stitch_1__4__data__63_, link_o_stitch_1__4__data__62_, link_o_stitch_1__4__data__61_, link_o_stitch_1__4__data__60_, link_o_stitch_1__4__data__59_, link_o_stitch_1__4__data__58_, link_o_stitch_1__4__data__57_, link_o_stitch_1__4__data__56_, link_o_stitch_1__4__data__55_, link_o_stitch_1__4__data__54_, link_o_stitch_1__4__data__53_, link_o_stitch_1__4__data__52_, link_o_stitch_1__4__data__51_, link_o_stitch_1__4__data__50_, link_o_stitch_1__4__data__49_, link_o_stitch_1__4__data__48_, link_o_stitch_1__4__data__47_, link_o_stitch_1__4__data__46_, link_o_stitch_1__4__data__45_, link_o_stitch_1__4__data__44_, link_o_stitch_1__4__data__43_, link_o_stitch_1__4__data__42_, link_o_stitch_1__4__data__41_, link_o_stitch_1__4__data__40_, link_o_stitch_1__4__data__39_, link_o_stitch_1__4__data__38_, link_o_stitch_1__4__data__37_, link_o_stitch_1__4__data__36_, link_o_stitch_1__4__data__35_, link_o_stitch_1__4__data__34_, link_o_stitch_1__4__data__33_, link_o_stitch_1__4__data__32_, link_o_stitch_1__4__data__31_, link_o_stitch_1__4__data__30_, link_o_stitch_1__4__data__29_, link_o_stitch_1__4__data__28_, link_o_stitch_1__4__data__27_, link_o_stitch_1__4__data__26_, link_o_stitch_1__4__data__25_, link_o_stitch_1__4__data__24_, link_o_stitch_1__4__data__23_, link_o_stitch_1__4__data__22_, link_o_stitch_1__4__data__21_, link_o_stitch_1__4__data__20_, link_o_stitch_1__4__data__19_, link_o_stitch_1__4__data__18_, link_o_stitch_1__4__data__17_, link_o_stitch_1__4__data__16_, link_o_stitch_1__4__data__15_, link_o_stitch_1__4__data__14_, link_o_stitch_1__4__data__13_, link_o_stitch_1__4__data__12_, link_o_stitch_1__4__data__11_, link_o_stitch_1__4__data__10_, link_o_stitch_1__4__data__9_, link_o_stitch_1__4__data__8_, link_o_stitch_1__4__data__7_, link_o_stitch_1__4__data__6_, link_o_stitch_1__4__data__5_, link_o_stitch_1__4__data__4_, link_o_stitch_1__4__data__3_, link_o_stitch_1__4__data__2_, link_o_stitch_1__4__data__1_, link_o_stitch_1__4__data__0_, link_o_stitch_1__3__v_, link_o_stitch_1__3__ready_then_rev_, link_o_stitch_1__3__data__98_, link_o_stitch_1__3__data__97_, link_o_stitch_1__3__data__96_, link_o_stitch_1__3__data__95_, link_o_stitch_1__3__data__94_, link_o_stitch_1__3__data__93_, link_o_stitch_1__3__data__92_, link_o_stitch_1__3__data__91_, link_o_stitch_1__3__data__90_, link_o_stitch_1__3__data__89_, link_o_stitch_1__3__data__88_, link_o_stitch_1__3__data__87_, link_o_stitch_1__3__data__86_, link_o_stitch_1__3__data__85_, link_o_stitch_1__3__data__84_, link_o_stitch_1__3__data__83_, link_o_stitch_1__3__data__82_, link_o_stitch_1__3__data__81_, link_o_stitch_1__3__data__80_, link_o_stitch_1__3__data__79_, link_o_stitch_1__3__data__78_, link_o_stitch_1__3__data__77_, link_o_stitch_1__3__data__76_, link_o_stitch_1__3__data__75_, link_o_stitch_1__3__data__74_, link_o_stitch_1__3__data__73_, link_o_stitch_1__3__data__72_, link_o_stitch_1__3__data__71_, link_o_stitch_1__3__data__70_, link_o_stitch_1__3__data__69_, link_o_stitch_1__3__data__68_, link_o_stitch_1__3__data__67_, link_o_stitch_1__3__data__66_, link_o_stitch_1__3__data__65_, link_o_stitch_1__3__data__64_, link_o_stitch_1__3__data__63_, link_o_stitch_1__3__data__62_, link_o_stitch_1__3__data__61_, link_o_stitch_1__3__data__60_, link_o_stitch_1__3__data__59_, link_o_stitch_1__3__data__58_, link_o_stitch_1__3__data__57_, link_o_stitch_1__3__data__56_, link_o_stitch_1__3__data__55_, link_o_stitch_1__3__data__54_, link_o_stitch_1__3__data__53_, link_o_stitch_1__3__data__52_, link_o_stitch_1__3__data__51_, link_o_stitch_1__3__data__50_, link_o_stitch_1__3__data__49_, link_o_stitch_1__3__data__48_, link_o_stitch_1__3__data__47_, link_o_stitch_1__3__data__46_, link_o_stitch_1__3__data__45_, link_o_stitch_1__3__data__44_, link_o_stitch_1__3__data__43_, link_o_stitch_1__3__data__42_, link_o_stitch_1__3__data__41_, link_o_stitch_1__3__data__40_, link_o_stitch_1__3__data__39_, link_o_stitch_1__3__data__38_, link_o_stitch_1__3__data__37_, link_o_stitch_1__3__data__36_, link_o_stitch_1__3__data__35_, link_o_stitch_1__3__data__34_, link_o_stitch_1__3__data__33_, link_o_stitch_1__3__data__32_, link_o_stitch_1__3__data__31_, link_o_stitch_1__3__data__30_, link_o_stitch_1__3__data__29_, link_o_stitch_1__3__data__28_, link_o_stitch_1__3__data__27_, link_o_stitch_1__3__data__26_, link_o_stitch_1__3__data__25_, link_o_stitch_1__3__data__24_, link_o_stitch_1__3__data__23_, link_o_stitch_1__3__data__22_, link_o_stitch_1__3__data__21_, link_o_stitch_1__3__data__20_, link_o_stitch_1__3__data__19_, link_o_stitch_1__3__data__18_, link_o_stitch_1__3__data__17_, link_o_stitch_1__3__data__16_, link_o_stitch_1__3__data__15_, link_o_stitch_1__3__data__14_, link_o_stitch_1__3__data__13_, link_o_stitch_1__3__data__12_, link_o_stitch_1__3__data__11_, link_o_stitch_1__3__data__10_, link_o_stitch_1__3__data__9_, link_o_stitch_1__3__data__8_, link_o_stitch_1__3__data__7_, link_o_stitch_1__3__data__6_, link_o_stitch_1__3__data__5_, link_o_stitch_1__3__data__4_, link_o_stitch_1__3__data__3_, link_o_stitch_1__3__data__2_, link_o_stitch_1__3__data__1_, link_o_stitch_1__3__data__0_, link_o_stitch_1__2__v_, link_o_stitch_1__2__ready_then_rev_, link_o_stitch_1__2__data__98_, link_o_stitch_1__2__data__97_, link_o_stitch_1__2__data__96_, link_o_stitch_1__2__data__95_, link_o_stitch_1__2__data__94_, link_o_stitch_1__2__data__93_, link_o_stitch_1__2__data__92_, link_o_stitch_1__2__data__91_, link_o_stitch_1__2__data__90_, link_o_stitch_1__2__data__89_, link_o_stitch_1__2__data__88_, link_o_stitch_1__2__data__87_, link_o_stitch_1__2__data__86_, link_o_stitch_1__2__data__85_, link_o_stitch_1__2__data__84_, link_o_stitch_1__2__data__83_, link_o_stitch_1__2__data__82_, link_o_stitch_1__2__data__81_, link_o_stitch_1__2__data__80_, link_o_stitch_1__2__data__79_, link_o_stitch_1__2__data__78_, link_o_stitch_1__2__data__77_, link_o_stitch_1__2__data__76_, link_o_stitch_1__2__data__75_, link_o_stitch_1__2__data__74_, link_o_stitch_1__2__data__73_, link_o_stitch_1__2__data__72_, link_o_stitch_1__2__data__71_, link_o_stitch_1__2__data__70_, link_o_stitch_1__2__data__69_, link_o_stitch_1__2__data__68_, link_o_stitch_1__2__data__67_, link_o_stitch_1__2__data__66_, link_o_stitch_1__2__data__65_, link_o_stitch_1__2__data__64_, link_o_stitch_1__2__data__63_, link_o_stitch_1__2__data__62_, link_o_stitch_1__2__data__61_, link_o_stitch_1__2__data__60_, link_o_stitch_1__2__data__59_, link_o_stitch_1__2__data__58_, link_o_stitch_1__2__data__57_, link_o_stitch_1__2__data__56_, link_o_stitch_1__2__data__55_, link_o_stitch_1__2__data__54_, link_o_stitch_1__2__data__53_, link_o_stitch_1__2__data__52_, link_o_stitch_1__2__data__51_, link_o_stitch_1__2__data__50_, link_o_stitch_1__2__data__49_, link_o_stitch_1__2__data__48_, link_o_stitch_1__2__data__47_, link_o_stitch_1__2__data__46_, link_o_stitch_1__2__data__45_, link_o_stitch_1__2__data__44_, link_o_stitch_1__2__data__43_, link_o_stitch_1__2__data__42_, link_o_stitch_1__2__data__41_, link_o_stitch_1__2__data__40_, link_o_stitch_1__2__data__39_, link_o_stitch_1__2__data__38_, link_o_stitch_1__2__data__37_, link_o_stitch_1__2__data__36_, link_o_stitch_1__2__data__35_, link_o_stitch_1__2__data__34_, link_o_stitch_1__2__data__33_, link_o_stitch_1__2__data__32_, link_o_stitch_1__2__data__31_, link_o_stitch_1__2__data__30_, link_o_stitch_1__2__data__29_, link_o_stitch_1__2__data__28_, link_o_stitch_1__2__data__27_, link_o_stitch_1__2__data__26_, link_o_stitch_1__2__data__25_, link_o_stitch_1__2__data__24_, link_o_stitch_1__2__data__23_, link_o_stitch_1__2__data__22_, link_o_stitch_1__2__data__21_, link_o_stitch_1__2__data__20_, link_o_stitch_1__2__data__19_, link_o_stitch_1__2__data__18_, link_o_stitch_1__2__data__17_, link_o_stitch_1__2__data__16_, link_o_stitch_1__2__data__15_, link_o_stitch_1__2__data__14_, link_o_stitch_1__2__data__13_, link_o_stitch_1__2__data__12_, link_o_stitch_1__2__data__11_, link_o_stitch_1__2__data__10_, link_o_stitch_1__2__data__9_, link_o_stitch_1__2__data__8_, link_o_stitch_1__2__data__7_, link_o_stitch_1__2__data__6_, link_o_stitch_1__2__data__5_, link_o_stitch_1__2__data__4_, link_o_stitch_1__2__data__3_, link_o_stitch_1__2__data__2_, link_o_stitch_1__2__data__1_, link_o_stitch_1__2__data__0_, link_i_stitch_0__2__v_, link_i_stitch_0__2__ready_then_rev_, link_i_stitch_0__2__data__98_, link_i_stitch_0__2__data__97_, link_i_stitch_0__2__data__96_, link_i_stitch_0__2__data__95_, link_i_stitch_0__2__data__94_, link_i_stitch_0__2__data__93_, link_i_stitch_0__2__data__92_, link_i_stitch_0__2__data__91_, link_i_stitch_0__2__data__90_, link_i_stitch_0__2__data__89_, link_i_stitch_0__2__data__88_, link_i_stitch_0__2__data__87_, link_i_stitch_0__2__data__86_, link_i_stitch_0__2__data__85_, link_i_stitch_0__2__data__84_, link_i_stitch_0__2__data__83_, link_i_stitch_0__2__data__82_, link_i_stitch_0__2__data__81_, link_i_stitch_0__2__data__80_, link_i_stitch_0__2__data__79_, link_i_stitch_0__2__data__78_, link_i_stitch_0__2__data__77_, link_i_stitch_0__2__data__76_, link_i_stitch_0__2__data__75_, link_i_stitch_0__2__data__74_, link_i_stitch_0__2__data__73_, link_i_stitch_0__2__data__72_, link_i_stitch_0__2__data__71_, link_i_stitch_0__2__data__70_, link_i_stitch_0__2__data__69_, link_i_stitch_0__2__data__68_, link_i_stitch_0__2__data__67_, link_i_stitch_0__2__data__66_, link_i_stitch_0__2__data__65_, link_i_stitch_0__2__data__64_, link_i_stitch_0__2__data__63_, link_i_stitch_0__2__data__62_, link_i_stitch_0__2__data__61_, link_i_stitch_0__2__data__60_, link_i_stitch_0__2__data__59_, link_i_stitch_0__2__data__58_, link_i_stitch_0__2__data__57_, link_i_stitch_0__2__data__56_, link_i_stitch_0__2__data__55_, link_i_stitch_0__2__data__54_, link_i_stitch_0__2__data__53_, link_i_stitch_0__2__data__52_, link_i_stitch_0__2__data__51_, link_i_stitch_0__2__data__50_, link_i_stitch_0__2__data__49_, link_i_stitch_0__2__data__48_, link_i_stitch_0__2__data__47_, link_i_stitch_0__2__data__46_, link_i_stitch_0__2__data__45_, link_i_stitch_0__2__data__44_, link_i_stitch_0__2__data__43_, link_i_stitch_0__2__data__42_, link_i_stitch_0__2__data__41_, link_i_stitch_0__2__data__40_, link_i_stitch_0__2__data__39_, link_i_stitch_0__2__data__38_, link_i_stitch_0__2__data__37_, link_i_stitch_0__2__data__36_, link_i_stitch_0__2__data__35_, link_i_stitch_0__2__data__34_, link_i_stitch_0__2__data__33_, link_i_stitch_0__2__data__32_, link_i_stitch_0__2__data__31_, link_i_stitch_0__2__data__30_, link_i_stitch_0__2__data__29_, link_i_stitch_0__2__data__28_, link_i_stitch_0__2__data__27_, link_i_stitch_0__2__data__26_, link_i_stitch_0__2__data__25_, link_i_stitch_0__2__data__24_, link_i_stitch_0__2__data__23_, link_i_stitch_0__2__data__22_, link_i_stitch_0__2__data__21_, link_i_stitch_0__2__data__20_, link_i_stitch_0__2__data__19_, link_i_stitch_0__2__data__18_, link_i_stitch_0__2__data__17_, link_i_stitch_0__2__data__16_, link_i_stitch_0__2__data__15_, link_i_stitch_0__2__data__14_, link_i_stitch_0__2__data__13_, link_i_stitch_0__2__data__12_, link_i_stitch_0__2__data__11_, link_i_stitch_0__2__data__10_, link_i_stitch_0__2__data__9_, link_i_stitch_0__2__data__8_, link_i_stitch_0__2__data__7_, link_i_stitch_0__2__data__6_, link_i_stitch_0__2__data__5_, link_i_stitch_0__2__data__4_, link_i_stitch_0__2__data__3_, link_i_stitch_0__2__data__2_, link_i_stitch_0__2__data__1_, link_i_stitch_0__2__data__0_, link_o_stitch_1__0__v_, link_o_stitch_1__0__ready_then_rev_, link_o_stitch_1__0__data__98_, link_o_stitch_1__0__data__97_, link_o_stitch_1__0__data__96_, link_o_stitch_1__0__data__95_, link_o_stitch_1__0__data__94_, link_o_stitch_1__0__data__93_, link_o_stitch_1__0__data__92_, link_o_stitch_1__0__data__91_, link_o_stitch_1__0__data__90_, link_o_stitch_1__0__data__89_, link_o_stitch_1__0__data__88_, link_o_stitch_1__0__data__87_, link_o_stitch_1__0__data__86_, link_o_stitch_1__0__data__85_, link_o_stitch_1__0__data__84_, link_o_stitch_1__0__data__83_, link_o_stitch_1__0__data__82_, link_o_stitch_1__0__data__81_, link_o_stitch_1__0__data__80_, link_o_stitch_1__0__data__79_, link_o_stitch_1__0__data__78_, link_o_stitch_1__0__data__77_, link_o_stitch_1__0__data__76_, link_o_stitch_1__0__data__75_, link_o_stitch_1__0__data__74_, link_o_stitch_1__0__data__73_, link_o_stitch_1__0__data__72_, link_o_stitch_1__0__data__71_, link_o_stitch_1__0__data__70_, link_o_stitch_1__0__data__69_, link_o_stitch_1__0__data__68_, link_o_stitch_1__0__data__67_, link_o_stitch_1__0__data__66_, link_o_stitch_1__0__data__65_, link_o_stitch_1__0__data__64_, link_o_stitch_1__0__data__63_, link_o_stitch_1__0__data__62_, link_o_stitch_1__0__data__61_, link_o_stitch_1__0__data__60_, link_o_stitch_1__0__data__59_, link_o_stitch_1__0__data__58_, link_o_stitch_1__0__data__57_, link_o_stitch_1__0__data__56_, link_o_stitch_1__0__data__55_, link_o_stitch_1__0__data__54_, link_o_stitch_1__0__data__53_, link_o_stitch_1__0__data__52_, link_o_stitch_1__0__data__51_, link_o_stitch_1__0__data__50_, link_o_stitch_1__0__data__49_, link_o_stitch_1__0__data__48_, link_o_stitch_1__0__data__47_, link_o_stitch_1__0__data__46_, link_o_stitch_1__0__data__45_, link_o_stitch_1__0__data__44_, link_o_stitch_1__0__data__43_, link_o_stitch_1__0__data__42_, link_o_stitch_1__0__data__41_, link_o_stitch_1__0__data__40_, link_o_stitch_1__0__data__39_, link_o_stitch_1__0__data__38_, link_o_stitch_1__0__data__37_, link_o_stitch_1__0__data__36_, link_o_stitch_1__0__data__35_, link_o_stitch_1__0__data__34_, link_o_stitch_1__0__data__33_, link_o_stitch_1__0__data__32_, link_o_stitch_1__0__data__31_, link_o_stitch_1__0__data__30_, link_o_stitch_1__0__data__29_, link_o_stitch_1__0__data__28_, link_o_stitch_1__0__data__27_, link_o_stitch_1__0__data__26_, link_o_stitch_1__0__data__25_, link_o_stitch_1__0__data__24_, link_o_stitch_1__0__data__23_, link_o_stitch_1__0__data__22_, link_o_stitch_1__0__data__21_, link_o_stitch_1__0__data__20_, link_o_stitch_1__0__data__19_, link_o_stitch_1__0__data__18_, link_o_stitch_1__0__data__17_, link_o_stitch_1__0__data__16_, link_o_stitch_1__0__data__15_, link_o_stitch_1__0__data__14_, link_o_stitch_1__0__data__13_, link_o_stitch_1__0__data__12_, link_o_stitch_1__0__data__11_, link_o_stitch_1__0__data__10_, link_o_stitch_1__0__data__9_, link_o_stitch_1__0__data__8_, link_o_stitch_1__0__data__7_, link_o_stitch_1__0__data__6_, link_o_stitch_1__0__data__5_, link_o_stitch_1__0__data__4_, link_o_stitch_1__0__data__3_, link_o_stitch_1__0__data__2_, link_o_stitch_1__0__data__1_, link_o_stitch_1__0__data__0_ }),
    .my_x_i(1'b1),
    .my_y_i(1'b1)
  );


endmodule



module bsg_mem_p28
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [27:0] w_data_i;
  input [0:0] r_addr_i;
  output [27:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [27:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  reg [55:0] mem;
  assign r_data_o[27] = (N3)? mem[27] :
                        (N0)? mem[55] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[26] = (N3)? mem[26] :
                        (N0)? mem[54] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] :
                        (N0)? mem[53] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] :
                        (N0)? mem[52] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] :
                        (N0)? mem[51] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] :
                        (N0)? mem[50] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] :
                        (N0)? mem[49] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] :
                        (N0)? mem[48] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] :
                        (N0)? mem[47] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] :
                        (N0)? mem[46] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] :
                        (N0)? mem[45] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] :
                        (N0)? mem[44] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] :
                        (N0)? mem[43] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] :
                        (N0)? mem[42] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] :
                        (N0)? mem[41] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] :
                        (N0)? mem[40] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] :
                        (N0)? mem[39] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] :
                        (N0)? mem[38] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] :
                       (N0)? mem[37] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] :
                       (N0)? mem[36] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] :
                       (N0)? mem[35] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] :
                       (N0)? mem[34] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] :
                       (N0)? mem[33] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] :
                       (N0)? mem[32] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] :
                       (N0)? mem[31] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] :
                       (N0)? mem[30] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] :
                       (N0)? mem[29] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] :
                       (N0)? mem[28] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } :
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      { mem[55:28] } <= { w_data_i[27:0] };
    end
    if(N7) begin
      { mem[27:0] } <= { w_data_i[27:0] };
    end
  end


endmodule



module bsg_mem_1r1w_width_p28_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [27:0] w_data_i;
  input [0:0] r_addr_i;
  output [27:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [27:0] r_data_o;

  bsg_mem_p28
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p28
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [27:0] data_i;
  output [27:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [27:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p28_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 :
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 :
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 :
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 :
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 :
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 :
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end
    if(N9) begin
      tail_r <= N10;
    end
    if(N11) begin
      head_r <= N12;
    end
  end


endmodule



module bsg_mux_one_hot_width_p28_els_p4
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [111:0] data_i;
  input [3:0] sel_one_hot_i;
  output [27:0] data_o;
  wire [27:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55;
  wire [111:0] data_masked;
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[1];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[1];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[1];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[1];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[1];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[1];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[1];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[1];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[1];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[1];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[1];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[1];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[1];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[1];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[1];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[1];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[1];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[1];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[1];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[1];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[1];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[1];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[1];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[1];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[1];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[1];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[1];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[2];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[2];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[2];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[2];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[2];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[2];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[2];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[2];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[2];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[2];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[2];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[2];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[2];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[2];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[2];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[2];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[2];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[2];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[2];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[2];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[2];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[2];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[2];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[2];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[2];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[2];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[2];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[2];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[3];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[3];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[3];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[3];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[3];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[3];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[3];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[3];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[3];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[3];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[3];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[3];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[3];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[3];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[3];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[3];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[3];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[3];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[3];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[3];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[3];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[3];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[3];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[3];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[3];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[3];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[3];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[3];
  assign data_o[0] = N1 | data_masked[0];
  assign N1 = N0 | data_masked[28];
  assign N0 = data_masked[84] | data_masked[56];
  assign data_o[1] = N3 | data_masked[1];
  assign N3 = N2 | data_masked[29];
  assign N2 = data_masked[85] | data_masked[57];
  assign data_o[2] = N5 | data_masked[2];
  assign N5 = N4 | data_masked[30];
  assign N4 = data_masked[86] | data_masked[58];
  assign data_o[3] = N7 | data_masked[3];
  assign N7 = N6 | data_masked[31];
  assign N6 = data_masked[87] | data_masked[59];
  assign data_o[4] = N9 | data_masked[4];
  assign N9 = N8 | data_masked[32];
  assign N8 = data_masked[88] | data_masked[60];
  assign data_o[5] = N11 | data_masked[5];
  assign N11 = N10 | data_masked[33];
  assign N10 = data_masked[89] | data_masked[61];
  assign data_o[6] = N13 | data_masked[6];
  assign N13 = N12 | data_masked[34];
  assign N12 = data_masked[90] | data_masked[62];
  assign data_o[7] = N15 | data_masked[7];
  assign N15 = N14 | data_masked[35];
  assign N14 = data_masked[91] | data_masked[63];
  assign data_o[8] = N17 | data_masked[8];
  assign N17 = N16 | data_masked[36];
  assign N16 = data_masked[92] | data_masked[64];
  assign data_o[9] = N19 | data_masked[9];
  assign N19 = N18 | data_masked[37];
  assign N18 = data_masked[93] | data_masked[65];
  assign data_o[10] = N21 | data_masked[10];
  assign N21 = N20 | data_masked[38];
  assign N20 = data_masked[94] | data_masked[66];
  assign data_o[11] = N23 | data_masked[11];
  assign N23 = N22 | data_masked[39];
  assign N22 = data_masked[95] | data_masked[67];
  assign data_o[12] = N25 | data_masked[12];
  assign N25 = N24 | data_masked[40];
  assign N24 = data_masked[96] | data_masked[68];
  assign data_o[13] = N27 | data_masked[13];
  assign N27 = N26 | data_masked[41];
  assign N26 = data_masked[97] | data_masked[69];
  assign data_o[14] = N29 | data_masked[14];
  assign N29 = N28 | data_masked[42];
  assign N28 = data_masked[98] | data_masked[70];
  assign data_o[15] = N31 | data_masked[15];
  assign N31 = N30 | data_masked[43];
  assign N30 = data_masked[99] | data_masked[71];
  assign data_o[16] = N33 | data_masked[16];
  assign N33 = N32 | data_masked[44];
  assign N32 = data_masked[100] | data_masked[72];
  assign data_o[17] = N35 | data_masked[17];
  assign N35 = N34 | data_masked[45];
  assign N34 = data_masked[101] | data_masked[73];
  assign data_o[18] = N37 | data_masked[18];
  assign N37 = N36 | data_masked[46];
  assign N36 = data_masked[102] | data_masked[74];
  assign data_o[19] = N39 | data_masked[19];
  assign N39 = N38 | data_masked[47];
  assign N38 = data_masked[103] | data_masked[75];
  assign data_o[20] = N41 | data_masked[20];
  assign N41 = N40 | data_masked[48];
  assign N40 = data_masked[104] | data_masked[76];
  assign data_o[21] = N43 | data_masked[21];
  assign N43 = N42 | data_masked[49];
  assign N42 = data_masked[105] | data_masked[77];
  assign data_o[22] = N45 | data_masked[22];
  assign N45 = N44 | data_masked[50];
  assign N44 = data_masked[106] | data_masked[78];
  assign data_o[23] = N47 | data_masked[23];
  assign N47 = N46 | data_masked[51];
  assign N46 = data_masked[107] | data_masked[79];
  assign data_o[24] = N49 | data_masked[24];
  assign N49 = N48 | data_masked[52];
  assign N48 = data_masked[108] | data_masked[80];
  assign data_o[25] = N51 | data_masked[25];
  assign N51 = N50 | data_masked[53];
  assign N50 = data_masked[109] | data_masked[81];
  assign data_o[26] = N53 | data_masked[26];
  assign N53 = N52 | data_masked[54];
  assign N52 = data_masked[110] | data_masked[82];
  assign data_o[27] = N55 | data_masked[27];
  assign N55 = N54 | data_masked[55];
  assign N54 = data_masked[111] | data_masked[83];

endmodule



module bsg_mux_one_hot_width_p28_els_p2
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [55:0] data_i;
  input [1:0] sel_one_hot_i;
  output [27:0] data_o;
  wire [27:0] data_o;
  wire [55:0] data_masked;
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[1];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[1];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[1];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[1];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[1];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[1];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[1];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[1];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[1];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[1];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[1];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[1];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[1];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[1];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[1];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[1];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[1];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[1];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[1];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[1];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[1];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[1];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[1];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[1];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[1];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[1];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[1];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[1];
  assign data_o[0] = data_masked[28] | data_masked[0];
  assign data_o[1] = data_masked[29] | data_masked[1];
  assign data_o[2] = data_masked[30] | data_masked[2];
  assign data_o[3] = data_masked[31] | data_masked[3];
  assign data_o[4] = data_masked[32] | data_masked[4];
  assign data_o[5] = data_masked[33] | data_masked[5];
  assign data_o[6] = data_masked[34] | data_masked[6];
  assign data_o[7] = data_masked[35] | data_masked[7];
  assign data_o[8] = data_masked[36] | data_masked[8];
  assign data_o[9] = data_masked[37] | data_masked[9];
  assign data_o[10] = data_masked[38] | data_masked[10];
  assign data_o[11] = data_masked[39] | data_masked[11];
  assign data_o[12] = data_masked[40] | data_masked[12];
  assign data_o[13] = data_masked[41] | data_masked[13];
  assign data_o[14] = data_masked[42] | data_masked[14];
  assign data_o[15] = data_masked[43] | data_masked[15];
  assign data_o[16] = data_masked[44] | data_masked[16];
  assign data_o[17] = data_masked[45] | data_masked[17];
  assign data_o[18] = data_masked[46] | data_masked[18];
  assign data_o[19] = data_masked[47] | data_masked[19];
  assign data_o[20] = data_masked[48] | data_masked[20];
  assign data_o[21] = data_masked[49] | data_masked[21];
  assign data_o[22] = data_masked[50] | data_masked[22];
  assign data_o[23] = data_masked[51] | data_masked[23];
  assign data_o[24] = data_masked[52] | data_masked[24];
  assign data_o[25] = data_masked[53] | data_masked[25];
  assign data_o[26] = data_masked[54] | data_masked[26];
  assign data_o[27] = data_masked[55] | data_masked[27];

endmodule



module bsg_mux_one_hot_width_p28_els_p5
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [139:0] data_i;
  input [4:0] sel_one_hot_i;
  output [27:0] data_o;
  wire [27:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83;
  wire [139:0] data_masked;
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[1];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[1];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[1];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[1];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[1];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[1];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[1];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[1];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[1];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[1];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[1];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[1];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[1];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[1];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[1];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[1];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[1];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[1];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[1];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[1];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[1];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[1];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[1];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[1];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[1];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[1];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[1];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[2];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[2];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[2];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[2];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[2];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[2];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[2];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[2];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[2];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[2];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[2];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[2];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[2];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[2];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[2];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[2];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[2];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[2];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[2];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[2];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[2];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[2];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[2];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[2];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[2];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[2];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[2];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[2];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[3];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[3];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[3];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[3];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[3];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[3];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[3];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[3];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[3];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[3];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[3];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[3];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[3];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[3];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[3];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[3];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[3];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[3];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[3];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[3];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[3];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[3];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[3];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[3];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[3];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[3];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[3];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[3];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[4];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[4];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[4];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[4];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[4];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[4];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[4];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[4];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[4];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[4];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[4];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[4];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[4];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[4];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[4];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[4];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[4];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[4];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[4];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[4];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[4];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[4];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[4];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[4];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[4];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[4];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[4];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[4];
  assign data_o[0] = N2 | data_masked[0];
  assign N2 = N1 | data_masked[28];
  assign N1 = N0 | data_masked[56];
  assign N0 = data_masked[112] | data_masked[84];
  assign data_o[1] = N5 | data_masked[1];
  assign N5 = N4 | data_masked[29];
  assign N4 = N3 | data_masked[57];
  assign N3 = data_masked[113] | data_masked[85];
  assign data_o[2] = N8 | data_masked[2];
  assign N8 = N7 | data_masked[30];
  assign N7 = N6 | data_masked[58];
  assign N6 = data_masked[114] | data_masked[86];
  assign data_o[3] = N11 | data_masked[3];
  assign N11 = N10 | data_masked[31];
  assign N10 = N9 | data_masked[59];
  assign N9 = data_masked[115] | data_masked[87];
  assign data_o[4] = N14 | data_masked[4];
  assign N14 = N13 | data_masked[32];
  assign N13 = N12 | data_masked[60];
  assign N12 = data_masked[116] | data_masked[88];
  assign data_o[5] = N17 | data_masked[5];
  assign N17 = N16 | data_masked[33];
  assign N16 = N15 | data_masked[61];
  assign N15 = data_masked[117] | data_masked[89];
  assign data_o[6] = N20 | data_masked[6];
  assign N20 = N19 | data_masked[34];
  assign N19 = N18 | data_masked[62];
  assign N18 = data_masked[118] | data_masked[90];
  assign data_o[7] = N23 | data_masked[7];
  assign N23 = N22 | data_masked[35];
  assign N22 = N21 | data_masked[63];
  assign N21 = data_masked[119] | data_masked[91];
  assign data_o[8] = N26 | data_masked[8];
  assign N26 = N25 | data_masked[36];
  assign N25 = N24 | data_masked[64];
  assign N24 = data_masked[120] | data_masked[92];
  assign data_o[9] = N29 | data_masked[9];
  assign N29 = N28 | data_masked[37];
  assign N28 = N27 | data_masked[65];
  assign N27 = data_masked[121] | data_masked[93];
  assign data_o[10] = N32 | data_masked[10];
  assign N32 = N31 | data_masked[38];
  assign N31 = N30 | data_masked[66];
  assign N30 = data_masked[122] | data_masked[94];
  assign data_o[11] = N35 | data_masked[11];
  assign N35 = N34 | data_masked[39];
  assign N34 = N33 | data_masked[67];
  assign N33 = data_masked[123] | data_masked[95];
  assign data_o[12] = N38 | data_masked[12];
  assign N38 = N37 | data_masked[40];
  assign N37 = N36 | data_masked[68];
  assign N36 = data_masked[124] | data_masked[96];
  assign data_o[13] = N41 | data_masked[13];
  assign N41 = N40 | data_masked[41];
  assign N40 = N39 | data_masked[69];
  assign N39 = data_masked[125] | data_masked[97];
  assign data_o[14] = N44 | data_masked[14];
  assign N44 = N43 | data_masked[42];
  assign N43 = N42 | data_masked[70];
  assign N42 = data_masked[126] | data_masked[98];
  assign data_o[15] = N47 | data_masked[15];
  assign N47 = N46 | data_masked[43];
  assign N46 = N45 | data_masked[71];
  assign N45 = data_masked[127] | data_masked[99];
  assign data_o[16] = N50 | data_masked[16];
  assign N50 = N49 | data_masked[44];
  assign N49 = N48 | data_masked[72];
  assign N48 = data_masked[128] | data_masked[100];
  assign data_o[17] = N53 | data_masked[17];
  assign N53 = N52 | data_masked[45];
  assign N52 = N51 | data_masked[73];
  assign N51 = data_masked[129] | data_masked[101];
  assign data_o[18] = N56 | data_masked[18];
  assign N56 = N55 | data_masked[46];
  assign N55 = N54 | data_masked[74];
  assign N54 = data_masked[130] | data_masked[102];
  assign data_o[19] = N59 | data_masked[19];
  assign N59 = N58 | data_masked[47];
  assign N58 = N57 | data_masked[75];
  assign N57 = data_masked[131] | data_masked[103];
  assign data_o[20] = N62 | data_masked[20];
  assign N62 = N61 | data_masked[48];
  assign N61 = N60 | data_masked[76];
  assign N60 = data_masked[132] | data_masked[104];
  assign data_o[21] = N65 | data_masked[21];
  assign N65 = N64 | data_masked[49];
  assign N64 = N63 | data_masked[77];
  assign N63 = data_masked[133] | data_masked[105];
  assign data_o[22] = N68 | data_masked[22];
  assign N68 = N67 | data_masked[50];
  assign N67 = N66 | data_masked[78];
  assign N66 = data_masked[134] | data_masked[106];
  assign data_o[23] = N71 | data_masked[23];
  assign N71 = N70 | data_masked[51];
  assign N70 = N69 | data_masked[79];
  assign N69 = data_masked[135] | data_masked[107];
  assign data_o[24] = N74 | data_masked[24];
  assign N74 = N73 | data_masked[52];
  assign N73 = N72 | data_masked[80];
  assign N72 = data_masked[136] | data_masked[108];
  assign data_o[25] = N77 | data_masked[25];
  assign N77 = N76 | data_masked[53];
  assign N76 = N75 | data_masked[81];
  assign N75 = data_masked[137] | data_masked[109];
  assign data_o[26] = N80 | data_masked[26];
  assign N80 = N79 | data_masked[54];
  assign N79 = N78 | data_masked[82];
  assign N78 = data_masked[138] | data_masked[110];
  assign data_o[27] = N83 | data_masked[27];
  assign N83 = N82 | data_masked[55];
  assign N82 = N81 | data_masked[83];
  assign N81 = data_masked[139] | data_masked[111];

endmodule



module bsg_mesh_router_28_1_1_0_0a_0
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  yumi_o,
  ready_i,
  data_o,
  v_o,
  my_x_i,
  my_y_i
);

  input [139:0] data_i;
  input [4:0] v_i;
  output [4:0] yumi_o;
  input [4:0] ready_i;
  output [139:0] data_o;
  output [4:0] v_o;
  input [0:0] my_x_i;
  input [0:0] my_y_i;
  input clk_i;
  input reset_i;
  wire [4:0] yumi_o,v_o;
  wire [139:0] data_o;
  wire n_3_net_,W_sel_e,W_sel_p,W_sel_n,W_sel_s,W_gnt_e,W_gnt_p,W_gnt_n,W_gnt_s,
  n_9_net_,E_sel_w,E_sel_p,E_sel_n,E_sel_s,E_gnt_w,E_gnt_p,E_gnt_n,E_gnt_s,n_15_net_,
  N_sel_s,N_sel_p,N_gnt_s,N_gnt_p,n_21_net_,S_sel_n,S_sel_p,S_gnt_n,S_gnt_p,n_27_net_,
  P_sel_s,P_sel_n,P_sel_e,P_sel_w,P_sel_p,P_gnt_s,P_gnt_n,P_gnt_e,P_gnt_w,P_gnt_p,
  N0,N1,N2,N3,N4,N5,N6,SV2V_UNCONNECTED_1,SV2V_UNCONNECTED_2,
  SV2V_UNCONNECTED_3,SV2V_UNCONNECTED_4,SV2V_UNCONNECTED_5,SV2V_UNCONNECTED_6,
  SV2V_UNCONNECTED_7,SV2V_UNCONNECTED_8,SV2V_UNCONNECTED_9;
  wire [24:0] req;

  bsg_mesh_router_dor_decoder_x_cord_width_p1_y_cord_width_p1_dirs_lp5_XY_order_p0
  dor_decoder
  (
    .clk_i(clk_i),
    .v_i({ v_i[4:4], 1'b0, v_i[2:2], 1'b0, v_i[0:0] }),
    .x_dirs_i({ data_i[112:112], data_i[84:84], data_i[56:56], data_i[28:28], data_i[0:0] }),
    .y_dirs_i({ data_i[113:113], data_i[85:85], data_i[57:57], data_i[29:29], data_i[1:1] }),
    .my_x_i(my_x_i[0]),
    .my_y_i(my_y_i[0]),
    .req_o(req)
  );


  bsg_round_robin_arb_inputs_p4
  genblk2_west_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ req[11:11], req[1:1], req[16:16], req[21:21] }),
    .grants_o({ W_gnt_e, W_gnt_p, W_gnt_n, W_gnt_s }),
    .sel_one_hot_o({ W_sel_e, W_sel_p, W_sel_n, W_sel_s }),
    .v_o(v_o[1]),
    .tag_o({ SV2V_UNCONNECTED_1, SV2V_UNCONNECTED_2 }),
    .yumi_i(n_3_net_)
  );


  bsg_mux_one_hot_width_p28_els_p4
  genblk2_mux_data_west
  (
    .data_i({ data_i[27:0], data_i[83:56], data_i[111:84], data_i[139:112] }),
    .sel_one_hot_i({ W_sel_p, W_sel_e, W_sel_n, W_sel_s }),
    .data_o(data_o[55:28])
  );


  bsg_round_robin_arb_inputs_p4
  genblk3_east_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[2]),
    .reqs_i({ req[7:7], req[2:2], req[17:17], req[22:22] }),
    .grants_o({ E_gnt_w, E_gnt_p, E_gnt_n, E_gnt_s }),
    .sel_one_hot_o({ E_sel_w, E_sel_p, E_sel_n, E_sel_s }),
    .v_o(v_o[2]),
    .tag_o({ SV2V_UNCONNECTED_3, SV2V_UNCONNECTED_4 }),
    .yumi_i(n_9_net_)
  );


  bsg_mux_one_hot_width_p28_els_p4
  genblk3_mux_data_east
  (
    .data_i({ data_i[27:0], data_i[55:28], data_i[111:84], data_i[139:112] }),
    .sel_one_hot_i({ E_sel_p, E_sel_w, E_sel_n, E_sel_s }),
    .data_o(data_o[83:56])
  );


  bsg_round_robin_arb_inputs_p2
  genblk4_north_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ req[23:23], req[3:3] }),
    .grants_o({ N_gnt_s, N_gnt_p }),
    .sel_one_hot_o({ N_sel_s, N_sel_p }),
    .v_o(v_o[3]),
    .tag_o(SV2V_UNCONNECTED_5),
    .yumi_i(n_15_net_)
  );


  bsg_mux_one_hot_width_p28_els_p2
  genblk4_mux_data_north
  (
    .data_i({ data_i[27:0], data_i[139:112] }),
    .sel_one_hot_i({ N_sel_p, N_sel_s }),
    .data_o(data_o[111:84])
  );


  bsg_round_robin_arb_inputs_p2
  genblk5_south_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[4]),
    .reqs_i({ req[19:19], req[4:4] }),
    .grants_o({ S_gnt_n, S_gnt_p }),
    .sel_one_hot_o({ S_sel_n, S_sel_p }),
    .v_o(v_o[4]),
    .tag_o(SV2V_UNCONNECTED_6),
    .yumi_i(n_21_net_)
  );


  bsg_mux_one_hot_width_p28_els_p2
  genblk5_mux_data_south
  (
    .data_i({ data_i[27:0], data_i[111:84] }),
    .sel_one_hot_i({ S_sel_p, S_sel_n }),
    .data_o(data_o[139:112])
  );


  bsg_round_robin_arb_inputs_p5
  proc_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[0]),
    .reqs_i({ req[20:20], req[15:15], req[10:10], req[5:5], req[0:0] }),
    .grants_o({ P_gnt_s, P_gnt_n, P_gnt_e, P_gnt_w, P_gnt_p }),
    .sel_one_hot_o({ P_sel_s, P_sel_n, P_sel_e, P_sel_w, P_sel_p }),
    .v_o(v_o[0]),
    .tag_o({ SV2V_UNCONNECTED_7, SV2V_UNCONNECTED_8, SV2V_UNCONNECTED_9 }),
    .yumi_i(n_27_net_)
  );


  bsg_mux_one_hot_width_p28_els_p5
  mux_data_proc
  (
    .data_i({ data_i[27:0], data_i[83:56], data_i[139:112], data_i[55:28], data_i[111:84] }),
    .sel_one_hot_i({ P_sel_p, P_sel_e, P_sel_s, P_sel_w, P_sel_n }),
    .data_o(data_o[27:0])
  );

  assign n_3_net_ = v_o[1] & 1'b1;
  assign n_9_net_ = v_o[2] & ready_i[2];
  assign n_15_net_ = v_o[3] & 1'b1;
  assign n_21_net_ = v_o[4] & ready_i[4];
  assign n_27_net_ = v_o[0] & ready_i[0];
  assign yumi_o[0] = N2 | W_gnt_p;
  assign N2 = N1 | P_gnt_p;
  assign N1 = N0 | S_gnt_p;
  assign N0 = E_gnt_p | N_gnt_p;
  assign yumi_o[1] = E_gnt_w | P_gnt_w;
  assign yumi_o[2] = W_gnt_e | P_gnt_e;
  assign yumi_o[3] = N4 | P_gnt_n;
  assign N4 = N3 | E_gnt_n;
  assign N3 = S_gnt_n | W_gnt_n;
  assign yumi_o[4] = N6 | P_gnt_s;
  assign N6 = N5 | E_gnt_s;
  assign N5 = N_gnt_s | W_gnt_s;

endmodule



module bsg_mesh_router_buffered_28_1_1_0_5_0a_0_30_00
(
  clk_i,
  reset_i,
  link_i,
  link_o,
  my_x_i,
  my_y_i
);

  input [149:0] link_i;
  output [149:0] link_o;
  input [0:0] my_x_i;
  input [0:0] my_y_i;
  input clk_i;
  input reset_i;
  wire [149:0] link_o;
  wire fifo_valid_2,fifo_valid_0,fifo_data_4__27_,fifo_data_4__26_,fifo_data_4__25_,
  fifo_data_4__24_,fifo_data_4__23_,fifo_data_4__22_,fifo_data_4__21_,
  fifo_data_4__20_,fifo_data_4__19_,fifo_data_4__18_,fifo_data_4__17_,fifo_data_4__16_,
  fifo_data_4__15_,fifo_data_4__14_,fifo_data_4__13_,fifo_data_4__12_,fifo_data_4__11_,
  fifo_data_4__10_,fifo_data_4__9_,fifo_data_4__8_,fifo_data_4__7_,fifo_data_4__6_,
  fifo_data_4__5_,fifo_data_4__4_,fifo_data_4__3_,fifo_data_4__2_,fifo_data_4__1_,
  fifo_data_4__0_,fifo_data_2__27_,fifo_data_2__26_,fifo_data_2__25_,fifo_data_2__24_,
  fifo_data_2__23_,fifo_data_2__22_,fifo_data_2__21_,fifo_data_2__20_,
  fifo_data_2__19_,fifo_data_2__18_,fifo_data_2__17_,fifo_data_2__16_,fifo_data_2__15_,
  fifo_data_2__14_,fifo_data_2__13_,fifo_data_2__12_,fifo_data_2__11_,fifo_data_2__10_,
  fifo_data_2__9_,fifo_data_2__8_,fifo_data_2__7_,fifo_data_2__6_,fifo_data_2__5_,
  fifo_data_2__4_,fifo_data_2__3_,fifo_data_2__2_,fifo_data_2__1_,fifo_data_2__0_,
  fifo_data_0__27_,fifo_data_0__26_,fifo_data_0__25_,fifo_data_0__24_,
  fifo_data_0__23_,fifo_data_0__22_,fifo_data_0__21_,fifo_data_0__20_,fifo_data_0__19_,
  fifo_data_0__18_,fifo_data_0__17_,fifo_data_0__16_,fifo_data_0__15_,fifo_data_0__14_,
  fifo_data_0__13_,fifo_data_0__12_,fifo_data_0__11_,fifo_data_0__10_,fifo_data_0__9_,
  fifo_data_0__8_,fifo_data_0__7_,fifo_data_0__6_,fifo_data_0__5_,fifo_data_0__4_,
  fifo_data_0__3_,fifo_data_0__2_,fifo_data_0__1_,fifo_data_0__0_;
  wire [4:4] fifo_valid;
  wire [4:0] fifo_yumi;
  assign link_o[58] = 1'b0;
  assign link_o[118] = 1'b0;

  bsg_two_fifo_width_p28
  rof_0__fi_twofer
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(link_o[28]),
    .data_i(link_i[27:0]),
    .v_i(link_i[29]),
    .v_o(fifo_valid_0),
    .data_o({ fifo_data_0__27_, fifo_data_0__26_, fifo_data_0__25_, fifo_data_0__24_, fifo_data_0__23_, fifo_data_0__22_, fifo_data_0__21_, fifo_data_0__20_, fifo_data_0__19_, fifo_data_0__18_, fifo_data_0__17_, fifo_data_0__16_, fifo_data_0__15_, fifo_data_0__14_, fifo_data_0__13_, fifo_data_0__12_, fifo_data_0__11_, fifo_data_0__10_, fifo_data_0__9_, fifo_data_0__8_, fifo_data_0__7_, fifo_data_0__6_, fifo_data_0__5_, fifo_data_0__4_, fifo_data_0__3_, fifo_data_0__2_, fifo_data_0__1_, fifo_data_0__0_ }),
    .yumi_i(fifo_yumi[0])
  );


  bsg_two_fifo_width_p28
  rof_2__fi_twofer
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(link_o[88]),
    .data_i(link_i[87:60]),
    .v_i(link_i[89]),
    .v_o(fifo_valid_2),
    .data_o({ fifo_data_2__27_, fifo_data_2__26_, fifo_data_2__25_, fifo_data_2__24_, fifo_data_2__23_, fifo_data_2__22_, fifo_data_2__21_, fifo_data_2__20_, fifo_data_2__19_, fifo_data_2__18_, fifo_data_2__17_, fifo_data_2__16_, fifo_data_2__15_, fifo_data_2__14_, fifo_data_2__13_, fifo_data_2__12_, fifo_data_2__11_, fifo_data_2__10_, fifo_data_2__9_, fifo_data_2__8_, fifo_data_2__7_, fifo_data_2__6_, fifo_data_2__5_, fifo_data_2__4_, fifo_data_2__3_, fifo_data_2__2_, fifo_data_2__1_, fifo_data_2__0_ }),
    .yumi_i(fifo_yumi[2])
  );


  bsg_two_fifo_width_p28
  rof_4__fi_twofer
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(link_o[148]),
    .data_i(link_i[147:120]),
    .v_i(link_i[149]),
    .v_o(fifo_valid[4]),
    .data_o({ fifo_data_4__27_, fifo_data_4__26_, fifo_data_4__25_, fifo_data_4__24_, fifo_data_4__23_, fifo_data_4__22_, fifo_data_4__21_, fifo_data_4__20_, fifo_data_4__19_, fifo_data_4__18_, fifo_data_4__17_, fifo_data_4__16_, fifo_data_4__15_, fifo_data_4__14_, fifo_data_4__13_, fifo_data_4__12_, fifo_data_4__11_, fifo_data_4__10_, fifo_data_4__9_, fifo_data_4__8_, fifo_data_4__7_, fifo_data_4__6_, fifo_data_4__5_, fifo_data_4__4_, fifo_data_4__3_, fifo_data_4__2_, fifo_data_4__1_, fifo_data_4__0_ }),
    .yumi_i(fifo_yumi[4])
  );


  bsg_mesh_router_28_1_1_0_0a_0
  bmr
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ fifo_data_4__27_, fifo_data_4__26_, fifo_data_4__25_, fifo_data_4__24_, fifo_data_4__23_, fifo_data_4__22_, fifo_data_4__21_, fifo_data_4__20_, fifo_data_4__19_, fifo_data_4__18_, fifo_data_4__17_, fifo_data_4__16_, fifo_data_4__15_, fifo_data_4__14_, fifo_data_4__13_, fifo_data_4__12_, fifo_data_4__11_, fifo_data_4__10_, fifo_data_4__9_, fifo_data_4__8_, fifo_data_4__7_, fifo_data_4__6_, fifo_data_4__5_, fifo_data_4__4_, fifo_data_4__3_, fifo_data_4__2_, fifo_data_4__1_, fifo_data_4__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_2__27_, fifo_data_2__26_, fifo_data_2__25_, fifo_data_2__24_, fifo_data_2__23_, fifo_data_2__22_, fifo_data_2__21_, fifo_data_2__20_, fifo_data_2__19_, fifo_data_2__18_, fifo_data_2__17_, fifo_data_2__16_, fifo_data_2__15_, fifo_data_2__14_, fifo_data_2__13_, fifo_data_2__12_, fifo_data_2__11_, fifo_data_2__10_, fifo_data_2__9_, fifo_data_2__8_, fifo_data_2__7_, fifo_data_2__6_, fifo_data_2__5_, fifo_data_2__4_, fifo_data_2__3_, fifo_data_2__2_, fifo_data_2__1_, fifo_data_2__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_0__27_, fifo_data_0__26_, fifo_data_0__25_, fifo_data_0__24_, fifo_data_0__23_, fifo_data_0__22_, fifo_data_0__21_, fifo_data_0__20_, fifo_data_0__19_, fifo_data_0__18_, fifo_data_0__17_, fifo_data_0__16_, fifo_data_0__15_, fifo_data_0__14_, fifo_data_0__13_, fifo_data_0__12_, fifo_data_0__11_, fifo_data_0__10_, fifo_data_0__9_, fifo_data_0__8_, fifo_data_0__7_, fifo_data_0__6_, fifo_data_0__5_, fifo_data_0__4_, fifo_data_0__3_, fifo_data_0__2_, fifo_data_0__1_, fifo_data_0__0_ }),
    .v_i({ fifo_valid[4:4], 1'b0, fifo_valid_2, 1'b0, fifo_valid_0 }),
    .yumi_o(fifo_yumi),
    .ready_i({ link_i[148:148], link_i[118:118], link_i[88:88], link_i[58:58], link_i[28:28] }),
    .data_o({ link_o[147:120], link_o[117:90], link_o[87:60], link_o[57:30], link_o[27:0] }),
    .v_o({ link_o[149:149], link_o[119:119], link_o[89:89], link_o[59:59], link_o[29:29] }),
    .my_x_i(my_x_i[0]),
    .my_y_i(my_y_i[0])
  );


endmodule



module bsg_mesh_router_28_1_1_0_0d_0
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  yumi_o,
  ready_i,
  data_o,
  v_o,
  my_x_i,
  my_y_i
);

  input [139:0] data_i;
  input [4:0] v_i;
  output [4:0] yumi_o;
  input [4:0] ready_i;
  output [139:0] data_o;
  output [4:0] v_o;
  input [0:0] my_x_i;
  input [0:0] my_y_i;
  input clk_i;
  input reset_i;
  wire [4:0] yumi_o,v_o;
  wire [139:0] data_o;
  wire n_3_net_,W_sel_e,W_sel_p,W_sel_n,W_sel_s,W_gnt_e,W_gnt_p,W_gnt_n,W_gnt_s,
  n_9_net_,E_sel_w,E_sel_p,E_sel_n,E_sel_s,E_gnt_w,E_gnt_p,E_gnt_n,E_gnt_s,n_15_net_,
  N_sel_s,N_sel_p,N_gnt_s,N_gnt_p,n_21_net_,S_sel_n,S_sel_p,S_gnt_n,S_gnt_p,n_27_net_,
  P_sel_s,P_sel_n,P_sel_e,P_sel_w,P_sel_p,P_gnt_s,P_gnt_n,P_gnt_e,P_gnt_w,P_gnt_p,
  N0,N1,N2,N3,N4,N5,N6,SV2V_UNCONNECTED_1,SV2V_UNCONNECTED_2,
  SV2V_UNCONNECTED_3,SV2V_UNCONNECTED_4,SV2V_UNCONNECTED_5,SV2V_UNCONNECTED_6,
  SV2V_UNCONNECTED_7,SV2V_UNCONNECTED_8,SV2V_UNCONNECTED_9;
  wire [24:0] req;

  bsg_mesh_router_dor_decoder_x_cord_width_p1_y_cord_width_p1_dirs_lp5_XY_order_p0
  dor_decoder
  (
    .clk_i(clk_i),
    .v_i({ v_i[4:4], 1'b0, 1'b0, v_i[1:1], 1'b0 }),
    .x_dirs_i({ data_i[112:112], data_i[84:84], data_i[56:56], data_i[28:28], data_i[0:0] }),
    .y_dirs_i({ data_i[113:113], data_i[85:85], data_i[57:57], data_i[29:29], data_i[1:1] }),
    .my_x_i(my_x_i[0]),
    .my_y_i(my_y_i[0]),
    .req_o(req)
  );


  bsg_round_robin_arb_inputs_p4
  genblk2_west_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[1]),
    .reqs_i({ req[11:11], req[1:1], req[16:16], req[21:21] }),
    .grants_o({ W_gnt_e, W_gnt_p, W_gnt_n, W_gnt_s }),
    .sel_one_hot_o({ W_sel_e, W_sel_p, W_sel_n, W_sel_s }),
    .v_o(v_o[1]),
    .tag_o({ SV2V_UNCONNECTED_1, SV2V_UNCONNECTED_2 }),
    .yumi_i(n_3_net_)
  );


  bsg_mux_one_hot_width_p28_els_p4
  genblk2_mux_data_west
  (
    .data_i({ data_i[27:0], data_i[83:56], data_i[111:84], data_i[139:112] }),
    .sel_one_hot_i({ W_sel_p, W_sel_e, W_sel_n, W_sel_s }),
    .data_o(data_o[55:28])
  );


  bsg_round_robin_arb_inputs_p4
  genblk3_east_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ req[7:7], req[2:2], req[17:17], req[22:22] }),
    .grants_o({ E_gnt_w, E_gnt_p, E_gnt_n, E_gnt_s }),
    .sel_one_hot_o({ E_sel_w, E_sel_p, E_sel_n, E_sel_s }),
    .v_o(v_o[2]),
    .tag_o({ SV2V_UNCONNECTED_3, SV2V_UNCONNECTED_4 }),
    .yumi_i(n_9_net_)
  );


  bsg_mux_one_hot_width_p28_els_p4
  genblk3_mux_data_east
  (
    .data_i({ data_i[27:0], data_i[55:28], data_i[111:84], data_i[139:112] }),
    .sel_one_hot_i({ E_sel_p, E_sel_w, E_sel_n, E_sel_s }),
    .data_o(data_o[83:56])
  );


  bsg_round_robin_arb_inputs_p2
  genblk4_north_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ req[23:23], req[3:3] }),
    .grants_o({ N_gnt_s, N_gnt_p }),
    .sel_one_hot_o({ N_sel_s, N_sel_p }),
    .v_o(v_o[3]),
    .tag_o(SV2V_UNCONNECTED_5),
    .yumi_i(n_15_net_)
  );


  bsg_mux_one_hot_width_p28_els_p2
  genblk4_mux_data_north
  (
    .data_i({ data_i[27:0], data_i[139:112] }),
    .sel_one_hot_i({ N_sel_p, N_sel_s }),
    .data_o(data_o[111:84])
  );


  bsg_round_robin_arb_inputs_p2
  genblk5_south_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[4]),
    .reqs_i({ req[19:19], req[4:4] }),
    .grants_o({ S_gnt_n, S_gnt_p }),
    .sel_one_hot_o({ S_sel_n, S_sel_p }),
    .v_o(v_o[4]),
    .tag_o(SV2V_UNCONNECTED_6),
    .yumi_i(n_21_net_)
  );


  bsg_mux_one_hot_width_p28_els_p2
  genblk5_mux_data_south
  (
    .data_i({ data_i[27:0], data_i[111:84] }),
    .sel_one_hot_i({ S_sel_p, S_sel_n }),
    .data_o(data_o[139:112])
  );


  bsg_round_robin_arb_inputs_p5
  proc_rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ req[20:20], req[15:15], req[10:10], req[5:5], req[0:0] }),
    .grants_o({ P_gnt_s, P_gnt_n, P_gnt_e, P_gnt_w, P_gnt_p }),
    .sel_one_hot_o({ P_sel_s, P_sel_n, P_sel_e, P_sel_w, P_sel_p }),
    .v_o(v_o[0]),
    .tag_o({ SV2V_UNCONNECTED_7, SV2V_UNCONNECTED_8, SV2V_UNCONNECTED_9 }),
    .yumi_i(n_27_net_)
  );


  bsg_mux_one_hot_width_p28_els_p5
  mux_data_proc
  (
    .data_i({ data_i[27:0], data_i[83:56], data_i[139:112], data_i[55:28], data_i[111:84] }),
    .sel_one_hot_i({ P_sel_p, P_sel_e, P_sel_s, P_sel_w, P_sel_n }),
    .data_o(data_o[27:0])
  );

  assign n_3_net_ = v_o[1] & ready_i[1];
  assign n_9_net_ = v_o[2] & 1'b1;
  assign n_15_net_ = v_o[3] & 1'b1;
  assign n_21_net_ = v_o[4] & ready_i[4];
  assign n_27_net_ = v_o[0] & 1'b1;
  assign yumi_o[0] = N2 | W_gnt_p;
  assign N2 = N1 | P_gnt_p;
  assign N1 = N0 | S_gnt_p;
  assign N0 = E_gnt_p | N_gnt_p;
  assign yumi_o[1] = E_gnt_w | P_gnt_w;
  assign yumi_o[2] = W_gnt_e | P_gnt_e;
  assign yumi_o[3] = N4 | P_gnt_n;
  assign N4 = N3 | E_gnt_n;
  assign N3 = S_gnt_n | W_gnt_n;
  assign yumi_o[4] = N6 | P_gnt_s;
  assign N6 = N5 | E_gnt_s;
  assign N5 = N_gnt_s | W_gnt_s;

endmodule



module bsg_mesh_router_buffered_28_1_1_0_5_0d_0_30_00
(
  clk_i,
  reset_i,
  link_i,
  link_o,
  my_x_i,
  my_y_i
);

  input [149:0] link_i;
  output [149:0] link_o;
  input [0:0] my_x_i;
  input [0:0] my_y_i;
  input clk_i;
  input reset_i;
  wire [149:0] link_o;
  wire fifo_data_4__27_,fifo_data_4__26_,fifo_data_4__25_,fifo_data_4__24_,
  fifo_data_4__23_,fifo_data_4__22_,fifo_data_4__21_,fifo_data_4__20_,fifo_data_4__19_,
  fifo_data_4__18_,fifo_data_4__17_,fifo_data_4__16_,fifo_data_4__15_,fifo_data_4__14_,
  fifo_data_4__13_,fifo_data_4__12_,fifo_data_4__11_,fifo_data_4__10_,
  fifo_data_4__9_,fifo_data_4__8_,fifo_data_4__7_,fifo_data_4__6_,fifo_data_4__5_,
  fifo_data_4__4_,fifo_data_4__3_,fifo_data_4__2_,fifo_data_4__1_,fifo_data_4__0_,
  fifo_data_1__27_,fifo_data_1__26_,fifo_data_1__25_,fifo_data_1__24_,fifo_data_1__23_,
  fifo_data_1__22_,fifo_data_1__21_,fifo_data_1__20_,fifo_data_1__19_,fifo_data_1__18_,
  fifo_data_1__17_,fifo_data_1__16_,fifo_data_1__15_,fifo_data_1__14_,
  fifo_data_1__13_,fifo_data_1__12_,fifo_data_1__11_,fifo_data_1__10_,fifo_data_1__9_,
  fifo_data_1__8_,fifo_data_1__7_,fifo_data_1__6_,fifo_data_1__5_,fifo_data_1__4_,
  fifo_data_1__3_,fifo_data_1__2_,fifo_data_1__1_,fifo_data_1__0_,fifo_valid_1;
  wire [4:4] fifo_valid;
  wire [4:0] fifo_yumi;
  assign link_o[28] = 1'b0;
  assign link_o[88] = 1'b0;
  assign link_o[118] = 1'b0;

  bsg_two_fifo_width_p28
  rof_1__fi_twofer
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(link_o[58]),
    .data_i(link_i[57:30]),
    .v_i(link_i[59]),
    .v_o(fifo_valid_1),
    .data_o({ fifo_data_1__27_, fifo_data_1__26_, fifo_data_1__25_, fifo_data_1__24_, fifo_data_1__23_, fifo_data_1__22_, fifo_data_1__21_, fifo_data_1__20_, fifo_data_1__19_, fifo_data_1__18_, fifo_data_1__17_, fifo_data_1__16_, fifo_data_1__15_, fifo_data_1__14_, fifo_data_1__13_, fifo_data_1__12_, fifo_data_1__11_, fifo_data_1__10_, fifo_data_1__9_, fifo_data_1__8_, fifo_data_1__7_, fifo_data_1__6_, fifo_data_1__5_, fifo_data_1__4_, fifo_data_1__3_, fifo_data_1__2_, fifo_data_1__1_, fifo_data_1__0_ }),
    .yumi_i(fifo_yumi[1])
  );


  bsg_two_fifo_width_p28
  rof_4__fi_twofer
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(link_o[148]),
    .data_i(link_i[147:120]),
    .v_i(link_i[149]),
    .v_o(fifo_valid[4]),
    .data_o({ fifo_data_4__27_, fifo_data_4__26_, fifo_data_4__25_, fifo_data_4__24_, fifo_data_4__23_, fifo_data_4__22_, fifo_data_4__21_, fifo_data_4__20_, fifo_data_4__19_, fifo_data_4__18_, fifo_data_4__17_, fifo_data_4__16_, fifo_data_4__15_, fifo_data_4__14_, fifo_data_4__13_, fifo_data_4__12_, fifo_data_4__11_, fifo_data_4__10_, fifo_data_4__9_, fifo_data_4__8_, fifo_data_4__7_, fifo_data_4__6_, fifo_data_4__5_, fifo_data_4__4_, fifo_data_4__3_, fifo_data_4__2_, fifo_data_4__1_, fifo_data_4__0_ }),
    .yumi_i(fifo_yumi[4])
  );


  bsg_mesh_router_28_1_1_0_0d_0
  bmr
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i({ fifo_data_4__27_, fifo_data_4__26_, fifo_data_4__25_, fifo_data_4__24_, fifo_data_4__23_, fifo_data_4__22_, fifo_data_4__21_, fifo_data_4__20_, fifo_data_4__19_, fifo_data_4__18_, fifo_data_4__17_, fifo_data_4__16_, fifo_data_4__15_, fifo_data_4__14_, fifo_data_4__13_, fifo_data_4__12_, fifo_data_4__11_, fifo_data_4__10_, fifo_data_4__9_, fifo_data_4__8_, fifo_data_4__7_, fifo_data_4__6_, fifo_data_4__5_, fifo_data_4__4_, fifo_data_4__3_, fifo_data_4__2_, fifo_data_4__1_, fifo_data_4__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_1__27_, fifo_data_1__26_, fifo_data_1__25_, fifo_data_1__24_, fifo_data_1__23_, fifo_data_1__22_, fifo_data_1__21_, fifo_data_1__20_, fifo_data_1__19_, fifo_data_1__18_, fifo_data_1__17_, fifo_data_1__16_, fifo_data_1__15_, fifo_data_1__14_, fifo_data_1__13_, fifo_data_1__12_, fifo_data_1__11_, fifo_data_1__10_, fifo_data_1__9_, fifo_data_1__8_, fifo_data_1__7_, fifo_data_1__6_, fifo_data_1__5_, fifo_data_1__4_, fifo_data_1__3_, fifo_data_1__2_, fifo_data_1__1_, fifo_data_1__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .v_i({ fifo_valid[4:4], 1'b0, 1'b0, fifo_valid_1, 1'b0 }),
    .yumi_o(fifo_yumi),
    .ready_i({ link_i[148:148], link_i[118:118], link_i[88:88], link_i[58:58], link_i[28:28] }),
    .data_o({ link_o[147:120], link_o[117:90], link_o[87:60], link_o[57:30], link_o[27:0] }),
    .v_o({ link_o[149:149], link_o[119:119], link_o[89:89], link_o[59:59], link_o[29:29] }),
    .my_x_i(my_x_i[0]),
    .my_y_i(my_y_i[0])
  );


endmodule



module bp_me_network_channel_mesh_packet_width_p26_num_src_p2_num_dst_p1_debug_p0
(
  clk_i,
  reset_i,
  src_data_i,
  src_v_i,
  src_ready_o,
  dst_data_o,
  dst_v_o,
  dst_ready_i
);

  input [51:0] src_data_i;
  input [1:0] src_v_i;
  output [1:0] src_ready_o;
  output [25:0] dst_data_o;
  output [0:0] dst_v_o;
  input [0:0] dst_ready_i;
  input clk_i;
  input reset_i;
  wire [1:0] src_ready_o;
  wire [25:0] dst_data_o;
  wire [0:0] dst_v_o;
  wire link_i_stitch_0__2__v_,link_i_stitch_0__2__ready_then_rev_,
  link_i_stitch_0__2__data__27_,link_i_stitch_0__2__data__26_,link_i_stitch_0__2__data__25_,
  link_i_stitch_0__2__data__24_,link_i_stitch_0__2__data__23_,link_i_stitch_0__2__data__22_,
  link_i_stitch_0__2__data__21_,link_i_stitch_0__2__data__20_,
  link_i_stitch_0__2__data__19_,link_i_stitch_0__2__data__18_,link_i_stitch_0__2__data__17_,
  link_i_stitch_0__2__data__16_,link_i_stitch_0__2__data__15_,link_i_stitch_0__2__data__14_,
  link_i_stitch_0__2__data__13_,link_i_stitch_0__2__data__12_,
  link_i_stitch_0__2__data__11_,link_i_stitch_0__2__data__10_,link_i_stitch_0__2__data__9_,
  link_i_stitch_0__2__data__8_,link_i_stitch_0__2__data__7_,link_i_stitch_0__2__data__6_,
  link_i_stitch_0__2__data__5_,link_i_stitch_0__2__data__4_,
  link_i_stitch_0__2__data__3_,link_i_stitch_0__2__data__2_,link_i_stitch_0__2__data__1_,
  link_i_stitch_0__2__data__0_,link_o_stitch_1__4__v_,link_o_stitch_1__4__data__27_,
  link_o_stitch_1__4__data__26_,link_o_stitch_1__4__data__25_,link_o_stitch_1__4__data__24_,
  link_o_stitch_1__4__data__23_,link_o_stitch_1__4__data__22_,
  link_o_stitch_1__4__data__21_,link_o_stitch_1__4__data__20_,link_o_stitch_1__4__data__19_,
  link_o_stitch_1__4__data__18_,link_o_stitch_1__4__data__17_,link_o_stitch_1__4__data__16_,
  link_o_stitch_1__4__data__15_,link_o_stitch_1__4__data__14_,
  link_o_stitch_1__4__data__13_,link_o_stitch_1__4__data__12_,link_o_stitch_1__4__data__11_,
  link_o_stitch_1__4__data__10_,link_o_stitch_1__4__data__9_,link_o_stitch_1__4__data__8_,
  link_o_stitch_1__4__data__7_,link_o_stitch_1__4__data__6_,link_o_stitch_1__4__data__5_,
  link_o_stitch_1__4__data__4_,link_o_stitch_1__4__data__3_,
  link_o_stitch_1__4__data__2_,link_o_stitch_1__4__data__1_,link_o_stitch_1__4__data__0_,
  link_o_stitch_1__3__v_,link_o_stitch_1__3__ready_then_rev_,link_o_stitch_1__3__data__27_,
  link_o_stitch_1__3__data__26_,link_o_stitch_1__3__data__25_,
  link_o_stitch_1__3__data__24_,link_o_stitch_1__3__data__23_,link_o_stitch_1__3__data__22_,
  link_o_stitch_1__3__data__21_,link_o_stitch_1__3__data__20_,link_o_stitch_1__3__data__19_,
  link_o_stitch_1__3__data__18_,link_o_stitch_1__3__data__17_,
  link_o_stitch_1__3__data__16_,link_o_stitch_1__3__data__15_,link_o_stitch_1__3__data__14_,
  link_o_stitch_1__3__data__13_,link_o_stitch_1__3__data__12_,link_o_stitch_1__3__data__11_,
  link_o_stitch_1__3__data__10_,link_o_stitch_1__3__data__9_,link_o_stitch_1__3__data__8_,
  link_o_stitch_1__3__data__7_,link_o_stitch_1__3__data__6_,
  link_o_stitch_1__3__data__5_,link_o_stitch_1__3__data__4_,link_o_stitch_1__3__data__3_,
  link_o_stitch_1__3__data__2_,link_o_stitch_1__3__data__1_,link_o_stitch_1__3__data__0_,
  link_o_stitch_1__2__v_,link_o_stitch_1__2__ready_then_rev_,link_o_stitch_1__2__data__27_,
  link_o_stitch_1__2__data__26_,link_o_stitch_1__2__data__25_,
  link_o_stitch_1__2__data__24_,link_o_stitch_1__2__data__23_,link_o_stitch_1__2__data__22_,
  link_o_stitch_1__2__data__21_,link_o_stitch_1__2__data__20_,link_o_stitch_1__2__data__19_,
  link_o_stitch_1__2__data__18_,link_o_stitch_1__2__data__17_,
  link_o_stitch_1__2__data__16_,link_o_stitch_1__2__data__15_,link_o_stitch_1__2__data__14_,
  link_o_stitch_1__2__data__13_,link_o_stitch_1__2__data__12_,link_o_stitch_1__2__data__11_,
  link_o_stitch_1__2__data__10_,link_o_stitch_1__2__data__9_,
  link_o_stitch_1__2__data__8_,link_o_stitch_1__2__data__7_,link_o_stitch_1__2__data__6_,
  link_o_stitch_1__2__data__5_,link_o_stitch_1__2__data__4_,link_o_stitch_1__2__data__3_,
  link_o_stitch_1__2__data__2_,link_o_stitch_1__2__data__1_,link_o_stitch_1__2__data__0_,
  link_o_stitch_1__0__v_,link_o_stitch_1__0__ready_then_rev_,
  link_o_stitch_1__0__data__27_,link_o_stitch_1__0__data__26_,link_o_stitch_1__0__data__25_,
  link_o_stitch_1__0__data__24_,link_o_stitch_1__0__data__23_,link_o_stitch_1__0__data__22_,
  link_o_stitch_1__0__data__21_,link_o_stitch_1__0__data__20_,
  link_o_stitch_1__0__data__19_,link_o_stitch_1__0__data__18_,link_o_stitch_1__0__data__17_,
  link_o_stitch_1__0__data__16_,link_o_stitch_1__0__data__15_,link_o_stitch_1__0__data__14_,
  link_o_stitch_1__0__data__13_,link_o_stitch_1__0__data__12_,
  link_o_stitch_1__0__data__11_,link_o_stitch_1__0__data__10_,link_o_stitch_1__0__data__9_,
  link_o_stitch_1__0__data__8_,link_o_stitch_1__0__data__7_,link_o_stitch_1__0__data__6_,
  link_o_stitch_1__0__data__5_,link_o_stitch_1__0__data__4_,
  link_o_stitch_1__0__data__3_,link_o_stitch_1__0__data__2_,link_o_stitch_1__0__data__1_,
  link_o_stitch_1__0__data__0_,link_o_stitch_0__4__v_,link_o_stitch_0__4__data__27_,
  link_o_stitch_0__4__data__26_,link_o_stitch_0__4__data__25_,link_o_stitch_0__4__data__24_,
  link_o_stitch_0__4__data__23_,link_o_stitch_0__4__data__22_,
  link_o_stitch_0__4__data__21_,link_o_stitch_0__4__data__20_,link_o_stitch_0__4__data__19_,
  link_o_stitch_0__4__data__18_,link_o_stitch_0__4__data__17_,link_o_stitch_0__4__data__16_,
  link_o_stitch_0__4__data__15_,link_o_stitch_0__4__data__14_,
  link_o_stitch_0__4__data__13_,link_o_stitch_0__4__data__12_,link_o_stitch_0__4__data__11_,
  link_o_stitch_0__4__data__10_,link_o_stitch_0__4__data__9_,link_o_stitch_0__4__data__8_,
  link_o_stitch_0__4__data__7_,link_o_stitch_0__4__data__6_,link_o_stitch_0__4__data__5_,
  link_o_stitch_0__4__data__4_,link_o_stitch_0__4__data__3_,
  link_o_stitch_0__4__data__2_,link_o_stitch_0__4__data__1_,link_o_stitch_0__4__data__0_,
  link_o_stitch_0__3__v_,link_o_stitch_0__3__ready_then_rev_,link_o_stitch_0__3__data__27_,
  link_o_stitch_0__3__data__26_,link_o_stitch_0__3__data__25_,
  link_o_stitch_0__3__data__24_,link_o_stitch_0__3__data__23_,link_o_stitch_0__3__data__22_,
  link_o_stitch_0__3__data__21_,link_o_stitch_0__3__data__20_,link_o_stitch_0__3__data__19_,
  link_o_stitch_0__3__data__18_,link_o_stitch_0__3__data__17_,
  link_o_stitch_0__3__data__16_,link_o_stitch_0__3__data__15_,link_o_stitch_0__3__data__14_,
  link_o_stitch_0__3__data__13_,link_o_stitch_0__3__data__12_,link_o_stitch_0__3__data__11_,
  link_o_stitch_0__3__data__10_,link_o_stitch_0__3__data__9_,link_o_stitch_0__3__data__8_,
  link_o_stitch_0__3__data__7_,link_o_stitch_0__3__data__6_,
  link_o_stitch_0__3__data__5_,link_o_stitch_0__3__data__4_,link_o_stitch_0__3__data__3_,
  link_o_stitch_0__3__data__2_,link_o_stitch_0__3__data__1_,link_o_stitch_0__3__data__0_,
  link_o_stitch_0__2__v_,link_o_stitch_0__2__ready_then_rev_,link_o_stitch_0__2__data__27_,
  link_o_stitch_0__2__data__26_,link_o_stitch_0__2__data__25_,
  link_o_stitch_0__2__data__24_,link_o_stitch_0__2__data__23_,link_o_stitch_0__2__data__22_,
  link_o_stitch_0__2__data__21_,link_o_stitch_0__2__data__20_,link_o_stitch_0__2__data__19_,
  link_o_stitch_0__2__data__18_,link_o_stitch_0__2__data__17_,
  link_o_stitch_0__2__data__16_,link_o_stitch_0__2__data__15_,link_o_stitch_0__2__data__14_,
  link_o_stitch_0__2__data__13_,link_o_stitch_0__2__data__12_,link_o_stitch_0__2__data__11_,
  link_o_stitch_0__2__data__10_,link_o_stitch_0__2__data__9_,
  link_o_stitch_0__2__data__8_,link_o_stitch_0__2__data__7_,link_o_stitch_0__2__data__6_,
  link_o_stitch_0__2__data__5_,link_o_stitch_0__2__data__4_,link_o_stitch_0__2__data__3_,
  link_o_stitch_0__2__data__2_,link_o_stitch_0__2__data__1_,link_o_stitch_0__2__data__0_,
  link_o_stitch_0__1__v_,link_o_stitch_0__1__ready_then_rev_,
  link_o_stitch_0__1__data__27_,link_o_stitch_0__1__data__26_,link_o_stitch_0__1__data__25_,
  link_o_stitch_0__1__data__24_,link_o_stitch_0__1__data__23_,link_o_stitch_0__1__data__22_,
  link_o_stitch_0__1__data__21_,link_o_stitch_0__1__data__20_,
  link_o_stitch_0__1__data__19_,link_o_stitch_0__1__data__18_,link_o_stitch_0__1__data__17_,
  link_o_stitch_0__1__data__16_,link_o_stitch_0__1__data__15_,link_o_stitch_0__1__data__14_,
  link_o_stitch_0__1__data__13_,link_o_stitch_0__1__data__12_,
  link_o_stitch_0__1__data__11_,link_o_stitch_0__1__data__10_,link_o_stitch_0__1__data__9_,
  link_o_stitch_0__1__data__8_,link_o_stitch_0__1__data__7_,link_o_stitch_0__1__data__6_,
  link_o_stitch_0__1__data__5_,link_o_stitch_0__1__data__4_,
  link_o_stitch_0__1__data__3_,link_o_stitch_0__1__data__2_,link_o_stitch_0__1__data__1_,
  link_o_stitch_0__1__data__0_,link_o_stitch_0__0__ready_then_rev_,link_o_stitch_0__0__data__1_,
  link_o_stitch_0__0__data__0_;

  bsg_mesh_router_buffered_28_1_1_0_5_0a_0_30_00
  rof_0__fi2_efi3_coherence_network_channel_node
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .link_i({ src_v_i[0:0], 1'b0, src_data_i[25:0], 1'b1, src_data_i[25:25], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, link_i_stitch_0__2__v_, link_i_stitch_0__2__ready_then_rev_, link_i_stitch_0__2__data__27_, link_i_stitch_0__2__data__26_, link_i_stitch_0__2__data__25_, link_i_stitch_0__2__data__24_, link_i_stitch_0__2__data__23_, link_i_stitch_0__2__data__22_, link_i_stitch_0__2__data__21_, link_i_stitch_0__2__data__20_, link_i_stitch_0__2__data__19_, link_i_stitch_0__2__data__18_, link_i_stitch_0__2__data__17_, link_i_stitch_0__2__data__16_, link_i_stitch_0__2__data__15_, link_i_stitch_0__2__data__14_, link_i_stitch_0__2__data__13_, link_i_stitch_0__2__data__12_, link_i_stitch_0__2__data__11_, link_i_stitch_0__2__data__10_, link_i_stitch_0__2__data__9_, link_i_stitch_0__2__data__8_, link_i_stitch_0__2__data__7_, link_i_stitch_0__2__data__6_, link_i_stitch_0__2__data__5_, link_i_stitch_0__2__data__4_, link_i_stitch_0__2__data__3_, link_i_stitch_0__2__data__2_, link_i_stitch_0__2__data__1_, link_i_stitch_0__2__data__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, dst_ready_i[0:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .link_o({ link_o_stitch_0__4__v_, src_ready_o[0:0], link_o_stitch_0__4__data__27_, link_o_stitch_0__4__data__26_, link_o_stitch_0__4__data__25_, link_o_stitch_0__4__data__24_, link_o_stitch_0__4__data__23_, link_o_stitch_0__4__data__22_, link_o_stitch_0__4__data__21_, link_o_stitch_0__4__data__20_, link_o_stitch_0__4__data__19_, link_o_stitch_0__4__data__18_, link_o_stitch_0__4__data__17_, link_o_stitch_0__4__data__16_, link_o_stitch_0__4__data__15_, link_o_stitch_0__4__data__14_, link_o_stitch_0__4__data__13_, link_o_stitch_0__4__data__12_, link_o_stitch_0__4__data__11_, link_o_stitch_0__4__data__10_, link_o_stitch_0__4__data__9_, link_o_stitch_0__4__data__8_, link_o_stitch_0__4__data__7_, link_o_stitch_0__4__data__6_, link_o_stitch_0__4__data__5_, link_o_stitch_0__4__data__4_, link_o_stitch_0__4__data__3_, link_o_stitch_0__4__data__2_, link_o_stitch_0__4__data__1_, link_o_stitch_0__4__data__0_, link_o_stitch_0__3__v_, link_o_stitch_0__3__ready_then_rev_, link_o_stitch_0__3__data__27_, link_o_stitch_0__3__data__26_, link_o_stitch_0__3__data__25_, link_o_stitch_0__3__data__24_, link_o_stitch_0__3__data__23_, link_o_stitch_0__3__data__22_, link_o_stitch_0__3__data__21_, link_o_stitch_0__3__data__20_, link_o_stitch_0__3__data__19_, link_o_stitch_0__3__data__18_, link_o_stitch_0__3__data__17_, link_o_stitch_0__3__data__16_, link_o_stitch_0__3__data__15_, link_o_stitch_0__3__data__14_, link_o_stitch_0__3__data__13_, link_o_stitch_0__3__data__12_, link_o_stitch_0__3__data__11_, link_o_stitch_0__3__data__10_, link_o_stitch_0__3__data__9_, link_o_stitch_0__3__data__8_, link_o_stitch_0__3__data__7_, link_o_stitch_0__3__data__6_, link_o_stitch_0__3__data__5_, link_o_stitch_0__3__data__4_, link_o_stitch_0__3__data__3_, link_o_stitch_0__3__data__2_, link_o_stitch_0__3__data__1_, link_o_stitch_0__3__data__0_, link_o_stitch_0__2__v_, link_o_stitch_0__2__ready_then_rev_, link_o_stitch_0__2__data__27_, link_o_stitch_0__2__data__26_, link_o_stitch_0__2__data__25_, link_o_stitch_0__2__data__24_, link_o_stitch_0__2__data__23_, link_o_stitch_0__2__data__22_, link_o_stitch_0__2__data__21_, link_o_stitch_0__2__data__20_, link_o_stitch_0__2__data__19_, link_o_stitch_0__2__data__18_, link_o_stitch_0__2__data__17_, link_o_stitch_0__2__data__16_, link_o_stitch_0__2__data__15_, link_o_stitch_0__2__data__14_, link_o_stitch_0__2__data__13_, link_o_stitch_0__2__data__12_, link_o_stitch_0__2__data__11_, link_o_stitch_0__2__data__10_, link_o_stitch_0__2__data__9_, link_o_stitch_0__2__data__8_, link_o_stitch_0__2__data__7_, link_o_stitch_0__2__data__6_, link_o_stitch_0__2__data__5_, link_o_stitch_0__2__data__4_, link_o_stitch_0__2__data__3_, link_o_stitch_0__2__data__2_, link_o_stitch_0__2__data__1_, link_o_stitch_0__2__data__0_, link_o_stitch_0__1__v_, link_o_stitch_0__1__ready_then_rev_, link_o_stitch_0__1__data__27_, link_o_stitch_0__1__data__26_, link_o_stitch_0__1__data__25_, link_o_stitch_0__1__data__24_, link_o_stitch_0__1__data__23_, link_o_stitch_0__1__data__22_, link_o_stitch_0__1__data__21_, link_o_stitch_0__1__data__20_, link_o_stitch_0__1__data__19_, link_o_stitch_0__1__data__18_, link_o_stitch_0__1__data__17_, link_o_stitch_0__1__data__16_, link_o_stitch_0__1__data__15_, link_o_stitch_0__1__data__14_, link_o_stitch_0__1__data__13_, link_o_stitch_0__1__data__12_, link_o_stitch_0__1__data__11_, link_o_stitch_0__1__data__10_, link_o_stitch_0__1__data__9_, link_o_stitch_0__1__data__8_, link_o_stitch_0__1__data__7_, link_o_stitch_0__1__data__6_, link_o_stitch_0__1__data__5_, link_o_stitch_0__1__data__4_, link_o_stitch_0__1__data__3_, link_o_stitch_0__1__data__2_, link_o_stitch_0__1__data__1_, link_o_stitch_0__1__data__0_, dst_v_o[0:0], link_o_stitch_0__0__ready_then_rev_, dst_data_o, link_o_stitch_0__0__data__1_, link_o_stitch_0__0__data__0_ }),
    .my_x_i(1'b0),
    .my_y_i(1'b1)
  );


  bsg_mesh_router_buffered_28_1_1_0_5_0d_0_30_00
  rof_1__efi2_fi7_coherence_network_channel_node
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .link_i({ src_v_i[1:1], 1'b0, src_data_i[51:26], 1'b1, src_data_i[51:51], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, link_o_stitch_0__2__v_, link_o_stitch_0__2__ready_then_rev_, link_o_stitch_0__2__data__27_, link_o_stitch_0__2__data__26_, link_o_stitch_0__2__data__25_, link_o_stitch_0__2__data__24_, link_o_stitch_0__2__data__23_, link_o_stitch_0__2__data__22_, link_o_stitch_0__2__data__21_, link_o_stitch_0__2__data__20_, link_o_stitch_0__2__data__19_, link_o_stitch_0__2__data__18_, link_o_stitch_0__2__data__17_, link_o_stitch_0__2__data__16_, link_o_stitch_0__2__data__15_, link_o_stitch_0__2__data__14_, link_o_stitch_0__2__data__13_, link_o_stitch_0__2__data__12_, link_o_stitch_0__2__data__11_, link_o_stitch_0__2__data__10_, link_o_stitch_0__2__data__9_, link_o_stitch_0__2__data__8_, link_o_stitch_0__2__data__7_, link_o_stitch_0__2__data__6_, link_o_stitch_0__2__data__5_, link_o_stitch_0__2__data__4_, link_o_stitch_0__2__data__3_, link_o_stitch_0__2__data__2_, link_o_stitch_0__2__data__1_, link_o_stitch_0__2__data__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .link_o({ link_o_stitch_1__4__v_, src_ready_o[1:1], link_o_stitch_1__4__data__27_, link_o_stitch_1__4__data__26_, link_o_stitch_1__4__data__25_, link_o_stitch_1__4__data__24_, link_o_stitch_1__4__data__23_, link_o_stitch_1__4__data__22_, link_o_stitch_1__4__data__21_, link_o_stitch_1__4__data__20_, link_o_stitch_1__4__data__19_, link_o_stitch_1__4__data__18_, link_o_stitch_1__4__data__17_, link_o_stitch_1__4__data__16_, link_o_stitch_1__4__data__15_, link_o_stitch_1__4__data__14_, link_o_stitch_1__4__data__13_, link_o_stitch_1__4__data__12_, link_o_stitch_1__4__data__11_, link_o_stitch_1__4__data__10_, link_o_stitch_1__4__data__9_, link_o_stitch_1__4__data__8_, link_o_stitch_1__4__data__7_, link_o_stitch_1__4__data__6_, link_o_stitch_1__4__data__5_, link_o_stitch_1__4__data__4_, link_o_stitch_1__4__data__3_, link_o_stitch_1__4__data__2_, link_o_stitch_1__4__data__1_, link_o_stitch_1__4__data__0_, link_o_stitch_1__3__v_, link_o_stitch_1__3__ready_then_rev_, link_o_stitch_1__3__data__27_, link_o_stitch_1__3__data__26_, link_o_stitch_1__3__data__25_, link_o_stitch_1__3__data__24_, link_o_stitch_1__3__data__23_, link_o_stitch_1__3__data__22_, link_o_stitch_1__3__data__21_, link_o_stitch_1__3__data__20_, link_o_stitch_1__3__data__19_, link_o_stitch_1__3__data__18_, link_o_stitch_1__3__data__17_, link_o_stitch_1__3__data__16_, link_o_stitch_1__3__data__15_, link_o_stitch_1__3__data__14_, link_o_stitch_1__3__data__13_, link_o_stitch_1__3__data__12_, link_o_stitch_1__3__data__11_, link_o_stitch_1__3__data__10_, link_o_stitch_1__3__data__9_, link_o_stitch_1__3__data__8_, link_o_stitch_1__3__data__7_, link_o_stitch_1__3__data__6_, link_o_stitch_1__3__data__5_, link_o_stitch_1__3__data__4_, link_o_stitch_1__3__data__3_, link_o_stitch_1__3__data__2_, link_o_stitch_1__3__data__1_, link_o_stitch_1__3__data__0_, link_o_stitch_1__2__v_, link_o_stitch_1__2__ready_then_rev_, link_o_stitch_1__2__data__27_, link_o_stitch_1__2__data__26_, link_o_stitch_1__2__data__25_, link_o_stitch_1__2__data__24_, link_o_stitch_1__2__data__23_, link_o_stitch_1__2__data__22_, link_o_stitch_1__2__data__21_, link_o_stitch_1__2__data__20_, link_o_stitch_1__2__data__19_, link_o_stitch_1__2__data__18_, link_o_stitch_1__2__data__17_, link_o_stitch_1__2__data__16_, link_o_stitch_1__2__data__15_, link_o_stitch_1__2__data__14_, link_o_stitch_1__2__data__13_, link_o_stitch_1__2__data__12_, link_o_stitch_1__2__data__11_, link_o_stitch_1__2__data__10_, link_o_stitch_1__2__data__9_, link_o_stitch_1__2__data__8_, link_o_stitch_1__2__data__7_, link_o_stitch_1__2__data__6_, link_o_stitch_1__2__data__5_, link_o_stitch_1__2__data__4_, link_o_stitch_1__2__data__3_, link_o_stitch_1__2__data__2_, link_o_stitch_1__2__data__1_, link_o_stitch_1__2__data__0_, link_i_stitch_0__2__v_, link_i_stitch_0__2__ready_then_rev_, link_i_stitch_0__2__data__27_, link_i_stitch_0__2__data__26_, link_i_stitch_0__2__data__25_, link_i_stitch_0__2__data__24_, link_i_stitch_0__2__data__23_, link_i_stitch_0__2__data__22_, link_i_stitch_0__2__data__21_, link_i_stitch_0__2__data__20_, link_i_stitch_0__2__data__19_, link_i_stitch_0__2__data__18_, link_i_stitch_0__2__data__17_, link_i_stitch_0__2__data__16_, link_i_stitch_0__2__data__15_, link_i_stitch_0__2__data__14_, link_i_stitch_0__2__data__13_, link_i_stitch_0__2__data__12_, link_i_stitch_0__2__data__11_, link_i_stitch_0__2__data__10_, link_i_stitch_0__2__data__9_, link_i_stitch_0__2__data__8_, link_i_stitch_0__2__data__7_, link_i_stitch_0__2__data__6_, link_i_stitch_0__2__data__5_, link_i_stitch_0__2__data__4_, link_i_stitch_0__2__data__3_, link_i_stitch_0__2__data__2_, link_i_stitch_0__2__data__1_, link_i_stitch_0__2__data__0_, link_o_stitch_1__0__v_, link_o_stitch_1__0__ready_then_rev_, link_o_stitch_1__0__data__27_, link_o_stitch_1__0__data__26_, link_o_stitch_1__0__data__25_, link_o_stitch_1__0__data__24_, link_o_stitch_1__0__data__23_, link_o_stitch_1__0__data__22_, link_o_stitch_1__0__data__21_, link_o_stitch_1__0__data__20_, link_o_stitch_1__0__data__19_, link_o_stitch_1__0__data__18_, link_o_stitch_1__0__data__17_, link_o_stitch_1__0__data__16_, link_o_stitch_1__0__data__15_, link_o_stitch_1__0__data__14_, link_o_stitch_1__0__data__13_, link_o_stitch_1__0__data__12_, link_o_stitch_1__0__data__11_, link_o_stitch_1__0__data__10_, link_o_stitch_1__0__data__9_, link_o_stitch_1__0__data__8_, link_o_stitch_1__0__data__7_, link_o_stitch_1__0__data__6_, link_o_stitch_1__0__data__5_, link_o_stitch_1__0__data__4_, link_o_stitch_1__0__data__3_, link_o_stitch_1__0__data__2_, link_o_stitch_1__0__data__1_, link_o_stitch_1__0__data__0_ }),
    .my_x_i(1'b1),
    .my_y_i(1'b1)
  );


endmodule



module bsg_mem_p136
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [135:0] w_data_i;
  input [0:0] r_addr_i;
  output [135:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [135:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10;
  reg [271:0] mem;
  assign r_data_o[135] = (N3)? mem[135] :
                         (N0)? mem[271] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[134] = (N3)? mem[134] :
                         (N0)? mem[270] : 1'b0;
  assign r_data_o[133] = (N3)? mem[133] :
                         (N0)? mem[269] : 1'b0;
  assign r_data_o[132] = (N3)? mem[132] :
                         (N0)? mem[268] : 1'b0;
  assign r_data_o[131] = (N3)? mem[131] :
                         (N0)? mem[267] : 1'b0;
  assign r_data_o[130] = (N3)? mem[130] :
                         (N0)? mem[266] : 1'b0;
  assign r_data_o[129] = (N3)? mem[129] :
                         (N0)? mem[265] : 1'b0;
  assign r_data_o[128] = (N3)? mem[128] :
                         (N0)? mem[264] : 1'b0;
  assign r_data_o[127] = (N3)? mem[127] :
                         (N0)? mem[263] : 1'b0;
  assign r_data_o[126] = (N3)? mem[126] :
                         (N0)? mem[262] : 1'b0;
  assign r_data_o[125] = (N3)? mem[125] :
                         (N0)? mem[261] : 1'b0;
  assign r_data_o[124] = (N3)? mem[124] :
                         (N0)? mem[260] : 1'b0;
  assign r_data_o[123] = (N3)? mem[123] :
                         (N0)? mem[259] : 1'b0;
  assign r_data_o[122] = (N3)? mem[122] :
                         (N0)? mem[258] : 1'b0;
  assign r_data_o[121] = (N3)? mem[121] :
                         (N0)? mem[257] : 1'b0;
  assign r_data_o[120] = (N3)? mem[120] :
                         (N0)? mem[256] : 1'b0;
  assign r_data_o[119] = (N3)? mem[119] :
                         (N0)? mem[255] : 1'b0;
  assign r_data_o[118] = (N3)? mem[118] :
                         (N0)? mem[254] : 1'b0;
  assign r_data_o[117] = (N3)? mem[117] :
                         (N0)? mem[253] : 1'b0;
  assign r_data_o[116] = (N3)? mem[116] :
                         (N0)? mem[252] : 1'b0;
  assign r_data_o[115] = (N3)? mem[115] :
                         (N0)? mem[251] : 1'b0;
  assign r_data_o[114] = (N3)? mem[114] :
                         (N0)? mem[250] : 1'b0;
  assign r_data_o[113] = (N3)? mem[113] :
                         (N0)? mem[249] : 1'b0;
  assign r_data_o[112] = (N3)? mem[112] :
                         (N0)? mem[248] : 1'b0;
  assign r_data_o[111] = (N3)? mem[111] :
                         (N0)? mem[247] : 1'b0;
  assign r_data_o[110] = (N3)? mem[110] :
                         (N0)? mem[246] : 1'b0;
  assign r_data_o[109] = (N3)? mem[109] :
                         (N0)? mem[245] : 1'b0;
  assign r_data_o[108] = (N3)? mem[108] :
                         (N0)? mem[244] : 1'b0;
  assign r_data_o[107] = (N3)? mem[107] :
                         (N0)? mem[243] : 1'b0;
  assign r_data_o[106] = (N3)? mem[106] :
                         (N0)? mem[242] : 1'b0;
  assign r_data_o[105] = (N3)? mem[105] :
                         (N0)? mem[241] : 1'b0;
  assign r_data_o[104] = (N3)? mem[104] :
                         (N0)? mem[240] : 1'b0;
  assign r_data_o[103] = (N3)? mem[103] :
                         (N0)? mem[239] : 1'b0;
  assign r_data_o[102] = (N3)? mem[102] :
                         (N0)? mem[238] : 1'b0;
  assign r_data_o[101] = (N3)? mem[101] :
                         (N0)? mem[237] : 1'b0;
  assign r_data_o[100] = (N3)? mem[100] :
                         (N0)? mem[236] : 1'b0;
  assign r_data_o[99] = (N3)? mem[99] :
                        (N0)? mem[235] : 1'b0;
  assign r_data_o[98] = (N3)? mem[98] :
                        (N0)? mem[234] : 1'b0;
  assign r_data_o[97] = (N3)? mem[97] :
                        (N0)? mem[233] : 1'b0;
  assign r_data_o[96] = (N3)? mem[96] :
                        (N0)? mem[232] : 1'b0;
  assign r_data_o[95] = (N3)? mem[95] :
                        (N0)? mem[231] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] :
                        (N0)? mem[230] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] :
                        (N0)? mem[229] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] :
                        (N0)? mem[228] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] :
                        (N0)? mem[227] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] :
                        (N0)? mem[226] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] :
                        (N0)? mem[225] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] :
                        (N0)? mem[224] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] :
                        (N0)? mem[223] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] :
                        (N0)? mem[222] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] :
                        (N0)? mem[221] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] :
                        (N0)? mem[220] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] :
                        (N0)? mem[219] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] :
                        (N0)? mem[218] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] :
                        (N0)? mem[217] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] :
                        (N0)? mem[216] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] :
                        (N0)? mem[215] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] :
                        (N0)? mem[214] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] :
                        (N0)? mem[213] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] :
                        (N0)? mem[212] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] :
                        (N0)? mem[211] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] :
                        (N0)? mem[210] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] :
                        (N0)? mem[209] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] :
                        (N0)? mem[208] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] :
                        (N0)? mem[207] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] :
                        (N0)? mem[206] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] :
                        (N0)? mem[205] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] :
                        (N0)? mem[204] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] :
                        (N0)? mem[203] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] :
                        (N0)? mem[202] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] :
                        (N0)? mem[201] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] :
                        (N0)? mem[200] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] :
                        (N0)? mem[199] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] :
                        (N0)? mem[198] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] :
                        (N0)? mem[197] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] :
                        (N0)? mem[196] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] :
                        (N0)? mem[195] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] :
                        (N0)? mem[194] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] :
                        (N0)? mem[193] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] :
                        (N0)? mem[192] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] :
                        (N0)? mem[191] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] :
                        (N0)? mem[190] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] :
                        (N0)? mem[189] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] :
                        (N0)? mem[188] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] :
                        (N0)? mem[187] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] :
                        (N0)? mem[186] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] :
                        (N0)? mem[185] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] :
                        (N0)? mem[184] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] :
                        (N0)? mem[183] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] :
                        (N0)? mem[182] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] :
                        (N0)? mem[181] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] :
                        (N0)? mem[180] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] :
                        (N0)? mem[179] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] :
                        (N0)? mem[178] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] :
                        (N0)? mem[177] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] :
                        (N0)? mem[176] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] :
                        (N0)? mem[175] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] :
                        (N0)? mem[174] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] :
                        (N0)? mem[173] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] :
                        (N0)? mem[172] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] :
                        (N0)? mem[171] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] :
                        (N0)? mem[170] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] :
                        (N0)? mem[169] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] :
                        (N0)? mem[168] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] :
                        (N0)? mem[167] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] :
                        (N0)? mem[166] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] :
                        (N0)? mem[165] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] :
                        (N0)? mem[164] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] :
                        (N0)? mem[163] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] :
                        (N0)? mem[162] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] :
                        (N0)? mem[161] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] :
                        (N0)? mem[160] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] :
                        (N0)? mem[159] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] :
                        (N0)? mem[158] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] :
                        (N0)? mem[157] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] :
                        (N0)? mem[156] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] :
                        (N0)? mem[155] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] :
                        (N0)? mem[154] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] :
                        (N0)? mem[153] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] :
                        (N0)? mem[152] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] :
                        (N0)? mem[151] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] :
                        (N0)? mem[150] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] :
                        (N0)? mem[149] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] :
                        (N0)? mem[148] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] :
                        (N0)? mem[147] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] :
                        (N0)? mem[146] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] :
                       (N0)? mem[145] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] :
                       (N0)? mem[144] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] :
                       (N0)? mem[143] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] :
                       (N0)? mem[142] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] :
                       (N0)? mem[141] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] :
                       (N0)? mem[140] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] :
                       (N0)? mem[139] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] :
                       (N0)? mem[138] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] :
                       (N0)? mem[137] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] :
                       (N0)? mem[136] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], N5, N5 } :
                               (N2)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N9) begin
      { mem[271:173], mem[136:136] } <= { w_data_i[135:37], w_data_i[0:0] };
    end
    if(N10) begin
      { mem[172:137] } <= { w_data_i[36:1] };
    end
    if(N7) begin
      { mem[135:37], mem[0:0] } <= { w_data_i[135:37], w_data_i[0:0] };
    end
    if(N8) begin
      { mem[36:1] } <= { w_data_i[36:1] };
    end
  end


endmodule



module bsg_mem_1r1w_width_p136_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [135:0] w_data_i;
  input [0:0] r_addr_i;
  output [135:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [135:0] r_data_o;

  bsg_mem_p136
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p136
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [135:0] data_i;
  output [135:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [135:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p136_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 :
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 :
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 :
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 :
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 :
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 :
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end
    if(N9) begin
      tail_r <= N10;
    end
    if(N11) begin
      head_r <= N12;
    end
  end


endmodule



module bsg_mux_one_hot_width_p136_els_p4
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [543:0] data_i;
  input [3:0] sel_one_hot_i;
  output [135:0] data_o;
  wire [135:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271;
  wire [543:0] data_masked;
  assign data_masked[135] = data_i[135] & sel_one_hot_i[0];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[0];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[0];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[0];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[0];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[0];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[0];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[0];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[0];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[0];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[0];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[0];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[0];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[0];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[0];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[0];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[0];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[0];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[0];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[0];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[0];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[0];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[0];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[0];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[0];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[0];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[0];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[0];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[0];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[0];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[0];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[0];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[0];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[0];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[0];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[0];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[0];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[0];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[0];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[0];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[0];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[0];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[0];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[0];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[0];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[0];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[0];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[0];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[0];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[0];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[0];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[0];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[0];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[0];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[0];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[0];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[0];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[0];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[0];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[0];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[0];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[0];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[0];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[0];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[0];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[0];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[0];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[0];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[1];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[1];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[1];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[1];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[1];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[1];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[1];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[1];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[1];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[1];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[1];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[1];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[1];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[1];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[1];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[1];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[1];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[1];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[1];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[1];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[1];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[1];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[1];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[1];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[1];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[1];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[1];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[1];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[1];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[1];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[1];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[1];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[1];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[1];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[1];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[1];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[1];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[1];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[1];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[1];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[1];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[1];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[1];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[1];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[1];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[1];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[1];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[1];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[1];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[1];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[1];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[1];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[1];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[1];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[1];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[1];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[1];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[1];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[1];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[1];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[1];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[1];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[1];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[1];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[1];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[1];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[1];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[1];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[1];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[1];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[1];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[1];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[1];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[1];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[1];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[1];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[1];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[1];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[1];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[1];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[1];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[1];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[1];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[1];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[1];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[1];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[1];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[1];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[1];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[1];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[1];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[1];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[1];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[1];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[1];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[1];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[1];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[1];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[1];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[1];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[1];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[1];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[1];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[1];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[1];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[1];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[1];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[1];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[1];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[1];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[1];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[1];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[1];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[1];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[1];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[1];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[1];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[1];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[1];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[1];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[1];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[1];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[1];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[1];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[1];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[1];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[1];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[1];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[1];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[1];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[1];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[1];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[1];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[1];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[1];
  assign data_masked[407] = data_i[407] & sel_one_hot_i[2];
  assign data_masked[406] = data_i[406] & sel_one_hot_i[2];
  assign data_masked[405] = data_i[405] & sel_one_hot_i[2];
  assign data_masked[404] = data_i[404] & sel_one_hot_i[2];
  assign data_masked[403] = data_i[403] & sel_one_hot_i[2];
  assign data_masked[402] = data_i[402] & sel_one_hot_i[2];
  assign data_masked[401] = data_i[401] & sel_one_hot_i[2];
  assign data_masked[400] = data_i[400] & sel_one_hot_i[2];
  assign data_masked[399] = data_i[399] & sel_one_hot_i[2];
  assign data_masked[398] = data_i[398] & sel_one_hot_i[2];
  assign data_masked[397] = data_i[397] & sel_one_hot_i[2];
  assign data_masked[396] = data_i[396] & sel_one_hot_i[2];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[2];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[2];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[2];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[2];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[2];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[2];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[2];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[2];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[2];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[2];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[2];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[2];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[2];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[2];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[2];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[2];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[2];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[2];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[2];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[2];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[2];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[2];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[2];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[2];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[2];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[2];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[2];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[2];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[2];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[2];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[2];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[2];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[2];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[2];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[2];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[2];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[2];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[2];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[2];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[2];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[2];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[2];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[2];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[2];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[2];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[2];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[2];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[2];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[2];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[2];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[2];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[2];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[2];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[2];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[2];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[2];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[2];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[2];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[2];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[2];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[2];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[2];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[2];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[2];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[2];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[2];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[2];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[2];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[2];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[2];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[2];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[2];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[2];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[2];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[2];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[2];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[2];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[2];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[2];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[2];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[2];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[2];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[2];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[2];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[2];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[2];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[2];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[2];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[2];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[2];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[2];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[2];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[2];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[2];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[2];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[2];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[2];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[2];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[2];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[2];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[2];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[2];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[2];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[2];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[2];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[2];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[2];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[2];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[2];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[2];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[2];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[2];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[2];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[2];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[2];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[2];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[2];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[2];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[2];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[2];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[2];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[2];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[2];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[2];
  assign data_masked[543] = data_i[543] & sel_one_hot_i[3];
  assign data_masked[542] = data_i[542] & sel_one_hot_i[3];
  assign data_masked[541] = data_i[541] & sel_one_hot_i[3];
  assign data_masked[540] = data_i[540] & sel_one_hot_i[3];
  assign data_masked[539] = data_i[539] & sel_one_hot_i[3];
  assign data_masked[538] = data_i[538] & sel_one_hot_i[3];
  assign data_masked[537] = data_i[537] & sel_one_hot_i[3];
  assign data_masked[536] = data_i[536] & sel_one_hot_i[3];
  assign data_masked[535] = data_i[535] & sel_one_hot_i[3];
  assign data_masked[534] = data_i[534] & sel_one_hot_i[3];
  assign data_masked[533] = data_i[533] & sel_one_hot_i[3];
  assign data_masked[532] = data_i[532] & sel_one_hot_i[3];
  assign data_masked[531] = data_i[531] & sel_one_hot_i[3];
  assign data_masked[530] = data_i[530] & sel_one_hot_i[3];
  assign data_masked[529] = data_i[529] & sel_one_hot_i[3];
  assign data_masked[528] = data_i[528] & sel_one_hot_i[3];
  assign data_masked[527] = data_i[527] & sel_one_hot_i[3];
  assign data_masked[526] = data_i[526] & sel_one_hot_i[3];
  assign data_masked[525] = data_i[525] & sel_one_hot_i[3];
  assign data_masked[524] = data_i[524] & sel_one_hot_i[3];
  assign data_masked[523] = data_i[523] & sel_one_hot_i[3];
  assign data_masked[522] = data_i[522] & sel_one_hot_i[3];
  assign data_masked[521] = data_i[521] & sel_one_hot_i[3];
  assign data_masked[520] = data_i[520] & sel_one_hot_i[3];
  assign data_masked[519] = data_i[519] & sel_one_hot_i[3];
  assign data_masked[518] = data_i[518] & sel_one_hot_i[3];
  assign data_masked[517] = data_i[517] & sel_one_hot_i[3];
  assign data_masked[516] = data_i[516] & sel_one_hot_i[3];
  assign data_masked[515] = data_i[515] & sel_one_hot_i[3];
  assign data_masked[514] = data_i[514] & sel_one_hot_i[3];
  assign data_masked[513] = data_i[513] & sel_one_hot_i[3];
  assign data_masked[512] = data_i[512] & sel_one_hot_i[3];
  assign data_masked[511] = data_i[511] & sel_one_hot_i[3];
  assign data_masked[510] = data_i[510] & sel_one_hot_i[3];
  assign data_masked[509] = data_i[509] & sel_one_hot_i[3];
  assign data_masked[508] = data_i[508] & sel_one_hot_i[3];
  assign data_masked[507] = data_i[507] & sel_one_hot_i[3];
  assign data_masked[506] = data_i[506] & sel_one_hot_i[3];
  assign data_masked[505] = data_i[505] & sel_one_hot_i[3];
  assign data_masked[504] = data_i[504] & sel_one_hot_i[3];
  assign data_masked[503] = data_i[503] & sel_one_hot_i[3];
  assign data_masked[502] = data_i[502] & sel_one_hot_i[3];
  assign data_masked[501] = data_i[501] & sel_one_hot_i[3];
  assign data_masked[500] = data_i[500] & sel_one_hot_i[3];
  assign data_masked[499] = data_i[499] & sel_one_hot_i[3];
  assign data_masked[498] = data_i[498] & sel_one_hot_i[3];
  assign data_masked[497] = data_i[497] & sel_one_hot_i[3];
  assign data_masked[496] = data_i[496] & sel_one_hot_i[3];
  assign data_masked[495] = data_i[495] & sel_one_hot_i[3];
  assign data_masked[494] = data_i[494] & sel_one_hot_i[3];
  assign data_masked[493] = data_i[493] & sel_one_hot_i[3];
  assign data_masked[492] = data_i[492] & sel_one_hot_i[3];
  assign data_masked[491] = data_i[491] & sel_one_hot_i[3];
  assign data_masked[490] = data_i[490] & sel_one_hot_i[3];
  assign data_masked[489] = data_i[489] & sel_one_hot_i[3];
  assign data_masked[488] = data_i[488] & sel_one_hot_i[3];
  assign data_masked[487] = data_i[487] & sel_one_hot_i[3];
  assign data_masked[486] = data_i[486] & sel_one_hot_i[3];
  assign data_masked[485] = data_i[485] & sel_one_hot_i[3];
  assign data_masked[484] = data_i[484] & sel_one_hot_i[3];
  assign data_masked[483] = data_i[483] & sel_one_hot_i[3];
  assign data_masked[482] = data_i[482] & sel_one_hot_i[3];
  assign data_masked[481] = data_i[481] & sel_one_hot_i[3];
  assign data_masked[480] = data_i[480] & sel_one_hot_i[3];
  assign data_masked[479] = data_i[479] & sel_one_hot_i[3];
  assign data_masked[478] = data_i[478] & sel_one_hot_i[3];
  assign data_masked[477] = data_i[477] & sel_one_hot_i[3];
  assign data_masked[476] = data_i[476] & sel_one_hot_i[3];
  assign data_masked[475] = data_i[475] & sel_one_hot_i[3];
  assign data_masked[474] = data_i[474] & sel_one_hot_i[3];
  assign data_masked[473] = data_i[473] & sel_one_hot_i[3];
  assign data_masked[472] = data_i[472] & sel_one_hot_i[3];
  assign data_masked[471] = data_i[471] & sel_one_hot_i[3];
  assign data_masked[470] = data_i[470] & sel_one_hot_i[3];
  assign data_masked[469] = data_i[469] & sel_one_hot_i[3];
  assign data_masked[468] = data_i[468] & sel_one_hot_i[3];
  assign data_masked[467] = data_i[467] & sel_one_hot_i[3];
  assign data_masked[466] = data_i[466] & sel_one_hot_i[3];
  assign data_masked[465] = data_i[465] & sel_one_hot_i[3];
  assign data_masked[464] = data_i[464] & sel_one_hot_i[3];
  assign data_masked[463] = data_i[463] & sel_one_hot_i[3];
  assign data_masked[462] = data_i[462] & sel_one_hot_i[3];
  assign data_masked[461] = data_i[461] & sel_one_hot_i[3];
  assign data_masked[460] = data_i[460] & sel_one_hot_i[3];
  assign data_masked[459] = data_i[459] & sel_one_hot_i[3];
  assign data_masked[458] = data_i[458] & sel_one_hot_i[3];
  assign data_masked[457] = data_i[457] & sel_one_hot_i[3];
  assign data_masked[456] = data_i[456] & sel_one_hot_i[3];
  assign data_masked[455] = data_i[455] & sel_one_hot_i[3];
  assign data_masked[454] = data_i[454] & sel_one_hot_i[3];
  assign data_masked[453] = data_i[453] & sel_one_hot_i[3];
  assign data_masked[452] = data_i[452] & sel_one_hot_i[3];
  assign data_masked[451] = data_i[451] & sel_one_hot_i[3];
  assign data_masked[450] = data_i[450] & sel_one_hot_i[3];
  assign data_masked[449] = data_i[449] & sel_one_hot_i[3];
  assign data_masked[448] = data_i[448] & sel_one_hot_i[3];
  assign data_masked[447] = data_i[447] & sel_one_hot_i[3];
  assign data_masked[446] = data_i[446] & sel_one_hot_i[3];
  assign data_masked[445] = data_i[445] & sel_one_hot_i[3];
  assign data_masked[444] = data_i[444] & sel_one_hot_i[3];
  assign data_masked[443] = data_i[443] & sel_one_hot_i[3];
  assign data_masked[442] = data_i[442] & sel_one_hot_i[3];
  assign data_masked[441] = data_i[441] & sel_one_hot_i[3];
  assign data_masked[440] = data_i[440] & sel_one_hot_i[3];
  assign data_masked[439] = data_i[439] & sel_one_hot_i[3];
  assign data_masked[438] = data_i[438] & sel_one_hot_i[3];
  assign data_masked[437] = data_i[437] & sel_one_hot_i[3];
  assign data_masked[436] = data_i[436] & sel_one_hot_i[3];
  assign data_masked[435] = data_i[435] & sel_one_hot_i[3];
  assign data_masked[434] = data_i[434] & sel_one_hot_i[3];
  assign data_masked[433] = data_i[433] & sel_one_hot_i[3];
  assign data_masked[432] = data_i[432] & sel_one_hot_i[3];
  assign data_masked[431] = data_i[431] & sel_one_hot_i[3];
  assign data_masked[430] = data_i[430] & sel_one_hot_i[3];
  assign data_masked[429] = data_i[429] & sel_one_hot_i[3];
  assign data_masked[428] = data_i[428] & sel_one_hot_i[3];
  assign data_masked[427] = data_i[427] & sel_one_hot_i[3];
  assign data_masked[426] = data_i[426] & sel_one_hot_i[3];
  assign data_masked[425] = data_i[425] & sel_one_hot_i[3];
  assign data_masked[424] = data_i[424] & sel_one_hot_i[3];
  assign data_masked[423] = data_i[423] & sel_one_hot_i[3];
  assign data_masked[422] = data_i[422] & sel_one_hot_i[3];
  assign data_masked[421] = data_i[421] & sel_one_hot_i[3];
  assign data_masked[420] = data_i[420] & sel_one_hot_i[3];
  assign data_masked[419] = data_i[419] & sel_one_hot_i[3];
  assign data_masked[418] = data_i[418] & sel_one_hot_i[3];
  assign data_masked[417] = data_i[417] & sel_one_hot_i[3];
  assign data_masked[416] = data_i[416] & sel_one_hot_i[3];
  assign data_masked[415] = data_i[415] & sel_one_hot_i[3];
  assign data_masked[414] = data_i[414] & sel_one_hot_i[3];
  assign data_masked[413] = data_i[413] & sel_one_hot_i[3];
  assign data_masked[412] = data_i[412] & sel_one_hot_i[3];
  assign data_masked[411] = data_i[411] & sel_one_hot_i[3];
  assign data_masked[410] = data_i[410] & sel_one_hot_i[3];
  assign data_masked[409] = data_i[409] & sel_one_hot_i[3];
  assign data_masked[408] = data_i[408] & sel_one_hot_i[3];
  assign data_o[0] = N1 | data_masked[0];
  assign N1 = N0 | data_masked[136];
  assign N0 = data_masked[408] | data_masked[272];
  assign data_o[1] = N3 | data_masked[1];
  assign N3 = N2 | data_masked[137];
  assign N2 = data_masked[409] | data_masked[273];
  assign data_o[2] = N5 | data_masked[2];
  assign N5 = N4 | data_masked[138];
  assign N4 = data_masked[410] | data_masked[274];
  assign data_o[3] = N7 | data_masked[3];
  assign N7 = N6 | data_masked[139];
  assign N6 = data_masked[411] | data_masked[275];
  assign data_o[4] = N9 | data_masked[4];
  assign N9 = N8 | data_masked[140];
  assign N8 = data_masked[412] | data_masked[276];
  assign data_o[5] = N11 | data_masked[5];
  assign N11 = N10 | data_masked[141];
  assign N10 = data_masked[413] | data_masked[277];
  assign data_o[6] = N13 | data_masked[6];
  assign N13 = N12 | data_masked[142];
  assign N12 = data_masked[414] | data_masked[278];
  assign data_o[7] = N15 | data_masked[7];
  assign N15 = N14 | data_masked[143];
  assign N14 = data_masked[415] | data_masked[279];
  assign data_o[8] = N17 | data_masked[8];
  assign N17 = N16 | data_masked[144];
  assign N16 = data_masked[416] | data_masked[280];
  assign data_o[9] = N19 | data_masked[9];
  assign N19 = N18 | data_masked[145];
  assign N18 = data_masked[417] | data_masked[281];
  assign data_o[10] = N21 | data_masked[10];
  assign N21 = N20 | data_masked[146];
  assign N20 = data_masked[418] | data_masked[282];
  assign data_o[11] = N23 | data_masked[11];
  assign N23 = N22 | data_masked[147];
  assign N22 = data_masked[419] | data_masked[283];
  assign data_o[12] = N25 | data_masked[12];
  assign N25 = N24 | data_masked[148];
  assign N24 = data_masked[420] | data_masked[284];
  assign data_o[13] = N27 | data_masked[13];
  assign N27 = N26 | data_masked[149];
  assign N26 = data_masked[421] | data_masked[285];
  assign data_o[14] = N29 | data_masked[14];
  assign N29 = N28 | data_masked[150];
  assign N28 = data_masked[422] | data_masked[286];
  assign data_o[15] = N31 | data_masked[15];
  assign N31 = N30 | data_masked[151];
  assign N30 = data_masked[423] | data_masked[287];
  assign data_o[16] = N33 | data_masked[16];
  assign N33 = N32 | data_masked[152];
  assign N32 = data_masked[424] | data_masked[288];
  assign data_o[17] = N35 | data_masked[17];
  assign N35 = N34 | data_masked[153];
  assign N34 = data_masked[425] | data_masked[289];
  assign data_o[18] = N37 | data_masked[18];
  assign N37 = N36 | data_masked[154];
  assign N36 = data_masked[426] | data_masked[290];
  assign data_o[19] = N39 | data_masked[19];
  assign N39 = N38 | data_masked[155];
  assign N38 = data_masked[427] | data_masked[291];
  assign data_o[20] = N41 | data_masked[20];
  assign N41 = N40 | data_masked[156];
  assign N40 = data_masked[428] | data_masked[292];
  assign data_o[21] = N43 | data_masked[21];
  assign N43 = N42 | data_masked[157];
  assign N42 = data_masked[429] | data_masked[293];
  assign data_o[22] = N45 | data_masked[22];
  assign N45 = N44 | data_masked[158];
  assign N44 = data_masked[430] | data_masked[294];
  assign data_o[23] = N47 | data_masked[23];
  assign N47 = N46 | data_masked[159];
  assign N46 = data_masked[431] | data_masked[295];
  assign data_o[24] = N49 | data_masked[24];
  assign N49 = N48 | data_masked[160];
  assign N48 = data_masked[432] | data_masked[296];
  assign data_o[25] = N51 | data_masked[25];
  assign N51 = N50 | data_masked[161];
  assign N50 = data_masked[433] | data_masked[297];
  assign data_o[26] = N53 | data_masked[26];
  assign N53 = N52 | data_masked[162];
  assign N52 = data_masked[434] | data_masked[298];
  assign data_o[27] = N55 | data_masked[27];
  assign N55 = N54 | data_masked[163];
  assign N54 = data_masked[435] | data_masked[299];
  assign data_o[28] = N57 | data_masked[28];
  assign N57 = N56 | data_masked[164];
  assign N56 = data_masked[436] | data_masked[300];
  assign data_o[29] = N59 | data_masked[29];
  assign N59 = N58 | data_masked[165];
  assign N58 = data_masked[437] | data_masked[301];
  assign data_o[30] = N61 | data_masked[30];
  assign N61 = N60 | data_masked[166];
  assign N60 = data_masked[438] | data_masked[302];
  assign data_o[31] = N63 | data_masked[31];
  assign N63 = N62 | data_masked[167];
  assign N62 = data_masked[439] | data_masked[303];
  assign data_o[32] = N65 | data_masked[32];
  assign N65 = N64 | data_masked[168];
  assign N64 = data_masked[440] | data_masked[304];
  assign data_o[33] = N67 | data_masked[33];
  assign N67 = N66 | data_masked[169];
  assign N66 = data_masked[441] | data_masked[305];
  assign data_o[34] = N69 | data_masked[34];
  assign N69 = N68 | data_masked[170];
  assign N68 = data_masked[442] | data_masked[306];
  assign data_o[35] = N71 | data_masked[35];
  assign N71 = N70 | data_masked[171];
  assign N70 = data_masked[443] | data_masked[307];
  assign data_o[36] = N73 | data_masked[36];
  assign N73 = N72 | data_masked[172];
  assign N72 = data_masked[444] | data_masked[308];
  assign data_o[37] = N75 | data_masked[37];
  assign N75 = N74 | data_masked[173];
  assign N74 = data_masked[445] | data_masked[309];
  assign data_o[38] = N77 | data_masked[38];
  assign N77 = N76 | data_masked[174];
  assign N76 = data_masked[446] | data_masked[310];
  assign data_o[39] = N79 | data_masked[39];
  assign N79 = N78 | data_masked[175];
  assign N78 = data_masked[447] | data_masked[311];
  assign data_o[40] = N81 | data_masked[40];
  assign N81 = N80 | data_masked[176];
  assign N80 = data_masked[448] | data_masked[312];
  assign data_o[41] = N83 | data_masked[41];
  assign N83 = N82 | data_masked[177];
  assign N82 = data_masked[449] | data_masked[313];
  assign data_o[42] = N85 | data_masked[42];
  assign N85 = N84 | data_masked[178];
  assign N84 = data_masked[450] | data_masked[314];
  assign data_o[43] = N87 | data_masked[43];
  assign N87 = N86 | data_masked[179];
  assign N86 = data_masked[451] | data_masked[315];
  assign data_o[44] = N89 | data_masked[44];
  assign N89 = N88 | data_masked[180];
  assign N88 = data_masked[452] | data_masked[316];
  assign data_o[45] = N91 | data_masked[45];
  assign N91 = N90 | data_masked[181];
  assign N90 = data_masked[453] | data_masked[317];
  assign data_o[46] = N93 | data_masked[46];
  assign N93 = N92 | data_masked[182];
  assign N92 = data_masked[454] | data_masked[318];
  assign data_o[47] = N95 | data_masked[47];
  assign N95 = N94 | data_masked[183];
  assign N94 = data_masked[455] | data_masked[319];
  assign data_o[48] = N97 | data_masked[48];
  assign N97 = N96 | data_masked[184];
  assign N96 = data_masked[456] | data_masked[320];
  assign data_o[49] = N99 | data_masked[49];
  assign N99 = N98 | data_masked[185];
  assign N98 = data_masked[457] | data_masked[321];
  assign data_o[50] = N101 | data_masked[50];
  assign N101 = N100 | data_masked[186];
  assign N100 = data_masked[458] | data_masked[322];
  assign data_o[51] = N103 | data_masked[51];
  assign N103 = N102 | data_masked[187];
  assign N102 = data_masked[459] | data_masked[323];
  assign data_o[52] = N105 | data_masked[52];
  assign N105 = N104 | data_masked[188];
  assign N104 = data_masked[460] | data_masked[324];
  assign data_o[53] = N107 | data_masked[53];
  assign N107 = N106 | data_masked[189];
  assign N106 = data_masked[461] | data_masked[325];
  assign data_o[54] = N109 | data_masked[54];
  assign N109 = N108 | data_masked[190];
  assign N108 = data_masked[462] | data_masked[326];
  assign data_o[55] = N111 | data_masked[55];
  assign N111 = N110 | data_masked[191];
  assign N110 = data_masked[463] | data_masked[327];
  assign data_o[56] = N113 | data_masked[56];
  assign N113 = N112 | data_masked[192];
  assign N112 = data_masked[464] | data_masked[328];
  assign data_o[57] = N115 | data_masked[57];
  assign N115 = N114 | data_masked[193];
  assign N114 = data_masked[465] | data_masked[329];
  assign data_o[58] = N117 | data_masked[58];
  assign N117 = N116 | data_masked[194];
  assign N116 = data_masked[466] | data_masked[330];
  assign data_o[59] = N119 | data_masked[59];
  assign N119 = N118 | data_masked[195];
  assign N118 = data_masked[467] | data_masked[331];
  assign data_o[60] = N121 | data_masked[60];
  assign N121 = N120 | data_masked[196];
  assign N120 = data_masked[468] | data_masked[332];
  assign data_o[61] = N123 | data_masked[61];
  assign N123 = N122 | data_masked[197];
  assign N122 = data_masked[469] | data_masked[333];
  assign data_o[62] = N125 | data_masked[62];
  assign N125 = N124 | data_masked[198];
  assign N124 = data_masked[470] | data_masked[334];
  assign data_o[63] = N127 | data_masked[63];
  assign N127 = N126 | data_masked[199];
  assign N126 = data_masked[471] | data_masked[335];
  assign data_o[64] = N129 | data_masked[64];
  assign N129 = N128 | data_masked[200];
  assign N128 = data_masked[472] | data_masked[336];
  assign data_o[65] = N131 | data_masked[65];
  assign N131 = N130 | data_masked[201];
  assign N130 = data_masked[473] | data_masked[337];
  assign data_o[66] = N133 | data_masked[66];
  assign N133 = N132 | data_masked[202];
  assign N132 = data_masked[474] | data_masked[338];
  assign data_o[67] = N135 | data_masked[67];
  assign N135 = N134 | data_masked[203];
  assign N134 = data_masked[475] | data_masked[339];
  assign data_o[68] = N137 | data_masked[68];
  assign N137 = N136 | data_masked[204];
  assign N136 = data_masked[476] | data_masked[340];
  assign data_o[69] = N139 | data_masked[69];
  assign N139 = N138 | data_masked[205];
  assign N138 = data_masked[477] | data_masked[341];
  assign data_o[70] = N141 | data_masked[70];
  assign N141 = N140 | data_masked[206];
  assign N140 = data_masked[478] | data_masked[342];
  assign data_o[71] = N143 | data_masked[71];
  assign N143 = N142 | data_masked[207];
  assign N142 = data_masked[479] | data_masked[343];
  assign data_o[72] = N145 | data_masked[72];
  assign N145 = N144 | data_masked[208];
  assign N144 = data_masked[480] | data_masked[344];
  assign data_o[73] = N147 | data_masked[73];
  assign N147 = N146 | data_masked[209];
  assign N146 = data_masked[481] | data_masked[345];
  assign data_o[74] = N149 | data_masked[74];
  assign N149 = N148 | data_masked[210];
  assign N148 = data_masked[482] | data_masked[346];
  assign data_o[75] = N151 | data_masked[75];
  assign N151 = N150 | data_masked[211];
  assign N150 = data_masked[483] | data_masked[347];
  assign data_o[76] = N153 | data_masked[76];
  assign N153 = N152 | data_masked[212];
  assign N152 = data_masked[484] | data_masked[348];
  assign data_o[77] = N155 | data_masked[77];
  assign N155 = N154 | data_masked[213];
  assign N154 = data_masked[485] | data_masked[349];
  assign data_o[78] = N157 | data_masked[78];
  assign N157 = N156 | data_masked[214];
  assign N156 = data_masked[486] | data_masked[350];
  assign data_o[79] = N159 | data_masked[79];
  assign N159 = N158 | data_masked[215];
  assign N158 = data_masked[487] | data_masked[351];
  assign data_o[80] = N161 | data_masked[80];
  assign N161 = N160 | data_masked[216];
  assign N160 = data_masked[488] | data_masked[352];
  assign data_o[81] = N163 | data_masked[81];
  assign N163 = N162 | data_masked[217];
  assign N162 = data_masked[489] | data_masked[353];
  assign data_o[82] = N165 | data_masked[82];
  assign N165 = N164 | data_masked[218];
  assign N164 = data_masked[490] | data_masked[354];
  assign data_o[83] = N167 | data_masked[83];
  assign N167 = N166 | data_masked[219];
  assign N166 = data_masked[491] | data_masked[355];
  assign data_o[84] = N169 | data_masked[84];
  assign N169 = N168 | data_masked[220];
  assign N168 = data_masked[492] | data_masked[356];
  assign data_o[85] = N171 | data_masked[85];
  assign N171 = N170 | data_masked[221];
  assign N170 = data_masked[493] | data_masked[357];
  assign data_o[86] = N173 | data_masked[86];
  assign N173 = N172 | data_masked[222];
  assign N172 = data_masked[494] | data_masked[358];
  assign data_o[87] = N175 | data_masked[87];
  assign N175 = N174 | data_masked[223];
  assign N174 = data_masked[495] | data_masked[359];
  assign data_o[88] = N177 | data_masked[88];
  assign N177 = N176 | data_masked[224];
  assign N176 = data_masked[496] | data_masked[360];
  assign data_o[89] = N179 | data_masked[89];
  assign N179 = N178 | data_masked[225];
  assign N178 = data_masked[497] | data_masked[361];
  assign data_o[90] = N181 | data_masked[90];
  assign N181 = N180 | data_masked[226];
  assign N180 = data_masked[498] | data_masked[362];
  assign data_o[91] = N183 | data_masked[91];
  assign N183 = N182 | data_masked[227];
  assign N182 = data_masked[499] | data_masked[363];
  assign data_o[92] = N185 | data_masked[92];
  assign N185 = N184 | data_masked[228];
  assign N184 = data_masked[500] | data_masked[364];
  assign data_o[93] = N187 | data_masked[93];
  assign N187 = N186 | data_masked[229];
  assign N186 = data_masked[501] | data_masked[365];
  assign data_o[94] = N189 | data_masked[94];
  assign N189 = N188 | data_masked[230];
  assign N188 = data_masked[502] | data_masked[366];
  assign data_o[95] = N191 | data_masked[95];
  assign N191 = N190 | data_masked[231];
  assign N190 = data_masked[503] | data_masked[367];
  assign data_o[96] = N193 | data_masked[96];
  assign N193 = N192 | data_masked[232];
  assign N192 = data_masked[504] | data_masked[368];
  assign data_o[97] = N195 | data_masked[97];
  assign N195 = N194 | data_masked[233];
  assign N194 = data_masked[505] | data_masked[369];
  assign data_o[98] = N197 | data_masked[98];
  assign N197 = N196 | data_masked[234];
  assign N196 = data_masked[506] | data_masked[370];
  assign data_o[99] = N199 | data_masked[99];
  assign N199 = N198 | data_masked[235];
  assign N198 = data_masked[507] | data_masked[371];
  assign data_o[100] = N201 | data_masked[100];
  assign N201 = N200 | data_masked[236];
  assign N200 = data_masked[508] | data_masked[372];
  assign data_o[101] = N203 | data_masked[101];
  assign N203 = N202 | data_masked[237];
  assign N202 = data_masked[509] | data_masked[373];
  assign data_o[102] = N205 | data_masked[102];
  assign N205 = N204 | data_masked[238];
  assign N204 = data_masked[510] | data_masked[374];
  assign data_o[103] = N207 | data_masked[103];
  assign N207 = N206 | data_masked[239];
  assign N206 = data_masked[511] | data_masked[375];
  assign data_o[104] = N209 | data_masked[104];
  assign N209 = N208 | data_masked[240];
  assign N208 = data_masked[512] | data_masked[376];
  assign data_o[105] = N211 | data_masked[105];
  assign N211 = N210 | data_masked[241];
  assign N210 = data_masked[513] | data_masked[377];
  assign data_o[106] = N213 | data_masked[106];
  assign N213 = N212 | data_masked[242];
  assign N212 = data_masked[514] | data_masked[378];
  assign data_o[107] = N215 | data_masked[107];
  assign N215 = N214 | data_masked[243];
  assign N214 = data_masked[515] | data_masked[379];
  assign data_o[108] = N217 | data_masked[108];
  assign N217 = N216 | data_masked[244];
  assign N216 = data_masked[516] | data_masked[380];
  assign data_o[109] = N219 | data_masked[109];
  assign N219 = N218 | data_masked[245];
  assign N218 = data_masked[517] | data_masked[381];
  assign data_o[110] = N221 | data_masked[110];
  assign N221 = N220 | data_masked[246];
  assign N220 = data_masked[518] | data_masked[382];
  assign data_o[111] = N223 | data_masked[111];
  assign N223 = N222 | data_masked[247];
  assign N222 = data_masked[519] | data_masked[383];
  assign data_o[112] = N225 | data_masked[112];
  assign N225 = N224 | data_masked[248];
  assign N224 = data_masked[520] | data_masked[384];
  assign data_o[113] = N227 | data_masked[113];
  assign N227 = N226 | data_masked[249];
  assign N226 = data_masked[521] | data_masked[385];
  assign data_o[114] = N229 | data_masked[114];
  assign N229 = N228 | data_masked[250];
  assign N228 = data_masked[522] | data_masked[386];
  assign data_o[115] = N231 | data_masked[115];
  assign N231 = N230 | data_masked[251];
  assign N230 = data_masked[523] | data_masked[387];
  assign data_o[116] = N233 | data_masked[116];
  assign N233 = N232 | data_masked[252];
  assign N232 = data_masked[524] | data_masked[388];
  assign data_o[117] = N235 | data_masked[117];
  assign N235 = N234 | data_masked[253];
  assign N234 = data_masked[525] | data_masked[389];
  assign data_o[118] = N237 | data_masked[118];
  assign N237 = N236 | data_masked[254];
  assign N236 = data_masked[526] | data_masked[390];
  assign data_o[119] = N239 | data_masked[119];
  assign N239 = N238 | data_masked[255];
  assign N238 = data_masked[527] | data_masked[391];
  assign data_o[120] = N241 | data_masked[120];
  assign N241 = N240 | data_masked[256];
  assign N240 = data_masked[528] | data_masked[392];
  assign data_o[121] = N243 | data_masked[121];
  assign N243 = N242 | data_masked[257];
  assign N242 = data_masked[529] | data_masked[393];
  assign data_o[122] = N245 | data_masked[122];
  assign N245 = N244 | data_masked[258];
  assign N244 = data_masked[530] | data_masked[394];
  assign data_o[123] = N247 | data_masked[123];
  assign N247 = N246 | data_masked[259];
  assign N246 = data_masked[531] | data_masked[395];
  assign data_o[124] = N249 | data_masked[124];
  assign N249 = N248 | data_masked[260];
  assign N248 = data_masked[532] | data_masked[396];
  assign data_o[125] = N251 | data_masked[125];
  assign N251 = N250 | data_masked[261];
  assign N250 = data_masked[533] | data_masked[397];
  assign data_o[126] = N253 | data_masked[126];
  assign N253 = N252 | data_masked[262];
  assign N252 = data_masked[534] | data_masked[398];
  assign data_o[127] = N255 | data_masked[127];
  assign N255 = N254 | data_masked[263];
  assign N254 = data_masked[535] | data_masked[399];
  assign data_o[128] = N257 | data_masked[128];
  assign N257 = N256 | data_masked[264];
  assign N256 = data_masked[536] | data_masked[400];
  assign data_o[129] = N259 | data_masked[129];
  assign N259 = N258 | data_masked[265];
  assign N258 = data_masked[537] | data_masked[401];
  assign data_o[130] = N261 | data_masked[130];
  assign N261 = N260 | data_masked[266];
  assign N260 = data_masked[538] | data_masked[402];
  assign data_o[131] = N263 | data_masked[131];
  assign N263 = N262 | data_masked[267];
  assign N262 = data_masked[539] | data_masked[403];
  assign data_o[132] = N265 | data_masked[132];
  assign N265 = N264 | data_masked[268];
  assign N264 = data_masked[540] | data_masked[404];
  assign data_o[133] = N267 | data_masked[133];
  assign N267 = N266 | data_masked[269];
  assign N266 = data_masked[541] | data_masked[405];
  assign data_o[134] = N269 | data_masked[134];
  assign N269 = N268 | data_masked[270];
  assign N268 = data_masked[542] | data_masked[406];
  assign data_o[135] = N271 | data_masked[135];
  assign N271 = N270 | data_masked[271];
  assign N270 = data_masked[543] | data_masked[407];

endmodule



module bsg_mux_one_hot_width_p136_els_p5
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [679:0] data_i;
  input [4:0] sel_one_hot_i;
  output [135:0] data_o;
  wire [135:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407;
  wire [679:0] data_masked;
  assign data_masked[135] = data_i[135] & sel_one_hot_i[0];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[0];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[0];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[0];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[0];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[0];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[0];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[0];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[0];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[0];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[0];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[0];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[0];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[0];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[0];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[0];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[0];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[0];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[0];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[0];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[0];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[0];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[0];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[0];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[0];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[0];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[0];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[0];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[0];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[0];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[0];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[0];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[0];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[0];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[0];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[0];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[0];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[0];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[0];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[0];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[0];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[0];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[0];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[0];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[0];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[0];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[0];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[0];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[0];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[0];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[0];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[0];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[0];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[0];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[0];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[0];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[0];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[0];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[0];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[0];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[0];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[0];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[0];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[0];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[0];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[0];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[0];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[0];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[1];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[1];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[1];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[1];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[1];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[1];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[1];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[1];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[1];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[1];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[1];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[1];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[1];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[1];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[1];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[1];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[1];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[1];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[1];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[1];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[1];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[1];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[1];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[1];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[1];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[1];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[1];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[1];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[1];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[1];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[1];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[1];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[1];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[1];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[1];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[1];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[1];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[1];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[1];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[1];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[1];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[1];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[1];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[1];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[1];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[1];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[1];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[1];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[1];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[1];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[1];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[1];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[1];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[1];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[1];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[1];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[1];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[1];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[1];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[1];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[1];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[1];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[1];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[1];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[1];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[1];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[1];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[1];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[1];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[1];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[1];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[1];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[1];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[1];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[1];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[1];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[1];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[1];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[1];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[1];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[1];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[1];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[1];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[1];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[1];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[1];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[1];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[1];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[1];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[1];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[1];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[1];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[1];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[1];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[1];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[1];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[1];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[1];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[1];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[1];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[1];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[1];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[1];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[1];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[1];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[1];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[1];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[1];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[1];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[1];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[1];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[1];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[1];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[1];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[1];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[1];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[1];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[1];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[1];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[1];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[1];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[1];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[1];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[1];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[1];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[1];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[1];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[1];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[1];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[1];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[1];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[1];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[1];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[1];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[1];
  assign data_masked[407] = data_i[407] & sel_one_hot_i[2];
  assign data_masked[406] = data_i[406] & sel_one_hot_i[2];
  assign data_masked[405] = data_i[405] & sel_one_hot_i[2];
  assign data_masked[404] = data_i[404] & sel_one_hot_i[2];
  assign data_masked[403] = data_i[403] & sel_one_hot_i[2];
  assign data_masked[402] = data_i[402] & sel_one_hot_i[2];
  assign data_masked[401] = data_i[401] & sel_one_hot_i[2];
  assign data_masked[400] = data_i[400] & sel_one_hot_i[2];
  assign data_masked[399] = data_i[399] & sel_one_hot_i[2];
  assign data_masked[398] = data_i[398] & sel_one_hot_i[2];
  assign data_masked[397] = data_i[397] & sel_one_hot_i[2];
  assign data_masked[396] = data_i[396] & sel_one_hot_i[2];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[2];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[2];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[2];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[2];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[2];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[2];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[2];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[2];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[2];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[2];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[2];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[2];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[2];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[2];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[2];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[2];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[2];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[2];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[2];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[2];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[2];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[2];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[2];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[2];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[2];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[2];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[2];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[2];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[2];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[2];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[2];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[2];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[2];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[2];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[2];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[2];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[2];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[2];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[2];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[2];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[2];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[2];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[2];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[2];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[2];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[2];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[2];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[2];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[2];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[2];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[2];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[2];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[2];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[2];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[2];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[2];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[2];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[2];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[2];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[2];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[2];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[2];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[2];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[2];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[2];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[2];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[2];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[2];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[2];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[2];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[2];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[2];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[2];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[2];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[2];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[2];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[2];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[2];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[2];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[2];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[2];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[2];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[2];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[2];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[2];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[2];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[2];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[2];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[2];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[2];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[2];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[2];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[2];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[2];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[2];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[2];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[2];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[2];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[2];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[2];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[2];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[2];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[2];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[2];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[2];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[2];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[2];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[2];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[2];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[2];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[2];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[2];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[2];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[2];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[2];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[2];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[2];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[2];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[2];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[2];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[2];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[2];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[2];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[2];
  assign data_masked[543] = data_i[543] & sel_one_hot_i[3];
  assign data_masked[542] = data_i[542] & sel_one_hot_i[3];
  assign data_masked[541] = data_i[541] & sel_one_hot_i[3];
  assign data_masked[540] = data_i[540] & sel_one_hot_i[3];
  assign data_masked[539] = data_i[539] & sel_one_hot_i[3];
  assign data_masked[538] = data_i[538] & sel_one_hot_i[3];
  assign data_masked[537] = data_i[537] & sel_one_hot_i[3];
  assign data_masked[536] = data_i[536] & sel_one_hot_i[3];
  assign data_masked[535] = data_i[535] & sel_one_hot_i[3];
  assign data_masked[534] = data_i[534] & sel_one_hot_i[3];
  assign data_masked[533] = data_i[533] & sel_one_hot_i[3];
  assign data_masked[532] = data_i[532] & sel_one_hot_i[3];
  assign data_masked[531] = data_i[531] & sel_one_hot_i[3];
  assign data_masked[530] = data_i[530] & sel_one_hot_i[3];
  assign data_masked[529] = data_i[529] & sel_one_hot_i[3];
  assign data_masked[528] = data_i[528] & sel_one_hot_i[3];
  assign data_masked[527] = data_i[527] & sel_one_hot_i[3];
  assign data_masked[526] = data_i[526] & sel_one_hot_i[3];
  assign data_masked[525] = data_i[525] & sel_one_hot_i[3];
  assign data_masked[524] = data_i[524] & sel_one_hot_i[3];
  assign data_masked[523] = data_i[523] & sel_one_hot_i[3];
  assign data_masked[522] = data_i[522] & sel_one_hot_i[3];
  assign data_masked[521] = data_i[521] & sel_one_hot_i[3];
  assign data_masked[520] = data_i[520] & sel_one_hot_i[3];
  assign data_masked[519] = data_i[519] & sel_one_hot_i[3];
  assign data_masked[518] = data_i[518] & sel_one_hot_i[3];
  assign data_masked[517] = data_i[517] & sel_one_hot_i[3];
  assign data_masked[516] = data_i[516] & sel_one_hot_i[3];
  assign data_masked[515] = data_i[515] & sel_one_hot_i[3];
  assign data_masked[514] = data_i[514] & sel_one_hot_i[3];
  assign data_masked[513] = data_i[513] & sel_one_hot_i[3];
  assign data_masked[512] = data_i[512] & sel_one_hot_i[3];
  assign data_masked[511] = data_i[511] & sel_one_hot_i[3];
  assign data_masked[510] = data_i[510] & sel_one_hot_i[3];
  assign data_masked[509] = data_i[509] & sel_one_hot_i[3];
  assign data_masked[508] = data_i[508] & sel_one_hot_i[3];
  assign data_masked[507] = data_i[507] & sel_one_hot_i[3];
  assign data_masked[506] = data_i[506] & sel_one_hot_i[3];
  assign data_masked[505] = data_i[505] & sel_one_hot_i[3];
  assign data_masked[504] = data_i[504] & sel_one_hot_i[3];
  assign data_masked[503] = data_i[503] & sel_one_hot_i[3];
  assign data_masked[502] = data_i[502] & sel_one_hot_i[3];
  assign data_masked[501] = data_i[501] & sel_one_hot_i[3];
  assign data_masked[500] = data_i[500] & sel_one_hot_i[3];
  assign data_masked[499] = data_i[499] & sel_one_hot_i[3];
  assign data_masked[498] = data_i[498] & sel_one_hot_i[3];
  assign data_masked[497] = data_i[497] & sel_one_hot_i[3];
  assign data_masked[496] = data_i[496] & sel_one_hot_i[3];
  assign data_masked[495] = data_i[495] & sel_one_hot_i[3];
  assign data_masked[494] = data_i[494] & sel_one_hot_i[3];
  assign data_masked[493] = data_i[493] & sel_one_hot_i[3];
  assign data_masked[492] = data_i[492] & sel_one_hot_i[3];
  assign data_masked[491] = data_i[491] & sel_one_hot_i[3];
  assign data_masked[490] = data_i[490] & sel_one_hot_i[3];
  assign data_masked[489] = data_i[489] & sel_one_hot_i[3];
  assign data_masked[488] = data_i[488] & sel_one_hot_i[3];
  assign data_masked[487] = data_i[487] & sel_one_hot_i[3];
  assign data_masked[486] = data_i[486] & sel_one_hot_i[3];
  assign data_masked[485] = data_i[485] & sel_one_hot_i[3];
  assign data_masked[484] = data_i[484] & sel_one_hot_i[3];
  assign data_masked[483] = data_i[483] & sel_one_hot_i[3];
  assign data_masked[482] = data_i[482] & sel_one_hot_i[3];
  assign data_masked[481] = data_i[481] & sel_one_hot_i[3];
  assign data_masked[480] = data_i[480] & sel_one_hot_i[3];
  assign data_masked[479] = data_i[479] & sel_one_hot_i[3];
  assign data_masked[478] = data_i[478] & sel_one_hot_i[3];
  assign data_masked[477] = data_i[477] & sel_one_hot_i[3];
  assign data_masked[476] = data_i[476] & sel_one_hot_i[3];
  assign data_masked[475] = data_i[475] & sel_one_hot_i[3];
  assign data_masked[474] = data_i[474] & sel_one_hot_i[3];
  assign data_masked[473] = data_i[473] & sel_one_hot_i[3];
  assign data_masked[472] = data_i[472] & sel_one_hot_i[3];
  assign data_masked[471] = data_i[471] & sel_one_hot_i[3];
  assign data_masked[470] = data_i[470] & sel_one_hot_i[3];
  assign data_masked[469] = data_i[469] & sel_one_hot_i[3];
  assign data_masked[468] = data_i[468] & sel_one_hot_i[3];
  assign data_masked[467] = data_i[467] & sel_one_hot_i[3];
  assign data_masked[466] = data_i[466] & sel_one_hot_i[3];
  assign data_masked[465] = data_i[465] & sel_one_hot_i[3];
  assign data_masked[464] = data_i[464] & sel_one_hot_i[3];
  assign data_masked[463] = data_i[463] & sel_one_hot_i[3];
  assign data_masked[462] = data_i[462] & sel_one_hot_i[3];
  assign data_masked[461] = data_i[461] & sel_one_hot_i[3];
  assign data_masked[460] = data_i[460] & sel_one_hot_i[3];
  assign data_masked[459] = data_i[459] & sel_one_hot_i[3];
  assign data_masked[458] = data_i[458] & sel_one_hot_i[3];
  assign data_masked[457] = data_i[457] & sel_one_hot_i[3];
  assign data_masked[456] = data_i[456] & sel_one_hot_i[3];
  assign data_masked[455] = data_i[455] & sel_one_hot_i[3];
  assign data_masked[454] = data_i[454] & sel_one_hot_i[3];
  assign data_masked[453] = data_i[453] & sel_one_hot_i[3];
  assign data_masked[452] = data_i[452] & sel_one_hot_i[3];
  assign data_masked[451] = data_i[451] & sel_one_hot_i[3];
  assign data_masked[450] = data_i[450] & sel_one_hot_i[3];
  assign data_masked[449] = data_i[449] & sel_one_hot_i[3];
  assign data_masked[448] = data_i[448] & sel_one_hot_i[3];
  assign data_masked[447] = data_i[447] & sel_one_hot_i[3];
  assign data_masked[446] = data_i[446] & sel_one_hot_i[3];
  assign data_masked[445] = data_i[445] & sel_one_hot_i[3];
  assign data_masked[444] = data_i[444] & sel_one_hot_i[3];
  assign data_masked[443] = data_i[443] & sel_one_hot_i[3];
  assign data_masked[442] = data_i[442] & sel_one_hot_i[3];
  assign data_masked[441] = data_i[441] & sel_one_hot_i[3];
  assign data_masked[440] = data_i[440] & sel_one_hot_i[3];
  assign data_masked[439] = data_i[439] & sel_one_hot_i[3];
  assign data_masked[438] = data_i[438] & sel_one_hot_i[3];
  assign data_masked[437] = data_i[437] & sel_one_hot_i[3];
  assign data_masked[436] = data_i[436] & sel_one_hot_i[3];
  assign data_masked[435] = data_i[435] & sel_one_hot_i[3];
  assign data_masked[434] = data_i[434] & sel_one_hot_i[3];
  assign data_masked[433] = data_i[433] & sel_one_hot_i[3];
  assign data_masked[432] = data_i[432] & sel_one_hot_i[3];
  assign data_masked[431] = data_i[431] & sel_one_hot_i[3];
  assign data_masked[430] = data_i[430] & sel_one_hot_i[3];
  assign data_masked[429] = data_i[429] & sel_one_hot_i[3];
  assign data_masked[428] = data_i[428] & sel_one_hot_i[3];
  assign data_masked[427] = data_i[427] & sel_one_hot_i[3];
  assign data_masked[426] = data_i[426] & sel_one_hot_i[3];
  assign data_masked[425] = data_i[425] & sel_one_hot_i[3];
  assign data_masked[424] = data_i[424] & sel_one_hot_i[3];
  assign data_masked[423] = data_i[423] & sel_one_hot_i[3];
  assign data_masked[422] = data_i[422] & sel_one_hot_i[3];
  assign data_masked[421] = data_i[421] & sel_one_hot_i[3];
  assign data_masked[420] = data_i[420] & sel_one_hot_i[3];
  assign data_masked[419] = data_i[419] & sel_one_hot_i[3];
  assign data_masked[418] = data_i[418] & sel_one_hot_i[3];
  assign data_masked[417] = data_i[417] & sel_one_hot_i[3];
  assign data_masked[416] = data_i[416] & sel_one_hot_i[3];
  assign data_masked[415] = data_i[415] & sel_one_hot_i[3];
  assign data_masked[414] = data_i[414] & sel_one_hot_i[3];
  assign data_masked[413] = data_i[413] & sel_one_hot_i[3];
  assign data_masked[412] = data_i[412] & sel_one_hot_i[3];
  assign data_masked[411] = data_i[411] & sel_one_hot_i[3];
  assign data_masked[410] = data_i[410] & sel_one_hot_i[3];
  assign data_masked[409] = data_i[409] & sel_one_hot_i[3];
  assign data_masked[408] = data_i[408] & sel_one_hot_i[3];
  assign data_masked[679] = data_i[679] & sel_one_hot_i[4];
  assign data_masked[678] = data_i[678] & sel_one_hot_i[4];
  assign data_masked[677] = data_i[677] & sel_one_hot_i[4];
  assign data_masked[676] = data_i[676] & sel_one_hot_i[4];
  assign data_masked[675] = data_i[675] & sel_one_hot_i[4];
  assign data_masked[674] = data_i[674] & sel_one_hot_i[4];
  assign data_masked[673] = data_i[673] & sel_one_hot_i[4];
  assign data_masked[672] = data_i[672] & sel_one_hot_i[4];
  assign data_masked[671] = data_i[671] & sel_one_hot_i[4];
  assign data_masked[670] = data_i[670] & sel_one_hot_i[4];
  assign data_masked[669] = data_i[669] & sel_one_hot_i[4];
  assign data_masked[668] = data_i[668] & sel_one_hot_i[4];
  assign data_masked[667] = data_i[667] & sel_one_hot_i[4];
  assign data_masked[666] = data_i[666] & sel_one_hot_i[4];
  assign data_masked[665] = data_i[665] & sel_one_hot_i[4];
  assign data_masked[664] = data_i[664] & sel_one_hot_i[4];
  assign data_masked[663] = data_i[663] & sel_one_hot_i[4];
  assign data_masked[662] = data_i[662] & sel_one_hot_i[4];
  assign data_masked[661] = data_i[661] & sel_one_hot_i[4];
  assign data_masked[660] = data_i[660] & sel_one_hot_i[4];
  assign data_masked[659] = data_i[659] & sel_one_hot_i[4];
  assign data_masked[658] = data_i[658] & sel_one_hot_i[4];
  assign data_masked[657] = data_i[657] & sel_one_hot_i[4];
  assign data_masked[656] = data_i[656] & sel_one_hot_i[4];
  assign data_masked[655] = data_i[655] & sel_one_hot_i[4];
  assign data_masked[654] = data_i[654] & sel_one_hot_i[4];
  assign data_masked[653] = data_i[653] & sel_one_hot_i[4];
  assign data_masked[652] = data_i[652] & sel_one_hot_i[4];
  assign data_masked[651] = data_i[651] & sel_one_hot_i[4];
  assign data_masked[650] = data_i[650] & sel_one_hot_i[4];
  assign data_masked[649] = data_i[649] & sel_one_hot_i[4];
  assign data_masked[648] = data_i[648] & sel_one_hot_i[4];
  assign data_masked[647] = data_i[647] & sel_one_hot_i[4];
  assign data_masked[646] = data_i[646] & sel_one_hot_i[4];
  assign data_masked[645] = data_i[645] & sel_one_hot_i[4];
  assign data_masked[644] = data_i[644] & sel_one_hot_i[4];
  assign data_masked[643] = data_i[643] & sel_one_hot_i[4];
  assign data_masked[642] = data_i[642] & sel_one_hot_i[4];
  assign data_masked[641] = data_i[641] & sel_one_hot_i[4];
  assign data_masked[640] = data_i[640] & sel_one_hot_i[4];
  assign data_masked[639] = data_i[639] & sel_one_hot_i[4];
  assign data_masked[638] = data_i[638] & sel_one_hot_i[4];
  assign data_masked[637] = data_i[637] & sel_one_hot_i[4];
  assign data_masked[636] = data_i[636] & sel_one_hot_i[4];
  assign data_masked[635] = data_i[635] & sel_one_hot_i[4];
  assign data_masked[634] = data_i[634] & sel_one_hot_i[4];
  assign data_masked[633] = data_i[633] & sel_one_hot_i[4];
  assign data_masked[632] = data_i[632] & sel_one_hot_i[4];
  assign data_masked[631] = data_i[631] & sel_one_hot_i[4];
  assign data_masked[630] = data_i[630] & sel_one_hot_i[4];
  assign data_masked[629] = data_i[629] & sel_one_hot_i[4];
  assign data_masked[628] = data_i[628] & sel_one_hot_i[4];
  assign data_masked[627] = data_i[627] & sel_one_hot_i[4];
  assign data_masked[626] = data_i[626] & sel_one_hot_i[4];
  assign data_masked[625] = data_i[625] & sel_one_hot_i[4];
  assign data_masked[624] = data_i[624] & sel_one_hot_i[4];
  assign data_masked[623] = data_i[623] & sel_one_hot_i[4];
  assign data_masked[622] = data_i[622] & sel_one_hot_i[4];
  assign data_masked[621] = data_i[621] & sel_one_hot_i[4];
  assign data_masked[620] = data_i[620] & sel_one_hot_i[4];
  assign data_masked[619] = data_i[619] & sel_one_hot_i[4];
  assign data_masked[618] = data_i[618] & sel_one_hot_i[4];
  assign data_masked[617] = data_i[617] & sel_one_hot_i[4];
  assign data_masked[616] = data_i[616] & sel_one_hot_i[4];
  assign data_masked[615] = data_i[615] & sel_one_hot_i[4];
  assign data_masked[614] = data_i[614] & sel_one_hot_i[4];
  assign data_masked[613] = data_i[613] & sel_one_hot_i[4];
  assign data_masked[612] = data_i[612] & sel_one_hot_i[4];
  assign data_masked[611] = data_i[611] & sel_one_hot_i[4];
  assign data_masked[610] = data_i[610] & sel_one_hot_i[4];
  assign data_masked[609] = data_i[609] & sel_one_hot_i[4];
  assign data_masked[608] = data_i[608] & sel_one_hot_i[4];
  assign data_masked[607] = data_i[607] & sel_one_hot_i[4];
  assign data_masked[606] = data_i[606] & sel_one_hot_i[4];
  assign data_masked[605] = data_i[605] & sel_one_hot_i[4];
  assign data_masked[604] = data_i[604] & sel_one_hot_i[4];
  assign data_masked[603] = data_i[603] & sel_one_hot_i[4];
  assign data_masked[602] = data_i[602] & sel_one_hot_i[4];
  assign data_masked[601] = data_i[601] & sel_one_hot_i[4];
  assign data_masked[600] = data_i[600] & sel_one_hot_i[4];
  assign data_masked[599] = data_i[599] & sel_one_hot_i[4];
  assign data_masked[598] = data_i[598] & sel_one_hot_i[4];
  assign data_masked[597] = data_i[597] & sel_one_hot_i[4];
  assign data_masked[596] = data_i[596] & sel_one_hot_i[4];
  assign data_masked[595] = data_i[595] & sel_one_hot_i[4];
  assign data_masked[594] = data_i[594] & sel_one_hot_i[4];
  assign data_masked[593] = data_i[593] & sel_one_hot_i[4];
  assign data_masked[592] = data_i[592] & sel_one_hot_i[4];
  assign data_masked[591] = data_i[591] & sel_one_hot_i[4];
  assign data_masked[590] = data_i[590] & sel_one_hot_i[4];
  assign data_masked[589] = data_i[589] & sel_one_hot_i[4];
  assign data_masked[588] = data_i[588] & sel_one_hot_i[4];
  assign data_masked[587] = data_i[587] & sel_one_hot_i[4];
  assign data_masked[586] = data_i[586] & sel_one_hot_i[4];
  assign data_masked[585] = data_i[585] & sel_one_hot_i[4];
  assign data_masked[584] = data_i[584] & sel_one_hot_i[4];
  assign data_masked[583] = data_i[583] & sel_one_hot_i[4];
  assign data_masked[582] = data_i[582] & sel_one_hot_i[4];
  assign data_masked[581] = data_i[581] & sel_one_hot_i[4];
  assign data_masked[580] = data_i[580] & sel_one_hot_i[4];
  assign data_masked[579] = data_i[579] & sel_one_hot_i[4];
  assign data_masked[578] = data_i[578] & sel_one_hot_i[4];
  assign data_masked[577] = data_i[577] & sel_one_hot_i[4];
  assign data_masked[576] = data_i[576] & sel_one_hot_i[4];
  assign data_masked[575] = data_i[575] & sel_one_hot_i[4];
  assign data_masked[574] = data_i[574] & sel_one_hot_i[4];
  assign data_masked[573] = data_i[573] & sel_one_hot_i[4];
  assign data_masked[572] = data_i[572] & sel_one_hot_i[4];
  assign data_masked[571] = data_i[571] & sel_one_hot_i[4];
  assign data_masked[570] = data_i[570] & sel_one_hot_i[4];
  assign data_masked[569] = data_i[569] & sel_one_hot_i[4];
  assign data_masked[568] = data_i[568] & sel_one_hot_i[4];
  assign data_masked[567] = data_i[567] & sel_one_hot_i[4];
  assign data_masked[566] = data_i[566] & sel_one_hot_i[4];
  assign data_masked[565] = data_i[565] & sel_one_hot_i[4];
  assign data_masked[564] = data_i[564] & sel_one_hot_i[4];
  assign data_masked[563] = data_i[563] & sel_one_hot_i[4];
  assign data_masked[562] = data_i[562] & sel_one_hot_i[4];
  assign data_masked[561] = data_i[561] & sel_one_hot_i[4];
  assign data_masked[560] = data_i[560] & sel_one_hot_i[4];
  assign data_masked[559] = data_i[559] & sel_one_hot_i[4];
  assign data_masked[558] = data_i[558] & sel_one_hot_i[4];
  assign data_masked[557] = data_i[557] & sel_one_hot_i[4];
  assign data_masked[556] = data_i[556] & sel_one_hot_i[4];
  assign data_masked[555] = data_i[555] & sel_one_hot_i[4];
  assign data_masked[554] = data_i[554] & sel_one_hot_i[4];
  assign data_masked[553] = data_i[553] & sel_one_hot_i[4];
  assign data_masked[552] = data_i[552] & sel_one_hot_i[4];
  assign data_masked[551] = data_i[551] & sel_one_hot_i[4];
  assign data_masked[550] = data_i[550] & sel_one_hot_i[4];
  assign data_masked[549] = data_i[549] & sel_one_hot_i[4];
  assign data_masked[548] = data_i[548] & sel_one_hot_i[4];
  assign data_masked[547] = data_i[547] & sel_one_hot_i[4];
  assign data_masked[546] = data_i[546] & sel_one_hot_i[4];
  assign data_masked[545] = data_i[545] & sel_one_hot_i[4];
  assign data_masked[544] = data_i[544] & sel_one_hot_i[4];
  assign data_o[0] = N2 | data_masked[0];
  assign N2 = N1 | data_masked[136];
  assign N1 = N0 | data_masked[272];
  assign N0 = data_masked[544] | data_masked[408];
  assign data_o[1] = N5 | data_masked[1];
  assign N5 = N4 | data_masked[137];
  assign N4 = N3 | data_masked[273];
  assign N3 = data_masked[545] | data_masked[409];
  assign data_o[2] = N8 | data_masked[2];
  assign N8 = N7 | data_masked[138];
  assign N7 = N6 | data_masked[274];
  assign N6 = data_masked[546] | data_masked[410];
  assign data_o[3] = N11 | data_masked[3];
  assign N11 = N10 | data_masked[139];
  assign N10 = N9 | data_masked[275];
  assign N9 = data_masked[547] | data_masked[411];
  assign data_o[4] = N14 | data_masked[4];
  assign N14 = N13 | data_masked[140];
  assign N13 = N12 | data_masked[276];
  assign N12 = data_masked[548] | data_masked[412];
  assign data_o[5] = N17 | data_masked[5];
  assign N17 = N16 | data_masked[141];
  assign N16 = N15 | data_masked[277];
  assign N15 = data_masked[549] | data_masked[413];
  assign data_o[6] = N20 | data_masked[6];
  assign N20 = N19 | data_masked[142];
  assign N19 = N18 | data_masked[278];
  assign N18 = data_masked[550] | data_masked[414];
  assign data_o[7] = N23 | data_masked[7];
  assign N23 = N22 | data_masked[143];
  assign N22 = N21 | data_masked[279];
  assign N21 = data_masked[551] | data_masked[415];
  assign data_o[8] = N26 | data_masked[8];
  assign N26 = N25 | data_masked[144];
  assign N25 = N24 | data_masked[280];
  assign N24 = data_masked[552] | data_masked[416];
  assign data_o[9] = N29 | data_masked[9];
  assign N29 = N28 | data_masked[145];
  assign N28 = N27 | data_masked[281];
  assign N27 = data_masked[553] | data_masked[417];
  assign data_o[10] = N32 | data_masked[10];
  assign N32 = N31 | data_masked[146];
  assign N31 = N30 | data_masked[282];
  assign N30 = data_masked[554] | data_masked[418];
  assign data_o[11] = N35 | data_masked[11];
  assign N35 = N34 | data_masked[147];
  assign N34 = N33 | data_masked[283];
  assign N33 = data_masked[555] | data_masked[419];
  assign data_o[12] = N38 | data_masked[12];
  assign N38 = N37 | data_masked[148];
  assign N37 = N36 | data_masked[284];
  assign N36 = data_masked[556] | data_masked[420];
  assign data_o[13] = N41 | data_masked[13];
  assign N41 = N40 | data_masked[149];
  assign N40 = N39 | data_masked[285];
  assign N39 = data_masked[557] | data_masked[421];
  assign data_o[14] = N44 | data_masked[14];
  assign N44 = N43 | data_masked[150];
  assign N43 = N42 | data_masked[286];
  assign N42 = data_masked[558] | data_masked[422];
  assign data_o[15] = N47 | data_masked[15];
  assign N47 = N46 | data_masked[151];
  assign N46 = N45 | data_masked[287];
  assign N45 = data_masked[559] | data_masked[423];
  assign data_o[16] = N50 | data_masked[16];
  assign N50 = N49 | data_masked[152];
  assign N49 = N48 | data_masked[288];
  assign N48 = data_masked[560] | data_masked[424];
  assign data_o[17] = N53 | data_masked[17];
  assign N53 = N52 | data_masked[153];
  assign N52 = N51 | data_masked[289];
  assign N51 = data_masked[561] | data_masked[425];
  assign data_o[18] = N56 | data_masked[18];
  assign N56 = N55 | data_masked[154];
  assign N55 = N54 | data_masked[290];
  assign N54 = data_masked[562] | data_masked[426];
  assign data_o[19] = N59 | data_masked[19];
  assign N59 = N58 | data_masked[155];
  assign N58 = N57 | data_masked[291];
  assign N57 = data_masked[563] | data_masked[427];
  assign data_o[20] = N62 | data_masked[20];
  assign N62 = N61 | data_masked[156];
  assign N61 = N60 | data_masked[292];
  assign N60 = data_masked[564] | data_masked[428];
  assign data_o[21] = N65 | data_masked[21];
  assign N65 = N64 | data_masked[157];
  assign N64 = N63 | data_masked[293];
  assign N63 = data_masked[565] | data_masked[429];
  assign data_o[22] = N68 | data_masked[22];
  assign N68 = N67 | data_masked[158];
  assign N67 = N66 | data_masked[294];
  assign N66 = data_masked[566] | data_masked[430];
  assign data_o[23] = N71 | data_masked[23];
  assign N71 = N70 | data_masked[159];
  assign N70 = N69 | data_masked[295];
  assign N69 = data_masked[567] | data_masked[431];
  assign data_o[24] = N74 | data_masked[24];
  assign N74 = N73 | data_masked[160];
  assign N73 = N72 | data_masked[296];
  assign N72 = data_masked[568] | data_masked[432];
  assign data_o[25] = N77 | data_masked[25];
  assign N77 = N76 | data_masked[161];
  assign N76 = N75 | data_masked[297];
  assign N75 = data_masked[569] | data_masked[433];
  assign data_o[26] = N80 | data_masked[26];
  assign N80 = N79 | data_masked[162];
  assign N79 = N78 | data_masked[298];
  assign N78 = data_masked[570] | data_masked[434];
  assign data_o[27] = N83 | data_masked[27];
  assign N83 = N82 | data_masked[163];
  assign N82 = N81 | data_masked[299];
  assign N81 = data_masked[571] | data_masked[435];
  assign data_o[28] = N86 | data_masked[28];
  assign N86 = N85 | data_masked[164];
  assign N85 = N84 | data_masked[300];
  assign N84 = data_masked[572] | data_masked[436];
  assign data_o[29] = N89 | data_masked[29];
  assign N89 = N88 | data_masked[165];
  assign N88 = N87 | data_masked[301];
  assign N87 = data_masked[573] | data_masked[437];
  assign data_o[30] = N92 | data_masked[30];
  assign N92 = N91 | data_masked[166];
  assign N91 = N90 | data_masked[302];
  assign N90 = data_masked[574] | data_masked[438];
  assign data_o[31] = N95 | data_masked[31];
  assign N95 = N94 | data_masked[167];
  assign N94 = N93 | data_masked[303];
  assign N93 = data_masked[575] | data_masked[439];
  assign data_o[32] = N98 | data_masked[32];
  assign N98 = N97 | data_masked[168];
  assign N97 = N96 | data_masked[304];
  assign N96 = data_masked[576] | data_masked[440];
  assign data_o[33] = N101 | data_masked[33];
  assign N101 = N100 | data_masked[169];
  assign N100 = N99 | data_masked[305];
  assign N99 = data_masked[577] | data_masked[441];
  assign data_o[34] = N104 | data_masked[34];
  assign N104 = N103 | data_masked[170];
  assign N103 = N102 | data_masked[306];
  assign N102 = data_masked[578] | data_masked[442];
  assign data_o[35] = N107 | data_masked[35];
  assign N107 = N106 | data_masked[171];
  assign N106 = N105 | data_masked[307];
  assign N105 = data_masked[579] | data_masked[443];
  assign data_o[36] = N110 | data_masked[36];
  assign N110 = N109 | data_masked[172];
  assign N109 = N108 | data_masked[308];
  assign N108 = data_masked[580] | data_masked[444];
  assign data_o[37] = N113 | data_masked[37];
  assign N113 = N112 | data_masked[173];
  assign N112 = N111 | data_masked[309];
  assign N111 = data_masked[581] | data_masked[445];
  assign data_o[38] = N116 | data_masked[38];
  assign N116 = N115 | data_masked[174];
  assign N115 = N114 | data_masked[310];
  assign N114 = data_masked[582] | data_masked[446];
  assign data_o[39] = N119 | data_masked[39];
  assign N119 = N118 | data_masked[175];
  assign N118 = N117 | data_masked[311];
  assign N117 = data_masked[583] | data_masked[447];
  assign data_o[40] = N122 | data_masked[40];
  assign N122 = N121 | data_masked[176];
  assign N121 = N120 | data_masked[312];
  assign N120 = data_masked[584] | data_masked[448];
  assign data_o[41] = N125 | data_masked[41];
  assign N125 = N124 | data_masked[177];
  assign N124 = N123 | data_masked[313];
  assign N123 = data_masked[585] | data_masked[449];
  assign data_o[42] = N128 | data_masked[42];
  assign N128 = N127 | data_masked[178];
  assign N127 = N126 | data_masked[314];
  assign N126 = data_masked[586] | data_masked[450];
  assign data_o[43] = N131 | data_masked[43];
  assign N131 = N130 | data_masked[179];
  assign N130 = N129 | data_masked[315];
  assign N129 = data_masked[587] | data_masked[451];
  assign data_o[44] = N134 | data_masked[44];
  assign N134 = N133 | data_masked[180];
  assign N133 = N132 | data_masked[316];
  assign N132 = data_masked[588] | data_masked[452];
  assign data_o[45] = N137 | data_masked[45];
  assign N137 = N136 | data_masked[181];
  assign N136 = N135 | data_masked[317];
  assign N135 = data_masked[589] | data_masked[453];
  assign data_o[46] = N140 | data_masked[46];
  assign N140 = N139 | data_masked[182];
  assign N139 = N138 | data_masked[318];
  assign N138 = data_masked[590] | data_masked[454];
  assign data_o[47] = N143 | data_masked[47];
  assign N143 = N142 | data_masked[183];
  assign N142 = N141 | data_masked[319];
  assign N141 = data_masked[591] | data_masked[455];
  assign data_o[48] = N146 | data_masked[48];
  assign N146 = N145 | data_masked[184];
  assign N145 = N144 | data_masked[320];
  assign N144 = data_masked[592] | data_masked[456];
  assign data_o[49] = N149 | data_masked[49];
  assign N149 = N148 | data_masked[185];
  assign N148 = N147 | data_masked[321];
  assign N147 = data_masked[593] | data_masked[457];
  assign data_o[50] = N152 | data_masked[50];
  assign N152 = N151 | data_masked[186];
  assign N151 = N150 | data_masked[322];
  assign N150 = data_masked[594] | data_masked[458];
  assign data_o[51] = N155 | data_masked[51];
  assign N155 = N154 | data_masked[187];
  assign N154 = N153 | data_masked[323];
  assign N153 = data_masked[595] | data_masked[459];
  assign data_o[52] = N158 | data_masked[52];
  assign N158 = N157 | data_masked[188];
  assign N157 = N156 | data_masked[324];
  assign N156 = data_masked[596] | data_masked[460];
  assign data_o[53] = N161 | data_masked[53];
  assign N161 = N160 | data_masked[189];
  assign N160 = N159 | data_masked[325];
  assign N159 = data_masked[597] | data_masked[461];
  assign data_o[54] = N164 | data_masked[54];
  assign N164 = N163 | data_masked[190];
  assign N163 = N162 | data_masked[326];
  assign N162 = data_masked[598] | data_masked[462];
  assign data_o[55] = N167 | data_masked[55];
  assign N167 = N166 | data_masked[191];
  assign N166 = N165 | data_masked[327];
  assign N165 = data_masked[599] | data_masked[463];
  assign data_o[56] = N170 | data_masked[56];
  assign N170 = N169 | data_masked[192];
  assign N169 = N168 | data_masked[328];
  assign N168 = data_masked[600] | data_masked[464];
  assign data_o[57] = N173 | data_masked[57];
  assign N173 = N172 | data_masked[193];
  assign N172 = N171 | data_masked[329];
  assign N171 = data_masked[601] | data_masked[465];
  assign data_o[58] = N176 | data_masked[58];
  assign N176 = N175 | data_masked[194];
  assign N175 = N174 | data_masked[330];
  assign N174 = data_masked[602] | data_masked[466];
  assign data_o[59] = N179 | data_masked[59];
  assign N179 = N178 | data_masked[195];
  assign N178 = N177 | data_masked[331];
  assign N177 = data_masked[603] | data_masked[467];
  assign data_o[60] = N182 | data_masked[60];
  assign N182 = N181 | data_masked[196];
  assign N181 = N180 | data_masked[332];
  assign N180 = data_masked[604] | data_masked[468];
  assign data_o[61] = N185 | data_masked[61];
  assign N185 = N184 | data_masked[197];
  assign N184 = N183 | data_masked[333];
  assign N183 = data_masked[605] | data_masked[469];
  assign data_o[62] = N188 | data_masked[62];
  assign N188 = N187 | data_masked[198];
  assign N187 = N186 | data_masked[334];
  assign N186 = data_masked[606] | data_masked[470];
  assign data_o[63] = N191 | data_masked[63];
  assign N191 = N190 | data_masked[199];
  assign N190 = N189 | data_masked[335];
  assign N189 = data_masked[607] | data_masked[471];
  assign data_o[64] = N194 | data_masked[64];
  assign N194 = N193 | data_masked[200];
  assign N193 = N192 | data_masked[336];
  assign N192 = data_masked[608] | data_masked[472];
  assign data_o[65] = N197 | data_masked[65];
  assign N197 = N196 | data_masked[201];
  assign N196 = N195 | data_masked[337];
  assign N195 = data_masked[609] | data_masked[473];
  assign data_o[66] = N200 | data_masked[66];
  assign N200 = N199 | data_masked[202];
  assign N199 = N198 | data_masked[338];
  assign N198 = data_masked[610] | data_masked[474];
  assign data_o[67] = N203 | data_masked[67];
  assign N203 = N202 | data_masked[203];
  assign N202 = N201 | data_masked[339];
  assign N201 = data_masked[611] | data_masked[475];
  assign data_o[68] = N206 | data_masked[68];
  assign N206 = N205 | data_masked[204];
  assign N205 = N204 | data_masked[340];
  assign N204 = data_masked[612] | data_masked[476];
  assign data_o[69] = N209 | data_masked[69];
  assign N209 = N208 | data_masked[205];
  assign N208 = N207 | data_masked[341];
  assign N207 = data_masked[613] | data_masked[477];
  assign data_o[70] = N212 | data_masked[70];
  assign N212 = N211 | data_masked[206];
  assign N211 = N210 | data_masked[342];
  assign N210 = data_masked[614] | data_masked[478];
  assign data_o[71] = N215 | data_masked[71];
  assign N215 = N214 | data_masked[207];
  assign N214 = N213 | data_masked[343];
  assign N213 = data_masked[615] | data_masked[479];
  assign data_o[72] = N218 | data_masked[72];
  assign N218 = N217 | data_masked[208];
  assign N217 = N216 | data_masked[344];
  assign N216 = data_masked[616] | data_masked[480];
  assign data_o[73] = N221 | data_masked[73];
  assign N221 = N220 | data_masked[209];
  assign N220 = N219 | data_masked[345];
  assign N219 = data_masked[617] | data_masked[481];
  assign data_o[74] = N224 | data_masked[74];
  assign N224 = N223 | data_masked[210];
  assign N223 = N222 | data_masked[346];
  assign N222 = data_masked[618] | data_masked[482];
  assign data_o[75] = N227 | data_masked[75];
  assign N227 = N226 | data_masked[211];
  assign N226 = N225 | data_masked[347];
  assign N225 = data_masked[619] | data_masked[483];
  assign data_o[76] = N230 | data_masked[76];
  assign N230 = N229 | data_masked[212];
  assign N229 = N228 | data_masked[348];
  assign N228 = data_masked[620] | data_masked[484];
  assign data_o[77] = N233 | data_masked[77];
  assign N233 = N232 | data_masked[213];
  assign N232 = N231 | data_masked[349];
  assign N231 = data_masked[621] | data_masked[485];
  assign data_o[78] = N236 | data_masked[78];
  assign N236 = N235 | data_masked[214];
  assign N235 = N234 | data_masked[350];
  assign N234 = data_masked[622] | data_masked[486];
  assign data_o[79] = N239 | data_masked[79];
  assign N239 = N238 | data_masked[215];
  assign N238 = N237 | data_masked[351];
  assign N237 = data_masked[623] | data_masked[487];
  assign data_o[80] = N242 | data_masked[80];
  assign N242 = N241 | data_masked[216];
  assign N241 = N240 | data_masked[352];
  assign N240 = data_masked[624] | data_masked[488];
  assign data_o[81] = N245 | data_masked[81];
  assign N245 = N244 | data_masked[217];
  assign N244 = N243 | data_masked[353];
  assign N243 = data_masked[625] | data_masked[489];
  assign data_o[82] = N248 | data_masked[82];
  assign N248 = N247 | data_masked[218];
  assign N247 = N246 | data_masked[354];
  assign N246 = data_masked[626] | data_masked[490];
  assign data_o[83] = N251 | data_masked[83];
  assign N251 = N250 | data_masked[219];
  assign N250 = N249 | data_masked[355];
  assign N249 = data_masked[627] | data_masked[491];
  assign data_o[84] = N254 | data_masked[84];
  assign N254 = N253 | data_masked[220];
  assign N253 = N252 | data_masked[356];
  assign N252 = data_masked[628] | data_masked[492];
  assign data_o[85] = N257 | data_masked[85];
  assign N257 = N256 | data_masked[221];
  assign N256 = N255 | data_masked[357];
  assign N255 = data_masked[629] | data_masked[493];
  assign data_o[86] = N260 | data_masked[86];
  assign N260 = N259 | data_masked[222];
  assign N259 = N258 | data_masked[358];
  assign N258 = data_masked[630] | data_masked[494];
  assign data_o[87] = N263 | data_masked[87];
  assign N263 = N262 | data_masked[223];
  assign N262 = N261 | data_masked[359];
  assign N261 = data_masked[631] | data_masked[495];
  assign data_o[88] = N266 | data_masked[88];
  assign N266 = N265 | data_masked[224];
  assign N265 = N264 | data_masked[360];
  assign N264 = data_masked[632] | data_masked[496];
  assign data_o[89] = N269 | data_masked[89];
  assign N269 = N268 | data_masked[225];
  assign N268 = N267 | data_masked[361];
  assign N267 = data_masked[633] | data_masked[497];
  assign data_o[90] = N272 | data_masked[90];
  assign N272 = N271 | data_masked[226];
  assign N271 = N270 | data_masked[362];
  assign N270 = data_masked[634] | data_masked[498];
  assign data_o[91] = N275 | data_masked[91];
  assign N275 = N274 | data_masked[227];
  assign N274 = N273 | data_masked[363];
  assign N273 = data_masked[635] | data_masked[499];
  assign data_o[92] = N278 | data_masked[92];
  assign N278 = N277 | data_masked[228];
  assign N277 = N276 | data_masked[364];
  assign N276 = data_masked[636] | data_masked[500];
  assign data_o[93] = N281 | data_masked[93];
  assign N281 = N280 | data_masked[229];
  assign N280 = N279 | data_masked[365];
  assign N279 = data_masked[637] | data_masked[501];
  assign data_o[94] = N284 | data_masked[94];
  assign N284 = N283 | data_masked[230];
  assign N283 = N282 | data_masked[366];
  assign N282 = data_masked[638] | data_masked[502];
  assign data_o[95] = N287 | data_masked[95];
  assign N287 = N286 | data_masked[231];
  assign N286 = N285 | data_masked[367];
  assign N285 = data_masked[639] | data_masked[503];
  assign data_o[96] = N290 | data_masked[96];
  assign N290 = N289 | data_masked[232];
  assign N289 = N288 | data_masked[368];
  assign N288 = data_masked[640] | data_masked[504];
  assign data_o[97] = N293 | data_masked[97];
  assign N293 = N292 | data_masked[233];
  assign N292 = N291 | data_masked[369];
  assign N291 = data_masked[641] | data_masked[505];
  assign data_o[98] = N296 | data_masked[98];
  assign N296 = N295 | data_masked[234];
  assign N295 = N294 | data_masked[370];
  assign N294 = data_masked[642] | data_masked[506];
  assign data_o[99] = N299 | data_masked[99];
  assign N299 = N298 | data_masked[235];
  assign N298 = N297 | data_masked[371];
  assign N297 = data_masked[643] | data_masked[507];
  assign data_o[100] = N302 | data_masked[100];
  assign N302 = N301 | data_masked[236];
  assign N301 = N300 | data_masked[372];
  assign N300 = data_masked[644] | data_masked[508];
  assign data_o[101] = N305 | data_masked[101];
  assign N305 = N304 | data_masked[237];
  assign N304 = N303 | data_masked[373];
  assign N303 = data_masked[645] | data_masked[509];
  assign data_o[102] = N308 | data_masked[102];
  assign N308 = N307 | data_masked[238];
  assign N307 = N306 | data_masked[374];
  assign N306 = data_masked[646] | data_masked[510];
  assign data_o[103] = N311 | data_masked[103];
  assign N311 = N310 | data_masked[239];
  assign N310 = N309 | data_masked[375];
  assign N309 = data_masked[647] | data_masked[511];
  assign data_o[104] = N314 | data_masked[104];
  assign N314 = N313 | data_masked[240];
  assign N313 = N312 | data_masked[376];
  assign N312 = data_masked[648] | data_masked[512];
  assign data_o[105] = N317 | data_masked[105];
  assign N317 = N316 | data_masked[241];
  assign N316 = N315 | data_masked[377];
  assign N315 = data_masked[649] | data_masked[513];
  assign data_o[106] = N320 | data_masked[106];
  assign N320 = N319 | data_masked[242];
  assign N319 = N318 | data_masked[378];
  assign N318 = data_masked[650] | data_masked[514];
  assign data_o[107] = N323 | data_masked[107];
  assign N323 = N322 | data_masked[243];
  assign N322 = N321 | data_masked[379];
  assign N321 = data_masked[651] | data_masked[515];
  assign data_o[108] = N326 | data_masked[108];
  assign N326 = N325 | data_masked[244];
  assign N325 = N324 | data_masked[380];
  assign N324 = data_masked[652] | data_masked[516];
  assign data_o[109] = N329 | data_masked[109];
  assign N329 = N328 | data_masked[245];
  assign N328 = N327 | data_masked[381];
  assign N327 = data_masked[653] | data_masked[517];
  assign data_o[110] = N332 | data_masked[110];
  assign N332 = N331 | data_masked[246];
  assign N331 = N330 | data_masked[382];
  assign N330 = data_masked[654] | data_masked[518];
  assign data_o[111] = N335 | data_masked[111];
  assign N335 = N334 | data_masked[247];
  assign N334 = N333 | data_masked[383];
  assign N333 = data_masked[655] | data_masked[519];
  assign data_o[112] = N338 | data_masked[112];
  assign N338 = N337 | data_masked[248];
  assign N337 = N336 | data_masked[384];
  assign N336 = data_masked[656] | data_masked[520];
  assign data_o[113] = N341 | data_masked[113];
  assign N341 = N340 | data_masked[249];
  assign N340 = N339 | data_masked[385];
  assign N339 = data_masked[657] | data_masked[521];
  assign data_o[114] = N344 | data_masked[114];
  assign N344 = N343 | data_masked[250];
  assign N343 = N342 | data_masked[386];
  assign N342 = data_masked[658] | data_masked[522];
  assign data_o[115] = N347 | data_masked[115];
  assign N347 = N346 | data_masked[251];
  assign N346 = N345 | data_masked[387];
  assign N345 = data_masked[659] | data_masked[523];
  assign data_o[116] = N350 | data_masked[116];
  assign N350 = N349 | data_masked[252];
  assign N349 = N348 | data_masked[388];
  assign N348 = data_masked[660] | data_masked[524];
  assign data_o[117] = N353 | data_masked[117];
  assign N353 = N352 | data_masked[253];
  assign N352 = N351 | data_masked[389];
  assign N351 = data_masked[661] | data_masked[525];
  assign data_o[118] = N356 | data_masked[118];
  assign N356 = N355 | data_masked[254];
  assign N355 = N354 | data_masked[390];
  assign N354 = data_masked[662] | data_masked[526];
  assign data_o[119] = N359 | data_masked[119];
  assign N359 = N358 | data_masked[255];
  assign N358 = N357 | data_masked[391];
  assign N357 = data_masked[663] | data_masked[527];
  assign data_o[120] = N362 | data_masked[120];
  assign N362 = N361 | data_masked[256];
  assign N361 = N360 | data_masked[392];
  assign N360 = data_masked[664] | data_masked[528];
  assign data_o[121] = N365 | data_masked[121];
  assign N365 = N364 | data_masked[257];
  assign N364 = N363 | data_masked[393];
  assign N363 = data_masked[665] | data_masked[529];
  assign data_o[122] = N368 | data_masked[122];
  assign N368 = N367 | data_masked[258];
  assign N367 = N366 | data_masked[394];
  assign N366 = data_masked[666] | data_masked[530];
  assign data_o[123] = N371 | data_masked[123];
  assign N371 = N370 | data_masked[259];
  assign N370 = N369 | data_masked[395];
  assign N369 = data_masked[667] | data_masked[531];
  assign data_o[124] = N374 | data_masked[124];
  assign N374 = N373 | data_masked[260];
  assign N373 = N372 | data_masked[396];
  assign N372 = data_masked[668] | data_masked[532];
  assign data_o[125] = N377 | data_masked[125];
  assign N377 = N376 | data_masked[261];
  assign N376 = N375 | data_masked[397];
  assign N375 = data_masked[669] | data_masked[533];
  assign data_o[126] = N380 | data_masked[126];
  assign N380 = N379 | data_masked[262];
  assign N379 = N378 | data_masked[398];
  assign N378 = data_masked[670] | data_masked[534];
  assign data_o[127] = N383 | data_masked[127];
  assign N383 = N382 | data_masked[263];
  assign N382 = N381 | data_masked[399];
  assign N381 = data_masked[671] | data_masked[535];
  assign data_o[128] = N386 | data_masked[128];
  assign N386 = N385 | data_masked[264];
  assign N385 = N384 | data_masked[400];
  assign N384 = data_masked[672] | data_masked[536];
  assign data_o[129] = N389 | data_masked[129];
  assign N389 = N388 | data_masked[265];
  assign N388 = N387 | data_masked[401];
  assign N387 = data_masked[673] | data_masked[537];
  assign data_o[130] = N392 | data_masked[130];
  assign N392 = N391 | data_masked[266];
  assign N391 = N390 | data_masked[402];
  assign N390 = data_masked[674] | data_masked[538];
  assign data_o[131] = N395 | data_masked[131];
  assign N395 = N394 | data_masked[267];
  assign N394 = N393 | data_masked[403];
  assign N393 = data_masked[675] | data_masked[539];
  assign data_o[132] = N398 | data_masked[132];
  assign N398 = N397 | data_masked[268];
  assign N397 = N396 | data_masked[404];
  assign N396 = data_masked[676] | data_masked[540];
  assign data_o[133] = N401 | data_masked[133];
  assign N401 = N400 | data_masked[269];
  assign N400 = N399 | data_masked[405];
  assign N399 = data_masked[677] | data_masked[541];
  assign data_o[134] = N404 | data_masked[134];
  assign N404 = N403 | data_masked[270];
  assign N403 = N402 | data_masked[406];
  assign N402 = data_masked[678] | data_masked[542];
  assign data_o[135] = N407 | data_masked[135];
  assign N407 = N406 | data_masked[271];
  assign N406 = N405 | data_masked[407];
  assign N405 = data_masked[679] | data_masked[543];

endmodule



module bsg_wormhole_router_136_1_1_2_1_1_1_00000013_0000001a
(
  clk_i,
  reset_i,
  local_x_cord_i,
  local_y_cord_i,
  valid_i,
  data_i,
  ready_o,
  valid_o,
  data_o,
  ready_i
);

  input [0:0] local_x_cord_i;
  input [0:0] local_y_cord_i;
  input [4:0] valid_i;
  input [679:0] data_i;
  output [4:0] ready_o;
  output [4:0] valid_o;
  output [679:0] data_o;
  input [4:0] ready_i;
  input clk_i;
  input reset_i;
  wire [4:0] ready_o,valid_o,fifo_yumi_i;
  wire [679:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,fifo_data_o_3__135_,fifo_data_o_3__134_,fifo_data_o_3__133_,
  fifo_data_o_3__132_,fifo_data_o_3__131_,fifo_data_o_3__130_,fifo_data_o_3__129_,
  fifo_data_o_3__128_,fifo_data_o_3__127_,fifo_data_o_3__126_,fifo_data_o_3__125_,
  fifo_data_o_3__124_,fifo_data_o_3__123_,fifo_data_o_3__122_,fifo_data_o_3__121_,
  fifo_data_o_3__120_,fifo_data_o_3__119_,fifo_data_o_3__118_,fifo_data_o_3__117_,
  fifo_data_o_3__116_,fifo_data_o_3__115_,fifo_data_o_3__114_,fifo_data_o_3__113_,
  fifo_data_o_3__112_,fifo_data_o_3__111_,fifo_data_o_3__110_,fifo_data_o_3__109_,
  fifo_data_o_3__108_,fifo_data_o_3__107_,fifo_data_o_3__106_,fifo_data_o_3__105_,
  fifo_data_o_3__104_,fifo_data_o_3__103_,fifo_data_o_3__102_,fifo_data_o_3__101_,
  fifo_data_o_3__100_,fifo_data_o_3__99_,fifo_data_o_3__98_,fifo_data_o_3__97_,
  fifo_data_o_3__96_,fifo_data_o_3__95_,fifo_data_o_3__94_,fifo_data_o_3__93_,
  fifo_data_o_3__92_,fifo_data_o_3__91_,fifo_data_o_3__90_,fifo_data_o_3__89_,fifo_data_o_3__88_,
  fifo_data_o_3__87_,fifo_data_o_3__86_,fifo_data_o_3__85_,fifo_data_o_3__84_,
  fifo_data_o_3__83_,fifo_data_o_3__82_,fifo_data_o_3__81_,fifo_data_o_3__80_,
  fifo_data_o_3__79_,fifo_data_o_3__78_,fifo_data_o_3__77_,fifo_data_o_3__76_,
  fifo_data_o_3__75_,fifo_data_o_3__74_,fifo_data_o_3__73_,fifo_data_o_3__72_,
  fifo_data_o_3__71_,fifo_data_o_3__70_,fifo_data_o_3__69_,fifo_data_o_3__68_,fifo_data_o_3__67_,
  fifo_data_o_3__66_,fifo_data_o_3__65_,fifo_data_o_3__64_,fifo_data_o_3__63_,
  fifo_data_o_3__62_,fifo_data_o_3__61_,fifo_data_o_3__60_,fifo_data_o_3__59_,
  fifo_data_o_3__58_,fifo_data_o_3__57_,fifo_data_o_3__56_,fifo_data_o_3__55_,
  fifo_data_o_3__54_,fifo_data_o_3__53_,fifo_data_o_3__52_,fifo_data_o_3__51_,fifo_data_o_3__50_,
  fifo_data_o_3__49_,fifo_data_o_3__48_,fifo_data_o_3__47_,fifo_data_o_3__46_,
  fifo_data_o_3__45_,fifo_data_o_3__44_,fifo_data_o_3__43_,fifo_data_o_3__42_,
  fifo_data_o_3__41_,fifo_data_o_3__40_,fifo_data_o_3__39_,fifo_data_o_3__38_,
  fifo_data_o_3__37_,fifo_data_o_3__36_,fifo_data_o_3__35_,fifo_data_o_3__34_,
  fifo_data_o_3__33_,fifo_data_o_3__32_,fifo_data_o_3__31_,fifo_data_o_3__30_,fifo_data_o_3__29_,
  fifo_data_o_3__28_,fifo_data_o_3__27_,fifo_data_o_3__26_,fifo_data_o_3__25_,
  fifo_data_o_3__24_,fifo_data_o_3__23_,fifo_data_o_3__22_,fifo_data_o_3__21_,
  fifo_data_o_3__20_,fifo_data_o_3__19_,fifo_data_o_3__18_,fifo_data_o_3__17_,
  fifo_data_o_3__16_,fifo_data_o_3__15_,fifo_data_o_3__14_,fifo_data_o_3__13_,
  fifo_data_o_3__12_,fifo_data_o_3__11_,fifo_data_o_3__10_,fifo_data_o_3__9_,fifo_data_o_3__8_,
  fifo_data_o_3__7_,fifo_data_o_3__6_,fifo_data_o_3__5_,fifo_data_o_3__4_,
  fifo_data_o_3__3_,fifo_data_o_3__2_,fifo_data_o_3__1_,fifo_data_o_3__0_,fifo_data_o_2__135_,
  fifo_data_o_2__134_,fifo_data_o_2__133_,fifo_data_o_2__132_,fifo_data_o_2__131_,
  fifo_data_o_2__130_,fifo_data_o_2__129_,fifo_data_o_2__128_,fifo_data_o_2__127_,
  fifo_data_o_2__126_,fifo_data_o_2__125_,fifo_data_o_2__124_,fifo_data_o_2__123_,
  fifo_data_o_2__122_,fifo_data_o_2__121_,fifo_data_o_2__120_,fifo_data_o_2__119_,
  fifo_data_o_2__118_,fifo_data_o_2__117_,fifo_data_o_2__116_,fifo_data_o_2__115_,
  fifo_data_o_2__114_,fifo_data_o_2__113_,fifo_data_o_2__112_,fifo_data_o_2__111_,
  fifo_data_o_2__110_,fifo_data_o_2__109_,fifo_data_o_2__108_,fifo_data_o_2__107_,
  fifo_data_o_2__106_,fifo_data_o_2__105_,fifo_data_o_2__104_,fifo_data_o_2__103_,
  fifo_data_o_2__102_,fifo_data_o_2__101_,fifo_data_o_2__100_,fifo_data_o_2__99_,
  fifo_data_o_2__98_,fifo_data_o_2__97_,fifo_data_o_2__96_,fifo_data_o_2__95_,
  fifo_data_o_2__94_,fifo_data_o_2__93_,fifo_data_o_2__92_,fifo_data_o_2__91_,
  fifo_data_o_2__90_,fifo_data_o_2__89_,fifo_data_o_2__88_,fifo_data_o_2__87_,
  fifo_data_o_2__86_,fifo_data_o_2__85_,fifo_data_o_2__84_,fifo_data_o_2__83_,
  fifo_data_o_2__82_,fifo_data_o_2__81_,fifo_data_o_2__80_,fifo_data_o_2__79_,fifo_data_o_2__78_,
  fifo_data_o_2__77_,fifo_data_o_2__76_,fifo_data_o_2__75_,fifo_data_o_2__74_,
  fifo_data_o_2__73_,fifo_data_o_2__72_,fifo_data_o_2__71_,fifo_data_o_2__70_,
  fifo_data_o_2__69_,fifo_data_o_2__68_,fifo_data_o_2__67_,fifo_data_o_2__66_,
  fifo_data_o_2__65_,fifo_data_o_2__64_,fifo_data_o_2__63_,fifo_data_o_2__62_,
  fifo_data_o_2__61_,fifo_data_o_2__60_,fifo_data_o_2__59_,fifo_data_o_2__58_,fifo_data_o_2__57_,
  fifo_data_o_2__56_,fifo_data_o_2__55_,fifo_data_o_2__54_,fifo_data_o_2__53_,
  fifo_data_o_2__52_,fifo_data_o_2__51_,fifo_data_o_2__50_,fifo_data_o_2__49_,
  fifo_data_o_2__48_,fifo_data_o_2__47_,fifo_data_o_2__46_,fifo_data_o_2__45_,
  fifo_data_o_2__44_,fifo_data_o_2__43_,fifo_data_o_2__42_,fifo_data_o_2__41_,fifo_data_o_2__40_,
  fifo_data_o_2__39_,fifo_data_o_2__38_,fifo_data_o_2__37_,fifo_data_o_2__36_,
  fifo_data_o_2__35_,fifo_data_o_2__34_,fifo_data_o_2__33_,fifo_data_o_2__32_,
  fifo_data_o_2__31_,fifo_data_o_2__30_,fifo_data_o_2__29_,fifo_data_o_2__28_,
  fifo_data_o_2__27_,fifo_data_o_2__26_,fifo_data_o_2__25_,fifo_data_o_2__24_,
  fifo_data_o_2__23_,fifo_data_o_2__22_,fifo_data_o_2__21_,fifo_data_o_2__20_,fifo_data_o_2__19_,
  fifo_data_o_2__18_,fifo_data_o_2__17_,fifo_data_o_2__16_,fifo_data_o_2__15_,
  fifo_data_o_2__14_,fifo_data_o_2__13_,fifo_data_o_2__12_,fifo_data_o_2__11_,
  fifo_data_o_2__10_,fifo_data_o_2__9_,fifo_data_o_2__8_,fifo_data_o_2__7_,
  fifo_data_o_2__6_,fifo_data_o_2__5_,fifo_data_o_2__4_,fifo_data_o_2__3_,fifo_data_o_2__2_,
  fifo_data_o_2__1_,fifo_data_o_2__0_,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,
  N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,
  N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,
  N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,
  N178,N179,N180,N181,N182,N183,N184,N185,N186,dest_n_4__3_,dest_n_4__2_,
  dest_n_4__1_,dest_n_4__0_,dest_n_3__4_,dest_n_3__2_,dest_n_3__1_,dest_n_3__0_,
  dest_n_2__4_,dest_n_2__3_,dest_n_2__1_,dest_n_2__0_,dest_n_1__4_,dest_n_1__3_,dest_n_1__2_,
  dest_n_1__0_,dest_n_0__4_,dest_n_0__3_,dest_n_0__2_,dest_n_0__1_,dest_n_0__0_,
  new_valid_4__3_,new_valid_4__2_,new_valid_4__1_,new_valid_4__0_,new_valid_3__4_,
  new_valid_3__2_,new_valid_3__1_,new_valid_3__0_,new_valid_2__4_,new_valid_2__3_,
  new_valid_2__1_,new_valid_2__0_,new_valid_1__4_,new_valid_1__3_,new_valid_1__2_,
  new_valid_1__0_,new_valid_0__4_,new_valid_0__3_,new_valid_0__2_,new_valid_0__1_,
  new_valid_0__0_,arb_grants_o_4__3_,arb_grants_o_4__2_,arb_grants_o_4__1_,
  arb_grants_o_4__0_,arb_grants_o_3__4_,arb_grants_o_3__2_,arb_grants_o_3__1_,
  arb_grants_o_3__0_,arb_grants_o_2__4_,arb_grants_o_2__3_,arb_grants_o_2__1_,
  arb_grants_o_2__0_,arb_grants_o_1__4_,arb_grants_o_1__3_,arb_grants_o_1__2_,arb_grants_o_1__0_,
  arb_grants_o_0__4_,arb_grants_o_0__3_,arb_grants_o_0__2_,arb_grants_o_0__1_,
  arb_grants_o_0__0_,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,
  N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,
  N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,
  N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,
  N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,arb_valid_4__3_,arb_valid_4__2_,
  arb_valid_4__1_,arb_valid_4__0_,arb_valid_3__4_,arb_valid_3__2_,arb_valid_3__1_,
  arb_valid_3__0_,arb_valid_2__4_,arb_valid_2__3_,arb_valid_2__1_,arb_valid_2__0_,
  arb_valid_1__4_,arb_valid_1__3_,arb_valid_1__2_,arb_valid_1__0_,arb_valid_0__4_,
  arb_valid_0__3_,arb_valid_0__2_,arb_valid_0__1_,arb_valid_0__0_,N258,N259,N260,
  N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,
  N277,n_3_net_,arb_sel_o_4__3_,arb_sel_o_4__2_,arb_sel_o_4__1_,arb_sel_o_4__0_,
  arb_sel_o_3__3_,arb_sel_o_3__2_,arb_sel_o_3__1_,arb_sel_o_3__0_,arb_sel_o_2__3_,
  arb_sel_o_2__2_,arb_sel_o_2__1_,arb_sel_o_2__0_,arb_sel_o_1__3_,arb_sel_o_1__2_,
  arb_sel_o_1__1_,arb_sel_o_1__0_,arb_sel_o_0__4_,arb_sel_o_0__3_,arb_sel_o_0__2_,
  arb_sel_o_0__1_,arb_sel_o_0__0_,n_9_net_,n_15_net_,n_21_net_,n_27_net_,N278,N279,
  N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,
  N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,
  N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,
  N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
  N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,
  N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,
  N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,
  N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,
  N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,
  N424,N425,N426,N427,N428,N429,N430,N431,N432,SV2V_UNCONNECTED_1,
  SV2V_UNCONNECTED_2,SV2V_UNCONNECTED_3,SV2V_UNCONNECTED_4,SV2V_UNCONNECTED_5,
  SV2V_UNCONNECTED_6,SV2V_UNCONNECTED_7,SV2V_UNCONNECTED_8,
  SV2V_UNCONNECTED_9,SV2V_UNCONNECTED_10,SV2V_UNCONNECTED_11;
  wire [3:2] fifo_valid_o;
  reg [9:0] count_r,out_count_r;
  reg dest_r_0__4_,dest_r_0__3_,dest_r_0__2_,dest_r_0__1_,dest_r_0__0_,dest_r_1__4_,
  dest_r_1__3_,dest_r_1__2_,dest_r_1__0_,dest_r_2__4_,dest_r_2__3_,dest_r_2__1_,
  dest_r_2__0_,dest_r_3__4_,dest_r_3__2_,dest_r_3__1_,dest_r_3__0_,dest_r_4__3_,
  dest_r_4__2_,dest_r_4__1_,dest_r_4__0_,arb_grants_r_0__0_,arb_grants_r_0__1_,
  arb_grants_r_0__2_,arb_grants_r_0__3_,arb_grants_r_0__4_,arb_grants_r_1__0_,
  arb_grants_r_1__2_,arb_grants_r_1__3_,arb_grants_r_1__4_,arb_grants_r_2__0_,
  arb_grants_r_2__1_,arb_grants_r_2__3_,arb_grants_r_2__4_,arb_grants_r_3__0_,arb_grants_r_3__1_,
  arb_grants_r_3__2_,arb_grants_r_3__4_,arb_grants_r_4__0_,arb_grants_r_4__1_,
  arb_grants_r_4__2_,arb_grants_r_4__3_;
  assign ready_o[4] = 1'b1;
  assign ready_o[1] = 1'b1;
  assign ready_o[0] = 1'b1;

  bsg_two_fifo_width_p136
  in_ff_2__no_stub_two_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(ready_o[2]),
    .data_i(data_i[407:272]),
    .v_i(valid_i[2]),
    .v_o(fifo_valid_o[2]),
    .data_o({ fifo_data_o_2__135_, fifo_data_o_2__134_, fifo_data_o_2__133_, fifo_data_o_2__132_, fifo_data_o_2__131_, fifo_data_o_2__130_, fifo_data_o_2__129_, fifo_data_o_2__128_, fifo_data_o_2__127_, fifo_data_o_2__126_, fifo_data_o_2__125_, fifo_data_o_2__124_, fifo_data_o_2__123_, fifo_data_o_2__122_, fifo_data_o_2__121_, fifo_data_o_2__120_, fifo_data_o_2__119_, fifo_data_o_2__118_, fifo_data_o_2__117_, fifo_data_o_2__116_, fifo_data_o_2__115_, fifo_data_o_2__114_, fifo_data_o_2__113_, fifo_data_o_2__112_, fifo_data_o_2__111_, fifo_data_o_2__110_, fifo_data_o_2__109_, fifo_data_o_2__108_, fifo_data_o_2__107_, fifo_data_o_2__106_, fifo_data_o_2__105_, fifo_data_o_2__104_, fifo_data_o_2__103_, fifo_data_o_2__102_, fifo_data_o_2__101_, fifo_data_o_2__100_, fifo_data_o_2__99_, fifo_data_o_2__98_, fifo_data_o_2__97_, fifo_data_o_2__96_, fifo_data_o_2__95_, fifo_data_o_2__94_, fifo_data_o_2__93_, fifo_data_o_2__92_, fifo_data_o_2__91_, fifo_data_o_2__90_, fifo_data_o_2__89_, fifo_data_o_2__88_, fifo_data_o_2__87_, fifo_data_o_2__86_, fifo_data_o_2__85_, fifo_data_o_2__84_, fifo_data_o_2__83_, fifo_data_o_2__82_, fifo_data_o_2__81_, fifo_data_o_2__80_, fifo_data_o_2__79_, fifo_data_o_2__78_, fifo_data_o_2__77_, fifo_data_o_2__76_, fifo_data_o_2__75_, fifo_data_o_2__74_, fifo_data_o_2__73_, fifo_data_o_2__72_, fifo_data_o_2__71_, fifo_data_o_2__70_, fifo_data_o_2__69_, fifo_data_o_2__68_, fifo_data_o_2__67_, fifo_data_o_2__66_, fifo_data_o_2__65_, fifo_data_o_2__64_, fifo_data_o_2__63_, fifo_data_o_2__62_, fifo_data_o_2__61_, fifo_data_o_2__60_, fifo_data_o_2__59_, fifo_data_o_2__58_, fifo_data_o_2__57_, fifo_data_o_2__56_, fifo_data_o_2__55_, fifo_data_o_2__54_, fifo_data_o_2__53_, fifo_data_o_2__52_, fifo_data_o_2__51_, fifo_data_o_2__50_, fifo_data_o_2__49_, fifo_data_o_2__48_, fifo_data_o_2__47_, fifo_data_o_2__46_, fifo_data_o_2__45_, fifo_data_o_2__44_, fifo_data_o_2__43_, fifo_data_o_2__42_, fifo_data_o_2__41_, fifo_data_o_2__40_, fifo_data_o_2__39_, fifo_data_o_2__38_, fifo_data_o_2__37_, fifo_data_o_2__36_, fifo_data_o_2__35_, fifo_data_o_2__34_, fifo_data_o_2__33_, fifo_data_o_2__32_, fifo_data_o_2__31_, fifo_data_o_2__30_, fifo_data_o_2__29_, fifo_data_o_2__28_, fifo_data_o_2__27_, fifo_data_o_2__26_, fifo_data_o_2__25_, fifo_data_o_2__24_, fifo_data_o_2__23_, fifo_data_o_2__22_, fifo_data_o_2__21_, fifo_data_o_2__20_, fifo_data_o_2__19_, fifo_data_o_2__18_, fifo_data_o_2__17_, fifo_data_o_2__16_, fifo_data_o_2__15_, fifo_data_o_2__14_, fifo_data_o_2__13_, fifo_data_o_2__12_, fifo_data_o_2__11_, fifo_data_o_2__10_, fifo_data_o_2__9_, fifo_data_o_2__8_, fifo_data_o_2__7_, fifo_data_o_2__6_, fifo_data_o_2__5_, fifo_data_o_2__4_, fifo_data_o_2__3_, fifo_data_o_2__2_, fifo_data_o_2__1_, fifo_data_o_2__0_ }),
    .yumi_i(fifo_yumi_i[2])
  );


  bsg_two_fifo_width_p136
  in_ff_3__no_stub_two_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(ready_o[3]),
    .data_i(data_i[543:408]),
    .v_i(valid_i[3]),
    .v_o(fifo_valid_o[3]),
    .data_o({ fifo_data_o_3__135_, fifo_data_o_3__134_, fifo_data_o_3__133_, fifo_data_o_3__132_, fifo_data_o_3__131_, fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_ }),
    .yumi_i(fifo_yumi_i[3])
  );


  bsg_round_robin_arb_inputs_p4
  out_side_1__rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ arb_valid_4__1_, arb_valid_3__1_, arb_valid_2__1_, arb_valid_0__1_ }),
    .grants_o({ arb_grants_o_4__1_, arb_grants_o_3__1_, arb_grants_o_2__1_, arb_grants_o_0__1_ }),
    .sel_one_hot_o({ arb_sel_o_1__3_, arb_sel_o_1__2_, arb_sel_o_1__1_, arb_sel_o_1__0_ }),
    .v_o(valid_o[1]),
    .tag_o({ SV2V_UNCONNECTED_1, SV2V_UNCONNECTED_2 }),
    .yumi_i(n_3_net_)
  );


  bsg_mux_one_hot_width_p136_els_p4
  out_side_1__mux
  (
    .data_i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_o_3__135_, fifo_data_o_3__134_, fifo_data_o_3__133_, fifo_data_o_3__132_, fifo_data_o_3__131_, fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_, fifo_data_o_2__135_, fifo_data_o_2__134_, fifo_data_o_2__133_, fifo_data_o_2__132_, fifo_data_o_2__131_, fifo_data_o_2__130_, fifo_data_o_2__129_, fifo_data_o_2__128_, fifo_data_o_2__127_, fifo_data_o_2__126_, fifo_data_o_2__125_, fifo_data_o_2__124_, fifo_data_o_2__123_, fifo_data_o_2__122_, fifo_data_o_2__121_, fifo_data_o_2__120_, fifo_data_o_2__119_, fifo_data_o_2__118_, fifo_data_o_2__117_, fifo_data_o_2__116_, fifo_data_o_2__115_, fifo_data_o_2__114_, fifo_data_o_2__113_, fifo_data_o_2__112_, fifo_data_o_2__111_, fifo_data_o_2__110_, fifo_data_o_2__109_, fifo_data_o_2__108_, fifo_data_o_2__107_, fifo_data_o_2__106_, fifo_data_o_2__105_, fifo_data_o_2__104_, fifo_data_o_2__103_, fifo_data_o_2__102_, fifo_data_o_2__101_, fifo_data_o_2__100_, fifo_data_o_2__99_, fifo_data_o_2__98_, fifo_data_o_2__97_, fifo_data_o_2__96_, fifo_data_o_2__95_, fifo_data_o_2__94_, fifo_data_o_2__93_, fifo_data_o_2__92_, fifo_data_o_2__91_, fifo_data_o_2__90_, fifo_data_o_2__89_, fifo_data_o_2__88_, fifo_data_o_2__87_, fifo_data_o_2__86_, fifo_data_o_2__85_, fifo_data_o_2__84_, fifo_data_o_2__83_, fifo_data_o_2__82_, fifo_data_o_2__81_, fifo_data_o_2__80_, fifo_data_o_2__79_, fifo_data_o_2__78_, fifo_data_o_2__77_, fifo_data_o_2__76_, fifo_data_o_2__75_, fifo_data_o_2__74_, fifo_data_o_2__73_, fifo_data_o_2__72_, fifo_data_o_2__71_, fifo_data_o_2__70_, fifo_data_o_2__69_, fifo_data_o_2__68_, fifo_data_o_2__67_, fifo_data_o_2__66_, fifo_data_o_2__65_, fifo_data_o_2__64_, fifo_data_o_2__63_, fifo_data_o_2__62_, fifo_data_o_2__61_, fifo_data_o_2__60_, fifo_data_o_2__59_, fifo_data_o_2__58_, fifo_data_o_2__57_, fifo_data_o_2__56_, fifo_data_o_2__55_, fifo_data_o_2__54_, fifo_data_o_2__53_, fifo_data_o_2__52_, fifo_data_o_2__51_, fifo_data_o_2__50_, fifo_data_o_2__49_, fifo_data_o_2__48_, fifo_data_o_2__47_, fifo_data_o_2__46_, fifo_data_o_2__45_, fifo_data_o_2__44_, fifo_data_o_2__43_, fifo_data_o_2__42_, fifo_data_o_2__41_, fifo_data_o_2__40_, fifo_data_o_2__39_, fifo_data_o_2__38_, fifo_data_o_2__37_, fifo_data_o_2__36_, fifo_data_o_2__35_, fifo_data_o_2__34_, fifo_data_o_2__33_, fifo_data_o_2__32_, fifo_data_o_2__31_, fifo_data_o_2__30_, fifo_data_o_2__29_, fifo_data_o_2__28_, fifo_data_o_2__27_, fifo_data_o_2__26_, fifo_data_o_2__25_, fifo_data_o_2__24_, fifo_data_o_2__23_, fifo_data_o_2__22_, fifo_data_o_2__21_, fifo_data_o_2__20_, fifo_data_o_2__19_, fifo_data_o_2__18_, fifo_data_o_2__17_, fifo_data_o_2__16_, fifo_data_o_2__15_, fifo_data_o_2__14_, fifo_data_o_2__13_, fifo_data_o_2__12_, fifo_data_o_2__11_, fifo_data_o_2__10_, fifo_data_o_2__9_, fifo_data_o_2__8_, fifo_data_o_2__7_, fifo_data_o_2__6_, fifo_data_o_2__5_, fifo_data_o_2__4_, fifo_data_o_2__3_, fifo_data_o_2__2_, fifo_data_o_2__1_, fifo_data_o_2__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_1__3_, arb_sel_o_1__2_, arb_sel_o_1__1_, arb_sel_o_1__0_ }),
    .data_o(data_o[271:136])
  );


  bsg_round_robin_arb_inputs_p4
  out_side_2__rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[2]),
    .reqs_i({ arb_valid_4__2_, arb_valid_3__2_, arb_valid_1__2_, arb_valid_0__2_ }),
    .grants_o({ arb_grants_o_4__2_, arb_grants_o_3__2_, arb_grants_o_1__2_, arb_grants_o_0__2_ }),
    .sel_one_hot_o({ arb_sel_o_2__3_, arb_sel_o_2__2_, arb_sel_o_2__1_, arb_sel_o_2__0_ }),
    .v_o(valid_o[2]),
    .tag_o({ SV2V_UNCONNECTED_3, SV2V_UNCONNECTED_4 }),
    .yumi_i(n_9_net_)
  );


  bsg_mux_one_hot_width_p136_els_p4
  out_side_2__mux
  (
    .data_i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_o_3__135_, fifo_data_o_3__134_, fifo_data_o_3__133_, fifo_data_o_3__132_, fifo_data_o_3__131_, fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_2__3_, arb_sel_o_2__2_, arb_sel_o_2__1_, arb_sel_o_2__0_ }),
    .data_o(data_o[407:272])
  );


  bsg_round_robin_arb_inputs_p4
  out_side_3__rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ arb_valid_4__3_, arb_valid_2__3_, arb_valid_1__3_, arb_valid_0__3_ }),
    .grants_o({ arb_grants_o_4__3_, arb_grants_o_2__3_, arb_grants_o_1__3_, arb_grants_o_0__3_ }),
    .sel_one_hot_o({ arb_sel_o_3__3_, arb_sel_o_3__2_, arb_sel_o_3__1_, arb_sel_o_3__0_ }),
    .v_o(valid_o[3]),
    .tag_o({ SV2V_UNCONNECTED_5, SV2V_UNCONNECTED_6 }),
    .yumi_i(n_15_net_)
  );


  bsg_mux_one_hot_width_p136_els_p4
  out_side_3__mux
  (
    .data_i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_o_2__135_, fifo_data_o_2__134_, fifo_data_o_2__133_, fifo_data_o_2__132_, fifo_data_o_2__131_, fifo_data_o_2__130_, fifo_data_o_2__129_, fifo_data_o_2__128_, fifo_data_o_2__127_, fifo_data_o_2__126_, fifo_data_o_2__125_, fifo_data_o_2__124_, fifo_data_o_2__123_, fifo_data_o_2__122_, fifo_data_o_2__121_, fifo_data_o_2__120_, fifo_data_o_2__119_, fifo_data_o_2__118_, fifo_data_o_2__117_, fifo_data_o_2__116_, fifo_data_o_2__115_, fifo_data_o_2__114_, fifo_data_o_2__113_, fifo_data_o_2__112_, fifo_data_o_2__111_, fifo_data_o_2__110_, fifo_data_o_2__109_, fifo_data_o_2__108_, fifo_data_o_2__107_, fifo_data_o_2__106_, fifo_data_o_2__105_, fifo_data_o_2__104_, fifo_data_o_2__103_, fifo_data_o_2__102_, fifo_data_o_2__101_, fifo_data_o_2__100_, fifo_data_o_2__99_, fifo_data_o_2__98_, fifo_data_o_2__97_, fifo_data_o_2__96_, fifo_data_o_2__95_, fifo_data_o_2__94_, fifo_data_o_2__93_, fifo_data_o_2__92_, fifo_data_o_2__91_, fifo_data_o_2__90_, fifo_data_o_2__89_, fifo_data_o_2__88_, fifo_data_o_2__87_, fifo_data_o_2__86_, fifo_data_o_2__85_, fifo_data_o_2__84_, fifo_data_o_2__83_, fifo_data_o_2__82_, fifo_data_o_2__81_, fifo_data_o_2__80_, fifo_data_o_2__79_, fifo_data_o_2__78_, fifo_data_o_2__77_, fifo_data_o_2__76_, fifo_data_o_2__75_, fifo_data_o_2__74_, fifo_data_o_2__73_, fifo_data_o_2__72_, fifo_data_o_2__71_, fifo_data_o_2__70_, fifo_data_o_2__69_, fifo_data_o_2__68_, fifo_data_o_2__67_, fifo_data_o_2__66_, fifo_data_o_2__65_, fifo_data_o_2__64_, fifo_data_o_2__63_, fifo_data_o_2__62_, fifo_data_o_2__61_, fifo_data_o_2__60_, fifo_data_o_2__59_, fifo_data_o_2__58_, fifo_data_o_2__57_, fifo_data_o_2__56_, fifo_data_o_2__55_, fifo_data_o_2__54_, fifo_data_o_2__53_, fifo_data_o_2__52_, fifo_data_o_2__51_, fifo_data_o_2__50_, fifo_data_o_2__49_, fifo_data_o_2__48_, fifo_data_o_2__47_, fifo_data_o_2__46_, fifo_data_o_2__45_, fifo_data_o_2__44_, fifo_data_o_2__43_, fifo_data_o_2__42_, fifo_data_o_2__41_, fifo_data_o_2__40_, fifo_data_o_2__39_, fifo_data_o_2__38_, fifo_data_o_2__37_, fifo_data_o_2__36_, fifo_data_o_2__35_, fifo_data_o_2__34_, fifo_data_o_2__33_, fifo_data_o_2__32_, fifo_data_o_2__31_, fifo_data_o_2__30_, fifo_data_o_2__29_, fifo_data_o_2__28_, fifo_data_o_2__27_, fifo_data_o_2__26_, fifo_data_o_2__25_, fifo_data_o_2__24_, fifo_data_o_2__23_, fifo_data_o_2__22_, fifo_data_o_2__21_, fifo_data_o_2__20_, fifo_data_o_2__19_, fifo_data_o_2__18_, fifo_data_o_2__17_, fifo_data_o_2__16_, fifo_data_o_2__15_, fifo_data_o_2__14_, fifo_data_o_2__13_, fifo_data_o_2__12_, fifo_data_o_2__11_, fifo_data_o_2__10_, fifo_data_o_2__9_, fifo_data_o_2__8_, fifo_data_o_2__7_, fifo_data_o_2__6_, fifo_data_o_2__5_, fifo_data_o_2__4_, fifo_data_o_2__3_, fifo_data_o_2__2_, fifo_data_o_2__1_, fifo_data_o_2__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_3__3_, arb_sel_o_3__2_, arb_sel_o_3__1_, arb_sel_o_3__0_ }),
    .data_o(data_o[543:408])
  );


  bsg_round_robin_arb_inputs_p4
  out_side_4__rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ arb_valid_3__4_, arb_valid_2__4_, arb_valid_1__4_, arb_valid_0__4_ }),
    .grants_o({ arb_grants_o_3__4_, arb_grants_o_2__4_, arb_grants_o_1__4_, arb_grants_o_0__4_ }),
    .sel_one_hot_o({ arb_sel_o_4__3_, arb_sel_o_4__2_, arb_sel_o_4__1_, arb_sel_o_4__0_ }),
    .v_o(valid_o[4]),
    .tag_o({ SV2V_UNCONNECTED_7, SV2V_UNCONNECTED_8 }),
    .yumi_i(n_21_net_)
  );


  bsg_mux_one_hot_width_p136_els_p4
  out_side_4__mux
  (
    .data_i({ fifo_data_o_3__135_, fifo_data_o_3__134_, fifo_data_o_3__133_, fifo_data_o_3__132_, fifo_data_o_3__131_, fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_, fifo_data_o_2__135_, fifo_data_o_2__134_, fifo_data_o_2__133_, fifo_data_o_2__132_, fifo_data_o_2__131_, fifo_data_o_2__130_, fifo_data_o_2__129_, fifo_data_o_2__128_, fifo_data_o_2__127_, fifo_data_o_2__126_, fifo_data_o_2__125_, fifo_data_o_2__124_, fifo_data_o_2__123_, fifo_data_o_2__122_, fifo_data_o_2__121_, fifo_data_o_2__120_, fifo_data_o_2__119_, fifo_data_o_2__118_, fifo_data_o_2__117_, fifo_data_o_2__116_, fifo_data_o_2__115_, fifo_data_o_2__114_, fifo_data_o_2__113_, fifo_data_o_2__112_, fifo_data_o_2__111_, fifo_data_o_2__110_, fifo_data_o_2__109_, fifo_data_o_2__108_, fifo_data_o_2__107_, fifo_data_o_2__106_, fifo_data_o_2__105_, fifo_data_o_2__104_, fifo_data_o_2__103_, fifo_data_o_2__102_, fifo_data_o_2__101_, fifo_data_o_2__100_, fifo_data_o_2__99_, fifo_data_o_2__98_, fifo_data_o_2__97_, fifo_data_o_2__96_, fifo_data_o_2__95_, fifo_data_o_2__94_, fifo_data_o_2__93_, fifo_data_o_2__92_, fifo_data_o_2__91_, fifo_data_o_2__90_, fifo_data_o_2__89_, fifo_data_o_2__88_, fifo_data_o_2__87_, fifo_data_o_2__86_, fifo_data_o_2__85_, fifo_data_o_2__84_, fifo_data_o_2__83_, fifo_data_o_2__82_, fifo_data_o_2__81_, fifo_data_o_2__80_, fifo_data_o_2__79_, fifo_data_o_2__78_, fifo_data_o_2__77_, fifo_data_o_2__76_, fifo_data_o_2__75_, fifo_data_o_2__74_, fifo_data_o_2__73_, fifo_data_o_2__72_, fifo_data_o_2__71_, fifo_data_o_2__70_, fifo_data_o_2__69_, fifo_data_o_2__68_, fifo_data_o_2__67_, fifo_data_o_2__66_, fifo_data_o_2__65_, fifo_data_o_2__64_, fifo_data_o_2__63_, fifo_data_o_2__62_, fifo_data_o_2__61_, fifo_data_o_2__60_, fifo_data_o_2__59_, fifo_data_o_2__58_, fifo_data_o_2__57_, fifo_data_o_2__56_, fifo_data_o_2__55_, fifo_data_o_2__54_, fifo_data_o_2__53_, fifo_data_o_2__52_, fifo_data_o_2__51_, fifo_data_o_2__50_, fifo_data_o_2__49_, fifo_data_o_2__48_, fifo_data_o_2__47_, fifo_data_o_2__46_, fifo_data_o_2__45_, fifo_data_o_2__44_, fifo_data_o_2__43_, fifo_data_o_2__42_, fifo_data_o_2__41_, fifo_data_o_2__40_, fifo_data_o_2__39_, fifo_data_o_2__38_, fifo_data_o_2__37_, fifo_data_o_2__36_, fifo_data_o_2__35_, fifo_data_o_2__34_, fifo_data_o_2__33_, fifo_data_o_2__32_, fifo_data_o_2__31_, fifo_data_o_2__30_, fifo_data_o_2__29_, fifo_data_o_2__28_, fifo_data_o_2__27_, fifo_data_o_2__26_, fifo_data_o_2__25_, fifo_data_o_2__24_, fifo_data_o_2__23_, fifo_data_o_2__22_, fifo_data_o_2__21_, fifo_data_o_2__20_, fifo_data_o_2__19_, fifo_data_o_2__18_, fifo_data_o_2__17_, fifo_data_o_2__16_, fifo_data_o_2__15_, fifo_data_o_2__14_, fifo_data_o_2__13_, fifo_data_o_2__12_, fifo_data_o_2__11_, fifo_data_o_2__10_, fifo_data_o_2__9_, fifo_data_o_2__8_, fifo_data_o_2__7_, fifo_data_o_2__6_, fifo_data_o_2__5_, fifo_data_o_2__4_, fifo_data_o_2__3_, fifo_data_o_2__2_, fifo_data_o_2__1_, fifo_data_o_2__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_4__3_, arb_sel_o_4__2_, arb_sel_o_4__1_, arb_sel_o_4__0_ }),
    .data_o(data_o[679:544])
  );


  bsg_round_robin_arb_inputs_p5
  rr_arb_proc
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[0]),
    .reqs_i({ arb_valid_4__0_, arb_valid_3__0_, arb_valid_2__0_, arb_valid_1__0_, arb_valid_0__0_ }),
    .grants_o({ arb_grants_o_4__0_, arb_grants_o_3__0_, arb_grants_o_2__0_, arb_grants_o_1__0_, arb_grants_o_0__0_ }),
    .sel_one_hot_o({ arb_sel_o_0__4_, arb_sel_o_0__3_, arb_sel_o_0__2_, arb_sel_o_0__1_, arb_sel_o_0__0_ }),
    .v_o(valid_o[0]),
    .tag_o({ SV2V_UNCONNECTED_9, SV2V_UNCONNECTED_10, SV2V_UNCONNECTED_11 }),
    .yumi_i(n_27_net_)
  );


  bsg_mux_one_hot_width_p136_els_p5
  mux_proc
  (
    .data_i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_o_3__135_, fifo_data_o_3__134_, fifo_data_o_3__133_, fifo_data_o_3__132_, fifo_data_o_3__131_, fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_, fifo_data_o_2__135_, fifo_data_o_2__134_, fifo_data_o_2__133_, fifo_data_o_2__132_, fifo_data_o_2__131_, fifo_data_o_2__130_, fifo_data_o_2__129_, fifo_data_o_2__128_, fifo_data_o_2__127_, fifo_data_o_2__126_, fifo_data_o_2__125_, fifo_data_o_2__124_, fifo_data_o_2__123_, fifo_data_o_2__122_, fifo_data_o_2__121_, fifo_data_o_2__120_, fifo_data_o_2__119_, fifo_data_o_2__118_, fifo_data_o_2__117_, fifo_data_o_2__116_, fifo_data_o_2__115_, fifo_data_o_2__114_, fifo_data_o_2__113_, fifo_data_o_2__112_, fifo_data_o_2__111_, fifo_data_o_2__110_, fifo_data_o_2__109_, fifo_data_o_2__108_, fifo_data_o_2__107_, fifo_data_o_2__106_, fifo_data_o_2__105_, fifo_data_o_2__104_, fifo_data_o_2__103_, fifo_data_o_2__102_, fifo_data_o_2__101_, fifo_data_o_2__100_, fifo_data_o_2__99_, fifo_data_o_2__98_, fifo_data_o_2__97_, fifo_data_o_2__96_, fifo_data_o_2__95_, fifo_data_o_2__94_, fifo_data_o_2__93_, fifo_data_o_2__92_, fifo_data_o_2__91_, fifo_data_o_2__90_, fifo_data_o_2__89_, fifo_data_o_2__88_, fifo_data_o_2__87_, fifo_data_o_2__86_, fifo_data_o_2__85_, fifo_data_o_2__84_, fifo_data_o_2__83_, fifo_data_o_2__82_, fifo_data_o_2__81_, fifo_data_o_2__80_, fifo_data_o_2__79_, fifo_data_o_2__78_, fifo_data_o_2__77_, fifo_data_o_2__76_, fifo_data_o_2__75_, fifo_data_o_2__74_, fifo_data_o_2__73_, fifo_data_o_2__72_, fifo_data_o_2__71_, fifo_data_o_2__70_, fifo_data_o_2__69_, fifo_data_o_2__68_, fifo_data_o_2__67_, fifo_data_o_2__66_, fifo_data_o_2__65_, fifo_data_o_2__64_, fifo_data_o_2__63_, fifo_data_o_2__62_, fifo_data_o_2__61_, fifo_data_o_2__60_, fifo_data_o_2__59_, fifo_data_o_2__58_, fifo_data_o_2__57_, fifo_data_o_2__56_, fifo_data_o_2__55_, fifo_data_o_2__54_, fifo_data_o_2__53_, fifo_data_o_2__52_, fifo_data_o_2__51_, fifo_data_o_2__50_, fifo_data_o_2__49_, fifo_data_o_2__48_, fifo_data_o_2__47_, fifo_data_o_2__46_, fifo_data_o_2__45_, fifo_data_o_2__44_, fifo_data_o_2__43_, fifo_data_o_2__42_, fifo_data_o_2__41_, fifo_data_o_2__40_, fifo_data_o_2__39_, fifo_data_o_2__38_, fifo_data_o_2__37_, fifo_data_o_2__36_, fifo_data_o_2__35_, fifo_data_o_2__34_, fifo_data_o_2__33_, fifo_data_o_2__32_, fifo_data_o_2__31_, fifo_data_o_2__30_, fifo_data_o_2__29_, fifo_data_o_2__28_, fifo_data_o_2__27_, fifo_data_o_2__26_, fifo_data_o_2__25_, fifo_data_o_2__24_, fifo_data_o_2__23_, fifo_data_o_2__22_, fifo_data_o_2__21_, fifo_data_o_2__20_, fifo_data_o_2__19_, fifo_data_o_2__18_, fifo_data_o_2__17_, fifo_data_o_2__16_, fifo_data_o_2__15_, fifo_data_o_2__14_, fifo_data_o_2__13_, fifo_data_o_2__12_, fifo_data_o_2__11_, fifo_data_o_2__10_, fifo_data_o_2__9_, fifo_data_o_2__8_, fifo_data_o_2__7_, fifo_data_o_2__6_, fifo_data_o_2__5_, fifo_data_o_2__4_, fifo_data_o_2__3_, fifo_data_o_2__2_, fifo_data_o_2__1_, fifo_data_o_2__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_0__4_, arb_sel_o_0__3_, arb_sel_o_0__2_, arb_sel_o_0__1_, arb_sel_o_0__0_ }),
    .data_o(data_o[135:0])
  );

  assign N278 = N0 & local_x_cord_i[0];
  assign N0 = ~1'b0;
  assign N279 = 1'b0 & N1;
  assign N1 = ~local_x_cord_i[0];
  assign N283 = N2 & local_y_cord_i[0];
  assign N2 = ~1'b0;
  assign N284 = 1'b0 & N3;
  assign N3 = ~local_y_cord_i[0];
  assign N4 = fifo_data_o_2__1_ ^ local_y_cord_i[0];
  assign N285 = ~N4;
  assign N5 = fifo_data_o_2__0_ ^ local_x_cord_i[0];
  assign N287 = ~N5;
  assign N288 = N6 & local_x_cord_i[0];
  assign N6 = ~fifo_data_o_2__0_;
  assign N291 = N7 & local_y_cord_i[0];
  assign N7 = ~fifo_data_o_2__1_;
  assign N292 = fifo_data_o_2__1_ & N8;
  assign N8 = ~local_y_cord_i[0];
  assign N9 = fifo_data_o_3__1_ ^ local_y_cord_i[0];
  assign N293 = ~N9;
  assign N10 = fifo_data_o_3__0_ ^ local_x_cord_i[0];
  assign N295 = ~N10;
  assign N296 = N11 & local_x_cord_i[0];
  assign N11 = ~fifo_data_o_3__0_;
  assign N297 = fifo_data_o_3__0_ & N12;
  assign N12 = ~local_x_cord_i[0];
  assign N301 = fifo_data_o_3__1_ & N13;
  assign N13 = ~local_y_cord_i[0];
  assign N323 = out_count_r[2] | out_count_r[3];
  assign N324 = ~N323;
  assign N325 = out_count_r[2] | out_count_r[3];
  assign N326 = ~N325;
  assign N327 = out_count_r[2] | out_count_r[3];
  assign N328 = ~N327;
  assign N329 = out_count_r[2] | out_count_r[3];
  assign N330 = ~N329;
  assign N331 = out_count_r[4] | out_count_r[5];
  assign N332 = ~N331;
  assign N333 = out_count_r[4] | out_count_r[5];
  assign N334 = ~N333;
  assign N335 = out_count_r[4] | out_count_r[5];
  assign N336 = ~N335;
  assign N337 = out_count_r[4] | out_count_r[5];
  assign N338 = ~N337;
  assign N339 = out_count_r[6] | out_count_r[7];
  assign N340 = ~N339;
  assign N341 = out_count_r[6] | out_count_r[7];
  assign N342 = ~N341;
  assign N343 = out_count_r[6] | out_count_r[7];
  assign N344 = ~N343;
  assign N345 = out_count_r[6] | out_count_r[7];
  assign N346 = ~N345;
  assign N347 = out_count_r[8] | out_count_r[9];
  assign N348 = ~N347;
  assign N349 = out_count_r[8] | out_count_r[9];
  assign N350 = ~N349;
  assign N351 = out_count_r[8] | out_count_r[9];
  assign N352 = ~N351;
  assign N353 = out_count_r[8] | out_count_r[9];
  assign N354 = ~N353;
  assign N355 = out_count_r[0] | out_count_r[1];
  assign N356 = ~N355;
  assign N357 = out_count_r[0] | out_count_r[1];
  assign N358 = ~N357;
  assign N359 = out_count_r[0] | out_count_r[1];
  assign N360 = ~N359;
  assign N361 = out_count_r[0] | out_count_r[1];
  assign N362 = ~N361;
  assign N363 = out_count_r[0] | out_count_r[1];
  assign N364 = ~N363;
  assign N365 = out_count_r[0] | out_count_r[1];
  assign N366 = out_count_r[2] | out_count_r[3];
  assign N367 = out_count_r[4] | out_count_r[5];
  assign N368 = out_count_r[6] | out_count_r[7];
  assign N369 = out_count_r[8] | out_count_r[9];
  assign N370 = out_count_r[0] | out_count_r[1];
  assign N371 = out_count_r[4] | out_count_r[5];
  assign N372 = out_count_r[6] | out_count_r[7];
  assign N373 = out_count_r[8] | out_count_r[9];
  assign N374 = out_count_r[0] | out_count_r[1];
  assign N375 = out_count_r[2] | out_count_r[3];
  assign N376 = out_count_r[6] | out_count_r[7];
  assign N377 = out_count_r[8] | out_count_r[9];
  assign N378 = out_count_r[0] | out_count_r[1];
  assign N379 = out_count_r[2] | out_count_r[3];
  assign N380 = out_count_r[4] | out_count_r[5];
  assign N381 = out_count_r[8] | out_count_r[9];
  assign N382 = out_count_r[0] | out_count_r[1];
  assign N383 = out_count_r[2] | out_count_r[3];
  assign N384 = out_count_r[4] | out_count_r[5];
  assign N385 = out_count_r[6] | out_count_r[7];
  assign N386 = count_r[8] | count_r[9];
  assign N387 = ~N386;
  assign N388 = count_r[6] | count_r[7];
  assign N389 = ~N388;
  assign N390 = count_r[4] | count_r[5];
  assign N391 = ~N390;
  assign N392 = count_r[2] | count_r[3];
  assign N393 = ~N392;
  assign N394 = count_r[0] | count_r[1];
  assign N395 = ~N394;
  assign N396 = ~local_y_cord_i[0];
  assign N397 = ~local_x_cord_i[0];
  assign N398 = count_r[0] | count_r[1];
  assign N399 = ~N398;
  assign N400 = count_r[2] | count_r[3];
  assign N401 = ~N400;
  assign N402 = count_r[4] | count_r[5];
  assign N403 = ~N402;
  assign N404 = count_r[6] | count_r[7];
  assign N405 = ~N404;
  assign N406 = count_r[8] | count_r[9];
  assign N407 = ~N406;
  assign N408 = out_count_r[0] | out_count_r[1];
  assign N409 = ~N408;
  assign N410 = out_count_r[2] | out_count_r[3];
  assign N411 = ~N410;
  assign N412 = out_count_r[4] | out_count_r[5];
  assign N413 = ~N412;
  assign N414 = out_count_r[6] | out_count_r[7];
  assign N415 = ~N414;
  assign N416 = out_count_r[8] | out_count_r[9];
  assign N417 = ~N416;
  assign { N126, N125 } = count_r[1:0] - 1'b1;
  assign { N139, N138 } = count_r[3:2] - 1'b1;
  assign { N153, N152 } = count_r[5:4] - 1'b1;
  assign { N167, N166 } = count_r[7:6] - 1'b1;
  assign { N180, N179 } = count_r[9:8] - 1'b1;
  assign { N194, N193 } = out_count_r[1:0] - 1'b1;
  assign { N208, N207 } = out_count_r[3:2] - 1'b1;
  assign { N222, N221 } = out_count_r[5:4] - 1'b1;
  assign { N236, N235 } = out_count_r[7:6] - 1'b1;
  assign { N250, N249 } = out_count_r[9:8] - 1'b1;
  assign { N128, N127 } = (N14)? { 1'b0, 1'b0 } :
                          (N15)? { N126, N125 } : 1'b0;
  assign N14 = N399;
  assign N15 = N398;
  assign { N130, N129 } = (N16)? { N128, N127 } :
                          (N123)? count_r[1:0] : 1'b0;
  assign N16 = fifo_yumi_i[0];
  assign { N132, N131 } = (N17)? { 1'b0, 1'b0 } :
                          (N18)? { N130, N129 } : 1'b0;
  assign N17 = N121;
  assign N18 = N120;
  assign { N141, N140 } = (N19)? { 1'b0, 1'b0 } :
                          (N20)? { N139, N138 } : 1'b0;
  assign N19 = N401;
  assign N20 = N400;
  assign { N143, N142 } = (N21)? { N141, N140 } :
                          (N136)? count_r[3:2] : 1'b0;
  assign N21 = fifo_yumi_i[1];
  assign { N145, N144 } = (N22)? { 1'b0, 1'b0 } :
                          (N23)? { N143, N142 } : 1'b0;
  assign N22 = N134;
  assign N23 = N133;
  assign { N155, N154 } = (N24)? { fifo_data_o_2__3_, fifo_data_o_2__2_ } :
                          (N25)? { N153, N152 } : 1'b0;
  assign N24 = N403;
  assign N25 = N402;
  assign { N157, N156 } = (N26)? { N155, N154 } :
                          (N150)? count_r[5:4] : 1'b0;
  assign N26 = N149;
  assign { N159, N158 } = (N27)? { 1'b0, 1'b0 } :
                          (N28)? { N157, N156 } : 1'b0;
  assign N27 = N147;
  assign N28 = N146;
  assign { N169, N168 } = (N29)? { fifo_data_o_3__3_, fifo_data_o_3__2_ } :
                          (N30)? { N167, N166 } : 1'b0;
  assign N29 = N405;
  assign N30 = N404;
  assign { N171, N170 } = (N31)? { N169, N168 } :
                          (N164)? count_r[7:6] : 1'b0;
  assign N31 = N163;
  assign { N173, N172 } = (N32)? { 1'b0, 1'b0 } :
                          (N33)? { N171, N170 } : 1'b0;
  assign N32 = N161;
  assign N33 = N160;
  assign { N182, N181 } = (N34)? { 1'b0, 1'b0 } :
                          (N35)? { N180, N179 } : 1'b0;
  assign N34 = N407;
  assign N35 = N406;
  assign { N184, N183 } = (N36)? { N182, N181 } :
                          (N177)? count_r[9:8] : 1'b0;
  assign N36 = fifo_yumi_i[4];
  assign { N186, N185 } = (N37)? { 1'b0, 1'b0 } :
                          (N38)? { N184, N183 } : 1'b0;
  assign N37 = N175;
  assign N38 = N174;
  assign { N196, N195 } = (N39)? data_o[3:2] :
                          (N40)? { N194, N193 } : 1'b0;
  assign N39 = N409;
  assign N40 = N408;
  assign { N198, N197 } = (N41)? { N196, N195 } :
                          (N191)? out_count_r[1:0] : 1'b0;
  assign N41 = N190;
  assign { N200, N199 } = (N42)? { 1'b0, 1'b0 } :
                          (N43)? { N198, N197 } : 1'b0;
  assign N42 = N188;
  assign N43 = N187;
  assign { N210, N209 } = (N44)? data_o[139:138] :
                          (N45)? { N208, N207 } : 1'b0;
  assign N44 = N411;
  assign N45 = N410;
  assign { N212, N211 } = (N46)? { N210, N209 } :
                          (N205)? out_count_r[3:2] : 1'b0;
  assign N46 = N204;
  assign { N214, N213 } = (N47)? { 1'b0, 1'b0 } :
                          (N48)? { N212, N211 } : 1'b0;
  assign N47 = N202;
  assign N48 = N201;
  assign { N224, N223 } = (N49)? data_o[275:274] :
                          (N50)? { N222, N221 } : 1'b0;
  assign N49 = N413;
  assign N50 = N412;
  assign { N226, N225 } = (N51)? { N224, N223 } :
                          (N219)? out_count_r[5:4] : 1'b0;
  assign N51 = N218;
  assign { N228, N227 } = (N52)? { 1'b0, 1'b0 } :
                          (N53)? { N226, N225 } : 1'b0;
  assign N52 = N216;
  assign N53 = N215;
  assign { N238, N237 } = (N54)? data_o[411:410] :
                          (N55)? { N236, N235 } : 1'b0;
  assign N54 = N415;
  assign N55 = N414;
  assign { N240, N239 } = (N56)? { N238, N237 } :
                          (N233)? out_count_r[7:6] : 1'b0;
  assign N56 = N232;
  assign { N242, N241 } = (N57)? { 1'b0, 1'b0 } :
                          (N58)? { N240, N239 } : 1'b0;
  assign N57 = N230;
  assign N58 = N229;
  assign { N252, N251 } = (N59)? data_o[547:546] :
                          (N60)? { N250, N249 } : 1'b0;
  assign N59 = N417;
  assign N60 = N416;
  assign { N254, N253 } = (N61)? { N252, N251 } :
                          (N247)? out_count_r[9:8] : 1'b0;
  assign N61 = N246;
  assign { N256, N255 } = (N62)? { 1'b0, 1'b0 } :
                          (N63)? { N254, N253 } : 1'b0;
  assign N62 = N244;
  assign N63 = N243;
  assign arb_valid_0__0_ = (N64)? new_valid_0__0_ :
                           (N65)? N257 : 1'b0;
  assign N64 = N364;
  assign N65 = N363;
  assign arb_valid_0__1_ = (N66)? new_valid_0__1_ :
                           (N67)? N258 : 1'b0;
  assign N66 = N330;
  assign N67 = N329;
  assign arb_valid_0__2_ = (N68)? new_valid_0__2_ :
                           (N69)? N259 : 1'b0;
  assign N68 = N338;
  assign N69 = N337;
  assign arb_valid_0__3_ = (N70)? new_valid_0__3_ :
                           (N71)? N260 : 1'b0;
  assign N70 = N346;
  assign N71 = N345;
  assign arb_valid_0__4_ = (N72)? new_valid_0__4_ :
                           (N73)? N261 : 1'b0;
  assign N72 = N354;
  assign N73 = N353;
  assign arb_valid_1__0_ = (N74)? new_valid_1__0_ :
                           (N75)? N262 : 1'b0;
  assign N74 = N362;
  assign N75 = N361;
  assign arb_valid_1__2_ = (N76)? new_valid_1__2_ :
                           (N77)? N263 : 1'b0;
  assign N76 = N336;
  assign N77 = N335;
  assign arb_valid_1__3_ = (N78)? new_valid_1__3_ :
                           (N79)? N264 : 1'b0;
  assign N78 = N344;
  assign N79 = N343;
  assign arb_valid_1__4_ = (N80)? new_valid_1__4_ :
                           (N81)? N265 : 1'b0;
  assign N80 = N352;
  assign N81 = N351;
  assign arb_valid_2__0_ = (N82)? new_valid_2__0_ :
                           (N83)? N266 : 1'b0;
  assign N82 = N360;
  assign N83 = N359;
  assign arb_valid_2__1_ = (N84)? new_valid_2__1_ :
                           (N85)? N267 : 1'b0;
  assign N84 = N328;
  assign N85 = N327;
  assign arb_valid_2__3_ = (N86)? new_valid_2__3_ :
                           (N87)? N268 : 1'b0;
  assign N86 = N342;
  assign N87 = N341;
  assign arb_valid_2__4_ = (N88)? new_valid_2__4_ :
                           (N89)? N269 : 1'b0;
  assign N88 = N350;
  assign N89 = N349;
  assign arb_valid_3__0_ = (N90)? new_valid_3__0_ :
                           (N91)? N270 : 1'b0;
  assign N90 = N358;
  assign N91 = N357;
  assign arb_valid_3__1_ = (N92)? new_valid_3__1_ :
                           (N93)? N271 : 1'b0;
  assign N92 = N326;
  assign N93 = N325;
  assign arb_valid_3__2_ = (N94)? new_valid_3__2_ :
                           (N95)? N272 : 1'b0;
  assign N94 = N334;
  assign N95 = N333;
  assign arb_valid_3__4_ = (N96)? new_valid_3__4_ :
                           (N97)? N273 : 1'b0;
  assign N96 = N348;
  assign N97 = N347;
  assign arb_valid_4__0_ = (N98)? new_valid_4__0_ :
                           (N99)? N274 : 1'b0;
  assign N98 = N356;
  assign N99 = N355;
  assign arb_valid_4__1_ = (N100)? new_valid_4__1_ :
                           (N101)? N275 : 1'b0;
  assign N100 = N324;
  assign N101 = N323;
  assign arb_valid_4__2_ = (N102)? new_valid_4__2_ :
                           (N103)? N276 : 1'b0;
  assign N102 = N332;
  assign N103 = N331;
  assign arb_valid_4__3_ = (N104)? new_valid_4__3_ :
                           (N105)? N277 : 1'b0;
  assign N104 = N340;
  assign N105 = N339;
  assign { N282, N281, N280 } = (N106)? { N279, N278, N397 } :
                                (N107)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N106 = N396;
  assign N107 = local_y_cord_i[0];
  assign { dest_n_0__4_, dest_n_0__3_, dest_n_0__2_, dest_n_0__1_, dest_n_0__0_ } = (N108)? { N284, N283, N282, N281, N280 } :
                                                                                    (N109)? { dest_r_0__4_, dest_r_0__3_, dest_r_0__2_, dest_r_0__1_, dest_r_0__0_ } : 1'b0;
  assign N108 = N395;
  assign N109 = N394;
  assign { dest_n_1__4_, dest_n_1__3_, dest_n_1__2_, dest_n_1__0_ } = (N110)? { N284, N283, N282, N280 } :
                                                                      (N111)? { dest_r_1__4_, dest_r_1__3_, dest_r_1__2_, dest_r_1__0_ } : 1'b0;
  assign N110 = N393;
  assign N111 = N392;
  assign { N290, N289 } = (N112)? { N288, N287 } :
                          (N286)? { 1'b0, 1'b0 } : 1'b0;
  assign N112 = N285;
  assign { dest_n_2__4_, dest_n_2__3_, dest_n_2__1_, dest_n_2__0_ } = (N113)? { N292, N291, N290, N289 } :
                                                                      (N114)? { dest_r_2__4_, dest_r_2__3_, dest_r_2__1_, dest_r_2__0_ } : 1'b0;
  assign N113 = N391;
  assign N114 = N390;
  assign { N300, N299, N298 } = (N115)? { N297, N296, N295 } :
                                (N294)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N115 = N293;
  assign { dest_n_3__4_, dest_n_3__2_, dest_n_3__1_, dest_n_3__0_ } = (N116)? { N301, N300, N299, N298 } :
                                                                      (N117)? { dest_r_3__4_, dest_r_3__2_, dest_r_3__1_, dest_r_3__0_ } : 1'b0;
  assign N116 = N389;
  assign N117 = N388;
  assign { dest_n_4__3_, dest_n_4__2_, dest_n_4__1_, dest_n_4__0_ } = (N118)? { N283, N282, N281, N280 } :
                                                                      (N119)? { dest_r_4__3_, dest_r_4__2_, dest_r_4__1_, dest_r_4__0_ } : 1'b0;
  assign N118 = N387;
  assign N119 = N386;
  assign N120 = ~reset_i;
  assign N121 = reset_i;
  assign N122 = N120;
  assign N123 = ~fifo_yumi_i[0];
  assign N124 = N122 & fifo_yumi_i[0];
  assign N133 = ~reset_i;
  assign N134 = reset_i;
  assign N135 = N133;
  assign N136 = ~fifo_yumi_i[1];
  assign N137 = N135 & fifo_yumi_i[1];
  assign N146 = ~reset_i;
  assign N147 = reset_i;
  assign N148 = N146;
  assign N149 = fifo_yumi_i[2];
  assign N150 = ~N149;
  assign N151 = N148 & N149;
  assign N160 = ~reset_i;
  assign N161 = reset_i;
  assign N162 = N160;
  assign N163 = fifo_yumi_i[3];
  assign N164 = ~N163;
  assign N165 = N162 & N163;
  assign N174 = ~reset_i;
  assign N175 = reset_i;
  assign N176 = N174;
  assign N177 = ~fifo_yumi_i[4];
  assign N178 = N176 & fifo_yumi_i[4];
  assign new_valid_0__0_ = 1'b0 & dest_n_0__0_;
  assign new_valid_0__1_ = 1'b0 & dest_n_0__1_;
  assign new_valid_0__2_ = 1'b0 & dest_n_0__2_;
  assign new_valid_0__3_ = 1'b0 & dest_n_0__3_;
  assign new_valid_0__4_ = 1'b0 & dest_n_0__4_;
  assign new_valid_1__0_ = 1'b0 & dest_n_1__0_;
  assign new_valid_1__2_ = 1'b0 & dest_n_1__2_;
  assign new_valid_1__3_ = 1'b0 & dest_n_1__3_;
  assign new_valid_1__4_ = 1'b0 & dest_n_1__4_;
  assign new_valid_2__0_ = fifo_valid_o[2] & dest_n_2__0_;
  assign new_valid_2__1_ = fifo_valid_o[2] & dest_n_2__1_;
  assign new_valid_2__3_ = fifo_valid_o[2] & dest_n_2__3_;
  assign new_valid_2__4_ = fifo_valid_o[2] & dest_n_2__4_;
  assign new_valid_3__0_ = fifo_valid_o[3] & dest_n_3__0_;
  assign new_valid_3__1_ = fifo_valid_o[3] & dest_n_3__1_;
  assign new_valid_3__2_ = fifo_valid_o[3] & dest_n_3__2_;
  assign new_valid_3__4_ = fifo_valid_o[3] & dest_n_3__4_;
  assign new_valid_4__0_ = 1'b0 & dest_n_4__0_;
  assign new_valid_4__1_ = 1'b0 & dest_n_4__1_;
  assign new_valid_4__2_ = 1'b0 & dest_n_4__2_;
  assign new_valid_4__3_ = 1'b0 & dest_n_4__3_;
  assign fifo_yumi_i[0] = N420 | arb_grants_o_0__0_;
  assign N420 = N419 | arb_grants_o_0__1_;
  assign N419 = N418 | arb_grants_o_0__2_;
  assign N418 = arb_grants_o_0__4_ | arb_grants_o_0__3_;
  assign fifo_yumi_i[1] = N423 | arb_grants_o_1__0_;
  assign N423 = N422 | 1'b0;
  assign N422 = N421 | arb_grants_o_1__2_;
  assign N421 = arb_grants_o_1__4_ | arb_grants_o_1__3_;
  assign fifo_yumi_i[2] = N426 | arb_grants_o_2__0_;
  assign N426 = N425 | arb_grants_o_2__1_;
  assign N425 = N424 | 1'b0;
  assign N424 = arb_grants_o_2__4_ | arb_grants_o_2__3_;
  assign fifo_yumi_i[3] = N429 | arb_grants_o_3__0_;
  assign N429 = N428 | arb_grants_o_3__1_;
  assign N428 = N427 | arb_grants_o_3__2_;
  assign N427 = arb_grants_o_3__4_ | 1'b0;
  assign fifo_yumi_i[4] = N432 | arb_grants_o_4__0_;
  assign N432 = N431 | arb_grants_o_4__1_;
  assign N431 = N430 | arb_grants_o_4__2_;
  assign N430 = 1'b0 | arb_grants_o_4__3_;
  assign N187 = ~reset_i;
  assign N188 = reset_i;
  assign N189 = N187;
  assign N190 = valid_o[0] & ready_i[0];
  assign N191 = ~N190;
  assign N192 = N189 & N190;
  assign N201 = ~reset_i;
  assign N202 = reset_i;
  assign N203 = N201;
  assign N204 = valid_o[1] & 1'b1;
  assign N205 = ~N204;
  assign N206 = N203 & N204;
  assign N215 = ~reset_i;
  assign N216 = reset_i;
  assign N217 = N215;
  assign N218 = valid_o[2] & ready_i[2];
  assign N219 = ~N218;
  assign N220 = N217 & N218;
  assign N229 = ~reset_i;
  assign N230 = reset_i;
  assign N231 = N229;
  assign N232 = valid_o[3] & 1'b1;
  assign N233 = ~N232;
  assign N234 = N231 & N232;
  assign N243 = ~reset_i;
  assign N244 = reset_i;
  assign N245 = N243;
  assign N246 = valid_o[4] & 1'b1;
  assign N247 = ~N246;
  assign N248 = N245 & N246;
  assign N257 = new_valid_0__0_ & arb_grants_r_0__0_;
  assign N258 = new_valid_0__1_ & arb_grants_r_0__1_;
  assign N259 = new_valid_0__2_ & arb_grants_r_0__2_;
  assign N260 = new_valid_0__3_ & arb_grants_r_0__3_;
  assign N261 = new_valid_0__4_ & arb_grants_r_0__4_;
  assign N262 = new_valid_1__0_ & arb_grants_r_1__0_;
  assign N263 = new_valid_1__2_ & arb_grants_r_1__2_;
  assign N264 = new_valid_1__3_ & arb_grants_r_1__3_;
  assign N265 = new_valid_1__4_ & arb_grants_r_1__4_;
  assign N266 = new_valid_2__0_ & arb_grants_r_2__0_;
  assign N267 = new_valid_2__1_ & arb_grants_r_2__1_;
  assign N268 = new_valid_2__3_ & arb_grants_r_2__3_;
  assign N269 = new_valid_2__4_ & arb_grants_r_2__4_;
  assign N270 = new_valid_3__0_ & arb_grants_r_3__0_;
  assign N271 = new_valid_3__1_ & arb_grants_r_3__1_;
  assign N272 = new_valid_3__2_ & arb_grants_r_3__2_;
  assign N273 = new_valid_3__4_ & arb_grants_r_3__4_;
  assign N274 = new_valid_4__0_ & arb_grants_r_4__0_;
  assign N275 = new_valid_4__1_ & arb_grants_r_4__1_;
  assign N276 = new_valid_4__2_ & arb_grants_r_4__2_;
  assign N277 = new_valid_4__3_ & arb_grants_r_4__3_;
  assign n_3_net_ = valid_o[1] & 1'b1;
  assign n_9_net_ = valid_o[2] & ready_i[2];
  assign n_15_net_ = valid_o[3] & 1'b1;
  assign n_21_net_ = valid_o[4] & 1'b1;
  assign n_27_net_ = valid_o[0] & ready_i[0];
  assign N286 = ~N285;
  assign N294 = ~N293;
  assign N302 = ~N365;
  assign N303 = ~N366;
  assign N304 = ~N367;
  assign N305 = ~N368;
  assign N306 = ~N369;
  assign N307 = ~N370;
  assign N308 = ~N371;
  assign N309 = ~N372;
  assign N310 = ~N373;
  assign N311 = ~N374;
  assign N312 = ~N375;
  assign N313 = ~N376;
  assign N314 = ~N377;
  assign N315 = ~N378;
  assign N316 = ~N379;
  assign N317 = ~N380;
  assign N318 = ~N381;
  assign N319 = ~N382;
  assign N320 = ~N383;
  assign N321 = ~N384;
  assign N322 = ~N385;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { count_r[9:0] } <= { N186, N185, N173, N172, N159, N158, N145, N144, N132, N131 };
      dest_r_0__4_ <= dest_n_0__4_;
      dest_r_0__3_ <= dest_n_0__3_;
      dest_r_0__2_ <= dest_n_0__2_;
      dest_r_0__1_ <= dest_n_0__1_;
      dest_r_0__0_ <= dest_n_0__0_;
      dest_r_1__4_ <= dest_n_1__4_;
      dest_r_1__3_ <= dest_n_1__3_;
      dest_r_1__2_ <= dest_n_1__2_;
      dest_r_1__0_ <= dest_n_1__0_;
      dest_r_2__4_ <= dest_n_2__4_;
      dest_r_2__3_ <= dest_n_2__3_;
      dest_r_2__1_ <= dest_n_2__1_;
      dest_r_2__0_ <= dest_n_2__0_;
      dest_r_3__4_ <= dest_n_3__4_;
      dest_r_3__2_ <= dest_n_3__2_;
      dest_r_3__1_ <= dest_n_3__1_;
      dest_r_3__0_ <= dest_n_3__0_;
      dest_r_4__3_ <= dest_n_4__3_;
      dest_r_4__2_ <= dest_n_4__2_;
      dest_r_4__1_ <= dest_n_4__1_;
      dest_r_4__0_ <= dest_n_4__0_;
      { out_count_r[9:0] } <= { N256, N255, N242, N241, N228, N227, N214, N213, N200, N199 };
    end
    if(N302) begin
      arb_grants_r_0__0_ <= arb_grants_o_0__0_;
    end
    if(N303) begin
      arb_grants_r_0__1_ <= arb_grants_o_0__1_;
    end
    if(N304) begin
      arb_grants_r_0__2_ <= arb_grants_o_0__2_;
    end
    if(N305) begin
      arb_grants_r_0__3_ <= arb_grants_o_0__3_;
    end
    if(N306) begin
      arb_grants_r_0__4_ <= arb_grants_o_0__4_;
    end
    if(N307) begin
      arb_grants_r_1__0_ <= arb_grants_o_1__0_;
    end
    if(N308) begin
      arb_grants_r_1__2_ <= arb_grants_o_1__2_;
    end
    if(N309) begin
      arb_grants_r_1__3_ <= arb_grants_o_1__3_;
    end
    if(N310) begin
      arb_grants_r_1__4_ <= arb_grants_o_1__4_;
    end
    if(N311) begin
      arb_grants_r_2__0_ <= arb_grants_o_2__0_;
    end
    if(N312) begin
      arb_grants_r_2__1_ <= arb_grants_o_2__1_;
    end
    if(N313) begin
      arb_grants_r_2__3_ <= arb_grants_o_2__3_;
    end
    if(N314) begin
      arb_grants_r_2__4_ <= arb_grants_o_2__4_;
    end
    if(N315) begin
      arb_grants_r_3__0_ <= arb_grants_o_3__0_;
    end
    if(N316) begin
      arb_grants_r_3__1_ <= arb_grants_o_3__1_;
    end
    if(N317) begin
      arb_grants_r_3__2_ <= arb_grants_o_3__2_;
    end
    if(N318) begin
      arb_grants_r_3__4_ <= arb_grants_o_3__4_;
    end
    if(N319) begin
      arb_grants_r_4__0_ <= arb_grants_o_4__0_;
    end
    if(N320) begin
      arb_grants_r_4__1_ <= arb_grants_o_4__1_;
    end
    if(N321) begin
      arb_grants_r_4__2_ <= arb_grants_o_4__2_;
    end
    if(N322) begin
      arb_grants_r_4__3_ <= arb_grants_o_4__3_;
    end
  end


endmodule



module bsg_wormhole_router_136_1_1_2_1_1_1_00000015_0000001c
(
  clk_i,
  reset_i,
  local_x_cord_i,
  local_y_cord_i,
  valid_i,
  data_i,
  ready_o,
  valid_o,
  data_o,
  ready_i
);

  input [0:0] local_x_cord_i;
  input [0:0] local_y_cord_i;
  input [4:0] valid_i;
  input [679:0] data_i;
  output [4:0] ready_o;
  output [4:0] valid_o;
  output [679:0] data_o;
  input [4:0] ready_i;
  input clk_i;
  input reset_i;
  wire [4:0] ready_o,valid_o,fifo_yumi_i;
  wire [679:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,fifo_valid_o_1,fifo_data_o_3__135_,fifo_data_o_3__134_,
  fifo_data_o_3__133_,fifo_data_o_3__132_,fifo_data_o_3__131_,fifo_data_o_3__130_,
  fifo_data_o_3__129_,fifo_data_o_3__128_,fifo_data_o_3__127_,fifo_data_o_3__126_,
  fifo_data_o_3__125_,fifo_data_o_3__124_,fifo_data_o_3__123_,fifo_data_o_3__122_,
  fifo_data_o_3__121_,fifo_data_o_3__120_,fifo_data_o_3__119_,fifo_data_o_3__118_,
  fifo_data_o_3__117_,fifo_data_o_3__116_,fifo_data_o_3__115_,fifo_data_o_3__114_,
  fifo_data_o_3__113_,fifo_data_o_3__112_,fifo_data_o_3__111_,fifo_data_o_3__110_,
  fifo_data_o_3__109_,fifo_data_o_3__108_,fifo_data_o_3__107_,fifo_data_o_3__106_,
  fifo_data_o_3__105_,fifo_data_o_3__104_,fifo_data_o_3__103_,fifo_data_o_3__102_,
  fifo_data_o_3__101_,fifo_data_o_3__100_,fifo_data_o_3__99_,fifo_data_o_3__98_,
  fifo_data_o_3__97_,fifo_data_o_3__96_,fifo_data_o_3__95_,fifo_data_o_3__94_,fifo_data_o_3__93_,
  fifo_data_o_3__92_,fifo_data_o_3__91_,fifo_data_o_3__90_,fifo_data_o_3__89_,
  fifo_data_o_3__88_,fifo_data_o_3__87_,fifo_data_o_3__86_,fifo_data_o_3__85_,
  fifo_data_o_3__84_,fifo_data_o_3__83_,fifo_data_o_3__82_,fifo_data_o_3__81_,
  fifo_data_o_3__80_,fifo_data_o_3__79_,fifo_data_o_3__78_,fifo_data_o_3__77_,
  fifo_data_o_3__76_,fifo_data_o_3__75_,fifo_data_o_3__74_,fifo_data_o_3__73_,fifo_data_o_3__72_,
  fifo_data_o_3__71_,fifo_data_o_3__70_,fifo_data_o_3__69_,fifo_data_o_3__68_,
  fifo_data_o_3__67_,fifo_data_o_3__66_,fifo_data_o_3__65_,fifo_data_o_3__64_,
  fifo_data_o_3__63_,fifo_data_o_3__62_,fifo_data_o_3__61_,fifo_data_o_3__60_,
  fifo_data_o_3__59_,fifo_data_o_3__58_,fifo_data_o_3__57_,fifo_data_o_3__56_,fifo_data_o_3__55_,
  fifo_data_o_3__54_,fifo_data_o_3__53_,fifo_data_o_3__52_,fifo_data_o_3__51_,
  fifo_data_o_3__50_,fifo_data_o_3__49_,fifo_data_o_3__48_,fifo_data_o_3__47_,
  fifo_data_o_3__46_,fifo_data_o_3__45_,fifo_data_o_3__44_,fifo_data_o_3__43_,
  fifo_data_o_3__42_,fifo_data_o_3__41_,fifo_data_o_3__40_,fifo_data_o_3__39_,
  fifo_data_o_3__38_,fifo_data_o_3__37_,fifo_data_o_3__36_,fifo_data_o_3__35_,fifo_data_o_3__34_,
  fifo_data_o_3__33_,fifo_data_o_3__32_,fifo_data_o_3__31_,fifo_data_o_3__30_,
  fifo_data_o_3__29_,fifo_data_o_3__28_,fifo_data_o_3__27_,fifo_data_o_3__26_,
  fifo_data_o_3__25_,fifo_data_o_3__24_,fifo_data_o_3__23_,fifo_data_o_3__22_,
  fifo_data_o_3__21_,fifo_data_o_3__20_,fifo_data_o_3__19_,fifo_data_o_3__18_,
  fifo_data_o_3__17_,fifo_data_o_3__16_,fifo_data_o_3__15_,fifo_data_o_3__14_,fifo_data_o_3__13_,
  fifo_data_o_3__12_,fifo_data_o_3__11_,fifo_data_o_3__10_,fifo_data_o_3__9_,
  fifo_data_o_3__8_,fifo_data_o_3__7_,fifo_data_o_3__6_,fifo_data_o_3__5_,
  fifo_data_o_3__4_,fifo_data_o_3__3_,fifo_data_o_3__2_,fifo_data_o_3__1_,fifo_data_o_3__0_,
  fifo_data_o_1__135_,fifo_data_o_1__134_,fifo_data_o_1__133_,fifo_data_o_1__132_,
  fifo_data_o_1__131_,fifo_data_o_1__130_,fifo_data_o_1__129_,fifo_data_o_1__128_,
  fifo_data_o_1__127_,fifo_data_o_1__126_,fifo_data_o_1__125_,fifo_data_o_1__124_,
  fifo_data_o_1__123_,fifo_data_o_1__122_,fifo_data_o_1__121_,fifo_data_o_1__120_,
  fifo_data_o_1__119_,fifo_data_o_1__118_,fifo_data_o_1__117_,fifo_data_o_1__116_,
  fifo_data_o_1__115_,fifo_data_o_1__114_,fifo_data_o_1__113_,fifo_data_o_1__112_,
  fifo_data_o_1__111_,fifo_data_o_1__110_,fifo_data_o_1__109_,fifo_data_o_1__108_,
  fifo_data_o_1__107_,fifo_data_o_1__106_,fifo_data_o_1__105_,fifo_data_o_1__104_,
  fifo_data_o_1__103_,fifo_data_o_1__102_,fifo_data_o_1__101_,fifo_data_o_1__100_,
  fifo_data_o_1__99_,fifo_data_o_1__98_,fifo_data_o_1__97_,fifo_data_o_1__96_,
  fifo_data_o_1__95_,fifo_data_o_1__94_,fifo_data_o_1__93_,fifo_data_o_1__92_,
  fifo_data_o_1__91_,fifo_data_o_1__90_,fifo_data_o_1__89_,fifo_data_o_1__88_,
  fifo_data_o_1__87_,fifo_data_o_1__86_,fifo_data_o_1__85_,fifo_data_o_1__84_,fifo_data_o_1__83_,
  fifo_data_o_1__82_,fifo_data_o_1__81_,fifo_data_o_1__80_,fifo_data_o_1__79_,
  fifo_data_o_1__78_,fifo_data_o_1__77_,fifo_data_o_1__76_,fifo_data_o_1__75_,
  fifo_data_o_1__74_,fifo_data_o_1__73_,fifo_data_o_1__72_,fifo_data_o_1__71_,
  fifo_data_o_1__70_,fifo_data_o_1__69_,fifo_data_o_1__68_,fifo_data_o_1__67_,
  fifo_data_o_1__66_,fifo_data_o_1__65_,fifo_data_o_1__64_,fifo_data_o_1__63_,fifo_data_o_1__62_,
  fifo_data_o_1__61_,fifo_data_o_1__60_,fifo_data_o_1__59_,fifo_data_o_1__58_,
  fifo_data_o_1__57_,fifo_data_o_1__56_,fifo_data_o_1__55_,fifo_data_o_1__54_,
  fifo_data_o_1__53_,fifo_data_o_1__52_,fifo_data_o_1__51_,fifo_data_o_1__50_,
  fifo_data_o_1__49_,fifo_data_o_1__48_,fifo_data_o_1__47_,fifo_data_o_1__46_,fifo_data_o_1__45_,
  fifo_data_o_1__44_,fifo_data_o_1__43_,fifo_data_o_1__42_,fifo_data_o_1__41_,
  fifo_data_o_1__40_,fifo_data_o_1__39_,fifo_data_o_1__38_,fifo_data_o_1__37_,
  fifo_data_o_1__36_,fifo_data_o_1__35_,fifo_data_o_1__34_,fifo_data_o_1__33_,
  fifo_data_o_1__32_,fifo_data_o_1__31_,fifo_data_o_1__30_,fifo_data_o_1__29_,
  fifo_data_o_1__28_,fifo_data_o_1__27_,fifo_data_o_1__26_,fifo_data_o_1__25_,fifo_data_o_1__24_,
  fifo_data_o_1__23_,fifo_data_o_1__22_,fifo_data_o_1__21_,fifo_data_o_1__20_,
  fifo_data_o_1__19_,fifo_data_o_1__18_,fifo_data_o_1__17_,fifo_data_o_1__16_,
  fifo_data_o_1__15_,fifo_data_o_1__14_,fifo_data_o_1__13_,fifo_data_o_1__12_,
  fifo_data_o_1__11_,fifo_data_o_1__10_,fifo_data_o_1__9_,fifo_data_o_1__8_,fifo_data_o_1__7_,
  fifo_data_o_1__6_,fifo_data_o_1__5_,fifo_data_o_1__4_,fifo_data_o_1__3_,
  fifo_data_o_1__2_,fifo_data_o_1__1_,fifo_data_o_1__0_,N120,N121,N122,N123,N124,N125,N126,
  N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,
  N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,
  N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,
  N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,dest_n_4__3_,
  dest_n_4__2_,dest_n_4__1_,dest_n_4__0_,dest_n_3__4_,dest_n_3__2_,dest_n_3__1_,
  dest_n_3__0_,dest_n_2__4_,dest_n_2__3_,dest_n_2__1_,dest_n_2__0_,dest_n_1__4_,
  dest_n_1__3_,dest_n_1__2_,dest_n_1__0_,dest_n_0__4_,dest_n_0__3_,dest_n_0__2_,dest_n_0__1_,
  dest_n_0__0_,new_valid_4__3_,new_valid_4__2_,new_valid_4__1_,new_valid_4__0_,
  new_valid_3__4_,new_valid_3__2_,new_valid_3__1_,new_valid_3__0_,new_valid_2__4_,
  new_valid_2__3_,new_valid_2__1_,new_valid_2__0_,new_valid_1__4_,new_valid_1__3_,
  new_valid_1__2_,new_valid_1__0_,new_valid_0__4_,new_valid_0__3_,new_valid_0__2_,
  new_valid_0__1_,new_valid_0__0_,arb_grants_o_4__3_,arb_grants_o_4__2_,
  arb_grants_o_4__1_,arb_grants_o_4__0_,arb_grants_o_3__4_,arb_grants_o_3__2_,
  arb_grants_o_3__1_,arb_grants_o_3__0_,arb_grants_o_2__4_,arb_grants_o_2__3_,arb_grants_o_2__1_,
  arb_grants_o_2__0_,arb_grants_o_1__4_,arb_grants_o_1__3_,arb_grants_o_1__2_,
  arb_grants_o_1__0_,arb_grants_o_0__4_,arb_grants_o_0__3_,arb_grants_o_0__2_,
  arb_grants_o_0__1_,arb_grants_o_0__0_,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
  N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,
  N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,
  N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,
  N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,arb_valid_4__3_,
  arb_valid_4__2_,arb_valid_4__1_,arb_valid_4__0_,arb_valid_3__4_,arb_valid_3__2_,
  arb_valid_3__1_,arb_valid_3__0_,arb_valid_2__4_,arb_valid_2__3_,arb_valid_2__1_,
  arb_valid_2__0_,arb_valid_1__4_,arb_valid_1__3_,arb_valid_1__2_,arb_valid_1__0_,
  arb_valid_0__4_,arb_valid_0__3_,arb_valid_0__2_,arb_valid_0__1_,arb_valid_0__0_,
  N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,
  N274,N275,N276,N277,n_3_net_,arb_sel_o_4__3_,arb_sel_o_4__2_,arb_sel_o_4__1_,
  arb_sel_o_4__0_,arb_sel_o_3__3_,arb_sel_o_3__2_,arb_sel_o_3__1_,arb_sel_o_3__0_,
  arb_sel_o_2__3_,arb_sel_o_2__2_,arb_sel_o_2__1_,arb_sel_o_2__0_,arb_sel_o_1__3_,
  arb_sel_o_1__2_,arb_sel_o_1__1_,arb_sel_o_1__0_,arb_sel_o_0__4_,arb_sel_o_0__3_,
  arb_sel_o_0__2_,arb_sel_o_0__1_,arb_sel_o_0__0_,n_9_net_,n_15_net_,n_21_net_,
  n_27_net_,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,
  N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,
  N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,
  N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,
  N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,
  N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,
  N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,
  N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,
  N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,
  N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,
  SV2V_UNCONNECTED_1,SV2V_UNCONNECTED_2,SV2V_UNCONNECTED_3,SV2V_UNCONNECTED_4,
  SV2V_UNCONNECTED_5,SV2V_UNCONNECTED_6,SV2V_UNCONNECTED_7,
  SV2V_UNCONNECTED_8,SV2V_UNCONNECTED_9,SV2V_UNCONNECTED_10,SV2V_UNCONNECTED_11;
  wire [3:3] fifo_valid_o;
  reg [9:0] count_r,out_count_r;
  reg dest_r_0__4_,dest_r_0__3_,dest_r_0__2_,dest_r_0__1_,dest_r_0__0_,dest_r_1__4_,
  dest_r_1__3_,dest_r_1__2_,dest_r_1__0_,dest_r_2__4_,dest_r_2__3_,dest_r_2__1_,
  dest_r_2__0_,dest_r_3__4_,dest_r_3__2_,dest_r_3__1_,dest_r_3__0_,dest_r_4__3_,
  dest_r_4__2_,dest_r_4__1_,dest_r_4__0_,arb_grants_r_0__0_,arb_grants_r_0__1_,
  arb_grants_r_0__2_,arb_grants_r_0__3_,arb_grants_r_0__4_,arb_grants_r_1__0_,
  arb_grants_r_1__2_,arb_grants_r_1__3_,arb_grants_r_1__4_,arb_grants_r_2__0_,
  arb_grants_r_2__1_,arb_grants_r_2__3_,arb_grants_r_2__4_,arb_grants_r_3__0_,arb_grants_r_3__1_,
  arb_grants_r_3__2_,arb_grants_r_3__4_,arb_grants_r_4__0_,arb_grants_r_4__1_,
  arb_grants_r_4__2_,arb_grants_r_4__3_;
  assign ready_o[4] = 1'b1;
  assign ready_o[2] = 1'b1;
  assign ready_o[0] = 1'b1;

  bsg_two_fifo_width_p136
  in_ff_1__no_stub_two_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(ready_o[1]),
    .data_i(data_i[271:136]),
    .v_i(valid_i[1]),
    .v_o(fifo_valid_o_1),
    .data_o({ fifo_data_o_1__135_, fifo_data_o_1__134_, fifo_data_o_1__133_, fifo_data_o_1__132_, fifo_data_o_1__131_, fifo_data_o_1__130_, fifo_data_o_1__129_, fifo_data_o_1__128_, fifo_data_o_1__127_, fifo_data_o_1__126_, fifo_data_o_1__125_, fifo_data_o_1__124_, fifo_data_o_1__123_, fifo_data_o_1__122_, fifo_data_o_1__121_, fifo_data_o_1__120_, fifo_data_o_1__119_, fifo_data_o_1__118_, fifo_data_o_1__117_, fifo_data_o_1__116_, fifo_data_o_1__115_, fifo_data_o_1__114_, fifo_data_o_1__113_, fifo_data_o_1__112_, fifo_data_o_1__111_, fifo_data_o_1__110_, fifo_data_o_1__109_, fifo_data_o_1__108_, fifo_data_o_1__107_, fifo_data_o_1__106_, fifo_data_o_1__105_, fifo_data_o_1__104_, fifo_data_o_1__103_, fifo_data_o_1__102_, fifo_data_o_1__101_, fifo_data_o_1__100_, fifo_data_o_1__99_, fifo_data_o_1__98_, fifo_data_o_1__97_, fifo_data_o_1__96_, fifo_data_o_1__95_, fifo_data_o_1__94_, fifo_data_o_1__93_, fifo_data_o_1__92_, fifo_data_o_1__91_, fifo_data_o_1__90_, fifo_data_o_1__89_, fifo_data_o_1__88_, fifo_data_o_1__87_, fifo_data_o_1__86_, fifo_data_o_1__85_, fifo_data_o_1__84_, fifo_data_o_1__83_, fifo_data_o_1__82_, fifo_data_o_1__81_, fifo_data_o_1__80_, fifo_data_o_1__79_, fifo_data_o_1__78_, fifo_data_o_1__77_, fifo_data_o_1__76_, fifo_data_o_1__75_, fifo_data_o_1__74_, fifo_data_o_1__73_, fifo_data_o_1__72_, fifo_data_o_1__71_, fifo_data_o_1__70_, fifo_data_o_1__69_, fifo_data_o_1__68_, fifo_data_o_1__67_, fifo_data_o_1__66_, fifo_data_o_1__65_, fifo_data_o_1__64_, fifo_data_o_1__63_, fifo_data_o_1__62_, fifo_data_o_1__61_, fifo_data_o_1__60_, fifo_data_o_1__59_, fifo_data_o_1__58_, fifo_data_o_1__57_, fifo_data_o_1__56_, fifo_data_o_1__55_, fifo_data_o_1__54_, fifo_data_o_1__53_, fifo_data_o_1__52_, fifo_data_o_1__51_, fifo_data_o_1__50_, fifo_data_o_1__49_, fifo_data_o_1__48_, fifo_data_o_1__47_, fifo_data_o_1__46_, fifo_data_o_1__45_, fifo_data_o_1__44_, fifo_data_o_1__43_, fifo_data_o_1__42_, fifo_data_o_1__41_, fifo_data_o_1__40_, fifo_data_o_1__39_, fifo_data_o_1__38_, fifo_data_o_1__37_, fifo_data_o_1__36_, fifo_data_o_1__35_, fifo_data_o_1__34_, fifo_data_o_1__33_, fifo_data_o_1__32_, fifo_data_o_1__31_, fifo_data_o_1__30_, fifo_data_o_1__29_, fifo_data_o_1__28_, fifo_data_o_1__27_, fifo_data_o_1__26_, fifo_data_o_1__25_, fifo_data_o_1__24_, fifo_data_o_1__23_, fifo_data_o_1__22_, fifo_data_o_1__21_, fifo_data_o_1__20_, fifo_data_o_1__19_, fifo_data_o_1__18_, fifo_data_o_1__17_, fifo_data_o_1__16_, fifo_data_o_1__15_, fifo_data_o_1__14_, fifo_data_o_1__13_, fifo_data_o_1__12_, fifo_data_o_1__11_, fifo_data_o_1__10_, fifo_data_o_1__9_, fifo_data_o_1__8_, fifo_data_o_1__7_, fifo_data_o_1__6_, fifo_data_o_1__5_, fifo_data_o_1__4_, fifo_data_o_1__3_, fifo_data_o_1__2_, fifo_data_o_1__1_, fifo_data_o_1__0_ }),
    .yumi_i(fifo_yumi_i[1])
  );


  bsg_two_fifo_width_p136
  in_ff_3__no_stub_two_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(ready_o[3]),
    .data_i(data_i[543:408]),
    .v_i(valid_i[3]),
    .v_o(fifo_valid_o[3]),
    .data_o({ fifo_data_o_3__135_, fifo_data_o_3__134_, fifo_data_o_3__133_, fifo_data_o_3__132_, fifo_data_o_3__131_, fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_ }),
    .yumi_i(fifo_yumi_i[3])
  );


  bsg_round_robin_arb_inputs_p4
  out_side_1__rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[1]),
    .reqs_i({ arb_valid_4__1_, arb_valid_3__1_, arb_valid_2__1_, arb_valid_0__1_ }),
    .grants_o({ arb_grants_o_4__1_, arb_grants_o_3__1_, arb_grants_o_2__1_, arb_grants_o_0__1_ }),
    .sel_one_hot_o({ arb_sel_o_1__3_, arb_sel_o_1__2_, arb_sel_o_1__1_, arb_sel_o_1__0_ }),
    .v_o(valid_o[1]),
    .tag_o({ SV2V_UNCONNECTED_1, SV2V_UNCONNECTED_2 }),
    .yumi_i(n_3_net_)
  );


  bsg_mux_one_hot_width_p136_els_p4
  out_side_1__mux
  (
    .data_i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_o_3__135_, fifo_data_o_3__134_, fifo_data_o_3__133_, fifo_data_o_3__132_, fifo_data_o_3__131_, fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_1__3_, arb_sel_o_1__2_, arb_sel_o_1__1_, arb_sel_o_1__0_ }),
    .data_o(data_o[271:136])
  );


  bsg_round_robin_arb_inputs_p4
  out_side_2__rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ arb_valid_4__2_, arb_valid_3__2_, arb_valid_1__2_, arb_valid_0__2_ }),
    .grants_o({ arb_grants_o_4__2_, arb_grants_o_3__2_, arb_grants_o_1__2_, arb_grants_o_0__2_ }),
    .sel_one_hot_o({ arb_sel_o_2__3_, arb_sel_o_2__2_, arb_sel_o_2__1_, arb_sel_o_2__0_ }),
    .v_o(valid_o[2]),
    .tag_o({ SV2V_UNCONNECTED_3, SV2V_UNCONNECTED_4 }),
    .yumi_i(n_9_net_)
  );


  bsg_mux_one_hot_width_p136_els_p4
  out_side_2__mux
  (
    .data_i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_o_3__135_, fifo_data_o_3__134_, fifo_data_o_3__133_, fifo_data_o_3__132_, fifo_data_o_3__131_, fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_, fifo_data_o_1__135_, fifo_data_o_1__134_, fifo_data_o_1__133_, fifo_data_o_1__132_, fifo_data_o_1__131_, fifo_data_o_1__130_, fifo_data_o_1__129_, fifo_data_o_1__128_, fifo_data_o_1__127_, fifo_data_o_1__126_, fifo_data_o_1__125_, fifo_data_o_1__124_, fifo_data_o_1__123_, fifo_data_o_1__122_, fifo_data_o_1__121_, fifo_data_o_1__120_, fifo_data_o_1__119_, fifo_data_o_1__118_, fifo_data_o_1__117_, fifo_data_o_1__116_, fifo_data_o_1__115_, fifo_data_o_1__114_, fifo_data_o_1__113_, fifo_data_o_1__112_, fifo_data_o_1__111_, fifo_data_o_1__110_, fifo_data_o_1__109_, fifo_data_o_1__108_, fifo_data_o_1__107_, fifo_data_o_1__106_, fifo_data_o_1__105_, fifo_data_o_1__104_, fifo_data_o_1__103_, fifo_data_o_1__102_, fifo_data_o_1__101_, fifo_data_o_1__100_, fifo_data_o_1__99_, fifo_data_o_1__98_, fifo_data_o_1__97_, fifo_data_o_1__96_, fifo_data_o_1__95_, fifo_data_o_1__94_, fifo_data_o_1__93_, fifo_data_o_1__92_, fifo_data_o_1__91_, fifo_data_o_1__90_, fifo_data_o_1__89_, fifo_data_o_1__88_, fifo_data_o_1__87_, fifo_data_o_1__86_, fifo_data_o_1__85_, fifo_data_o_1__84_, fifo_data_o_1__83_, fifo_data_o_1__82_, fifo_data_o_1__81_, fifo_data_o_1__80_, fifo_data_o_1__79_, fifo_data_o_1__78_, fifo_data_o_1__77_, fifo_data_o_1__76_, fifo_data_o_1__75_, fifo_data_o_1__74_, fifo_data_o_1__73_, fifo_data_o_1__72_, fifo_data_o_1__71_, fifo_data_o_1__70_, fifo_data_o_1__69_, fifo_data_o_1__68_, fifo_data_o_1__67_, fifo_data_o_1__66_, fifo_data_o_1__65_, fifo_data_o_1__64_, fifo_data_o_1__63_, fifo_data_o_1__62_, fifo_data_o_1__61_, fifo_data_o_1__60_, fifo_data_o_1__59_, fifo_data_o_1__58_, fifo_data_o_1__57_, fifo_data_o_1__56_, fifo_data_o_1__55_, fifo_data_o_1__54_, fifo_data_o_1__53_, fifo_data_o_1__52_, fifo_data_o_1__51_, fifo_data_o_1__50_, fifo_data_o_1__49_, fifo_data_o_1__48_, fifo_data_o_1__47_, fifo_data_o_1__46_, fifo_data_o_1__45_, fifo_data_o_1__44_, fifo_data_o_1__43_, fifo_data_o_1__42_, fifo_data_o_1__41_, fifo_data_o_1__40_, fifo_data_o_1__39_, fifo_data_o_1__38_, fifo_data_o_1__37_, fifo_data_o_1__36_, fifo_data_o_1__35_, fifo_data_o_1__34_, fifo_data_o_1__33_, fifo_data_o_1__32_, fifo_data_o_1__31_, fifo_data_o_1__30_, fifo_data_o_1__29_, fifo_data_o_1__28_, fifo_data_o_1__27_, fifo_data_o_1__26_, fifo_data_o_1__25_, fifo_data_o_1__24_, fifo_data_o_1__23_, fifo_data_o_1__22_, fifo_data_o_1__21_, fifo_data_o_1__20_, fifo_data_o_1__19_, fifo_data_o_1__18_, fifo_data_o_1__17_, fifo_data_o_1__16_, fifo_data_o_1__15_, fifo_data_o_1__14_, fifo_data_o_1__13_, fifo_data_o_1__12_, fifo_data_o_1__11_, fifo_data_o_1__10_, fifo_data_o_1__9_, fifo_data_o_1__8_, fifo_data_o_1__7_, fifo_data_o_1__6_, fifo_data_o_1__5_, fifo_data_o_1__4_, fifo_data_o_1__3_, fifo_data_o_1__2_, fifo_data_o_1__1_, fifo_data_o_1__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_2__3_, arb_sel_o_2__2_, arb_sel_o_2__1_, arb_sel_o_2__0_ }),
    .data_o(data_o[407:272])
  );


  bsg_round_robin_arb_inputs_p4
  out_side_3__rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ arb_valid_4__3_, arb_valid_2__3_, arb_valid_1__3_, arb_valid_0__3_ }),
    .grants_o({ arb_grants_o_4__3_, arb_grants_o_2__3_, arb_grants_o_1__3_, arb_grants_o_0__3_ }),
    .sel_one_hot_o({ arb_sel_o_3__3_, arb_sel_o_3__2_, arb_sel_o_3__1_, arb_sel_o_3__0_ }),
    .v_o(valid_o[3]),
    .tag_o({ SV2V_UNCONNECTED_5, SV2V_UNCONNECTED_6 }),
    .yumi_i(n_15_net_)
  );


  bsg_mux_one_hot_width_p136_els_p4
  out_side_3__mux
  (
    .data_i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_o_1__135_, fifo_data_o_1__134_, fifo_data_o_1__133_, fifo_data_o_1__132_, fifo_data_o_1__131_, fifo_data_o_1__130_, fifo_data_o_1__129_, fifo_data_o_1__128_, fifo_data_o_1__127_, fifo_data_o_1__126_, fifo_data_o_1__125_, fifo_data_o_1__124_, fifo_data_o_1__123_, fifo_data_o_1__122_, fifo_data_o_1__121_, fifo_data_o_1__120_, fifo_data_o_1__119_, fifo_data_o_1__118_, fifo_data_o_1__117_, fifo_data_o_1__116_, fifo_data_o_1__115_, fifo_data_o_1__114_, fifo_data_o_1__113_, fifo_data_o_1__112_, fifo_data_o_1__111_, fifo_data_o_1__110_, fifo_data_o_1__109_, fifo_data_o_1__108_, fifo_data_o_1__107_, fifo_data_o_1__106_, fifo_data_o_1__105_, fifo_data_o_1__104_, fifo_data_o_1__103_, fifo_data_o_1__102_, fifo_data_o_1__101_, fifo_data_o_1__100_, fifo_data_o_1__99_, fifo_data_o_1__98_, fifo_data_o_1__97_, fifo_data_o_1__96_, fifo_data_o_1__95_, fifo_data_o_1__94_, fifo_data_o_1__93_, fifo_data_o_1__92_, fifo_data_o_1__91_, fifo_data_o_1__90_, fifo_data_o_1__89_, fifo_data_o_1__88_, fifo_data_o_1__87_, fifo_data_o_1__86_, fifo_data_o_1__85_, fifo_data_o_1__84_, fifo_data_o_1__83_, fifo_data_o_1__82_, fifo_data_o_1__81_, fifo_data_o_1__80_, fifo_data_o_1__79_, fifo_data_o_1__78_, fifo_data_o_1__77_, fifo_data_o_1__76_, fifo_data_o_1__75_, fifo_data_o_1__74_, fifo_data_o_1__73_, fifo_data_o_1__72_, fifo_data_o_1__71_, fifo_data_o_1__70_, fifo_data_o_1__69_, fifo_data_o_1__68_, fifo_data_o_1__67_, fifo_data_o_1__66_, fifo_data_o_1__65_, fifo_data_o_1__64_, fifo_data_o_1__63_, fifo_data_o_1__62_, fifo_data_o_1__61_, fifo_data_o_1__60_, fifo_data_o_1__59_, fifo_data_o_1__58_, fifo_data_o_1__57_, fifo_data_o_1__56_, fifo_data_o_1__55_, fifo_data_o_1__54_, fifo_data_o_1__53_, fifo_data_o_1__52_, fifo_data_o_1__51_, fifo_data_o_1__50_, fifo_data_o_1__49_, fifo_data_o_1__48_, fifo_data_o_1__47_, fifo_data_o_1__46_, fifo_data_o_1__45_, fifo_data_o_1__44_, fifo_data_o_1__43_, fifo_data_o_1__42_, fifo_data_o_1__41_, fifo_data_o_1__40_, fifo_data_o_1__39_, fifo_data_o_1__38_, fifo_data_o_1__37_, fifo_data_o_1__36_, fifo_data_o_1__35_, fifo_data_o_1__34_, fifo_data_o_1__33_, fifo_data_o_1__32_, fifo_data_o_1__31_, fifo_data_o_1__30_, fifo_data_o_1__29_, fifo_data_o_1__28_, fifo_data_o_1__27_, fifo_data_o_1__26_, fifo_data_o_1__25_, fifo_data_o_1__24_, fifo_data_o_1__23_, fifo_data_o_1__22_, fifo_data_o_1__21_, fifo_data_o_1__20_, fifo_data_o_1__19_, fifo_data_o_1__18_, fifo_data_o_1__17_, fifo_data_o_1__16_, fifo_data_o_1__15_, fifo_data_o_1__14_, fifo_data_o_1__13_, fifo_data_o_1__12_, fifo_data_o_1__11_, fifo_data_o_1__10_, fifo_data_o_1__9_, fifo_data_o_1__8_, fifo_data_o_1__7_, fifo_data_o_1__6_, fifo_data_o_1__5_, fifo_data_o_1__4_, fifo_data_o_1__3_, fifo_data_o_1__2_, fifo_data_o_1__1_, fifo_data_o_1__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_3__3_, arb_sel_o_3__2_, arb_sel_o_3__1_, arb_sel_o_3__0_ }),
    .data_o(data_o[543:408])
  );


  bsg_round_robin_arb_inputs_p4
  out_side_4__rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ arb_valid_3__4_, arb_valid_2__4_, arb_valid_1__4_, arb_valid_0__4_ }),
    .grants_o({ arb_grants_o_3__4_, arb_grants_o_2__4_, arb_grants_o_1__4_, arb_grants_o_0__4_ }),
    .sel_one_hot_o({ arb_sel_o_4__3_, arb_sel_o_4__2_, arb_sel_o_4__1_, arb_sel_o_4__0_ }),
    .v_o(valid_o[4]),
    .tag_o({ SV2V_UNCONNECTED_7, SV2V_UNCONNECTED_8 }),
    .yumi_i(n_21_net_)
  );


  bsg_mux_one_hot_width_p136_els_p4
  out_side_4__mux
  (
    .data_i({ fifo_data_o_3__135_, fifo_data_o_3__134_, fifo_data_o_3__133_, fifo_data_o_3__132_, fifo_data_o_3__131_, fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_o_1__135_, fifo_data_o_1__134_, fifo_data_o_1__133_, fifo_data_o_1__132_, fifo_data_o_1__131_, fifo_data_o_1__130_, fifo_data_o_1__129_, fifo_data_o_1__128_, fifo_data_o_1__127_, fifo_data_o_1__126_, fifo_data_o_1__125_, fifo_data_o_1__124_, fifo_data_o_1__123_, fifo_data_o_1__122_, fifo_data_o_1__121_, fifo_data_o_1__120_, fifo_data_o_1__119_, fifo_data_o_1__118_, fifo_data_o_1__117_, fifo_data_o_1__116_, fifo_data_o_1__115_, fifo_data_o_1__114_, fifo_data_o_1__113_, fifo_data_o_1__112_, fifo_data_o_1__111_, fifo_data_o_1__110_, fifo_data_o_1__109_, fifo_data_o_1__108_, fifo_data_o_1__107_, fifo_data_o_1__106_, fifo_data_o_1__105_, fifo_data_o_1__104_, fifo_data_o_1__103_, fifo_data_o_1__102_, fifo_data_o_1__101_, fifo_data_o_1__100_, fifo_data_o_1__99_, fifo_data_o_1__98_, fifo_data_o_1__97_, fifo_data_o_1__96_, fifo_data_o_1__95_, fifo_data_o_1__94_, fifo_data_o_1__93_, fifo_data_o_1__92_, fifo_data_o_1__91_, fifo_data_o_1__90_, fifo_data_o_1__89_, fifo_data_o_1__88_, fifo_data_o_1__87_, fifo_data_o_1__86_, fifo_data_o_1__85_, fifo_data_o_1__84_, fifo_data_o_1__83_, fifo_data_o_1__82_, fifo_data_o_1__81_, fifo_data_o_1__80_, fifo_data_o_1__79_, fifo_data_o_1__78_, fifo_data_o_1__77_, fifo_data_o_1__76_, fifo_data_o_1__75_, fifo_data_o_1__74_, fifo_data_o_1__73_, fifo_data_o_1__72_, fifo_data_o_1__71_, fifo_data_o_1__70_, fifo_data_o_1__69_, fifo_data_o_1__68_, fifo_data_o_1__67_, fifo_data_o_1__66_, fifo_data_o_1__65_, fifo_data_o_1__64_, fifo_data_o_1__63_, fifo_data_o_1__62_, fifo_data_o_1__61_, fifo_data_o_1__60_, fifo_data_o_1__59_, fifo_data_o_1__58_, fifo_data_o_1__57_, fifo_data_o_1__56_, fifo_data_o_1__55_, fifo_data_o_1__54_, fifo_data_o_1__53_, fifo_data_o_1__52_, fifo_data_o_1__51_, fifo_data_o_1__50_, fifo_data_o_1__49_, fifo_data_o_1__48_, fifo_data_o_1__47_, fifo_data_o_1__46_, fifo_data_o_1__45_, fifo_data_o_1__44_, fifo_data_o_1__43_, fifo_data_o_1__42_, fifo_data_o_1__41_, fifo_data_o_1__40_, fifo_data_o_1__39_, fifo_data_o_1__38_, fifo_data_o_1__37_, fifo_data_o_1__36_, fifo_data_o_1__35_, fifo_data_o_1__34_, fifo_data_o_1__33_, fifo_data_o_1__32_, fifo_data_o_1__31_, fifo_data_o_1__30_, fifo_data_o_1__29_, fifo_data_o_1__28_, fifo_data_o_1__27_, fifo_data_o_1__26_, fifo_data_o_1__25_, fifo_data_o_1__24_, fifo_data_o_1__23_, fifo_data_o_1__22_, fifo_data_o_1__21_, fifo_data_o_1__20_, fifo_data_o_1__19_, fifo_data_o_1__18_, fifo_data_o_1__17_, fifo_data_o_1__16_, fifo_data_o_1__15_, fifo_data_o_1__14_, fifo_data_o_1__13_, fifo_data_o_1__12_, fifo_data_o_1__11_, fifo_data_o_1__10_, fifo_data_o_1__9_, fifo_data_o_1__8_, fifo_data_o_1__7_, fifo_data_o_1__6_, fifo_data_o_1__5_, fifo_data_o_1__4_, fifo_data_o_1__3_, fifo_data_o_1__2_, fifo_data_o_1__1_, fifo_data_o_1__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_4__3_, arb_sel_o_4__2_, arb_sel_o_4__1_, arb_sel_o_4__0_ }),
    .data_o(data_o[679:544])
  );


  bsg_round_robin_arb_inputs_p5
  rr_arb_proc
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[0]),
    .reqs_i({ arb_valid_4__0_, arb_valid_3__0_, arb_valid_2__0_, arb_valid_1__0_, arb_valid_0__0_ }),
    .grants_o({ arb_grants_o_4__0_, arb_grants_o_3__0_, arb_grants_o_2__0_, arb_grants_o_1__0_, arb_grants_o_0__0_ }),
    .sel_one_hot_o({ arb_sel_o_0__4_, arb_sel_o_0__3_, arb_sel_o_0__2_, arb_sel_o_0__1_, arb_sel_o_0__0_ }),
    .v_o(valid_o[0]),
    .tag_o({ SV2V_UNCONNECTED_9, SV2V_UNCONNECTED_10, SV2V_UNCONNECTED_11 }),
    .yumi_i(n_27_net_)
  );


  bsg_mux_one_hot_width_p136_els_p5
  mux_proc
  (
    .data_i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_o_3__135_, fifo_data_o_3__134_, fifo_data_o_3__133_, fifo_data_o_3__132_, fifo_data_o_3__131_, fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_o_1__135_, fifo_data_o_1__134_, fifo_data_o_1__133_, fifo_data_o_1__132_, fifo_data_o_1__131_, fifo_data_o_1__130_, fifo_data_o_1__129_, fifo_data_o_1__128_, fifo_data_o_1__127_, fifo_data_o_1__126_, fifo_data_o_1__125_, fifo_data_o_1__124_, fifo_data_o_1__123_, fifo_data_o_1__122_, fifo_data_o_1__121_, fifo_data_o_1__120_, fifo_data_o_1__119_, fifo_data_o_1__118_, fifo_data_o_1__117_, fifo_data_o_1__116_, fifo_data_o_1__115_, fifo_data_o_1__114_, fifo_data_o_1__113_, fifo_data_o_1__112_, fifo_data_o_1__111_, fifo_data_o_1__110_, fifo_data_o_1__109_, fifo_data_o_1__108_, fifo_data_o_1__107_, fifo_data_o_1__106_, fifo_data_o_1__105_, fifo_data_o_1__104_, fifo_data_o_1__103_, fifo_data_o_1__102_, fifo_data_o_1__101_, fifo_data_o_1__100_, fifo_data_o_1__99_, fifo_data_o_1__98_, fifo_data_o_1__97_, fifo_data_o_1__96_, fifo_data_o_1__95_, fifo_data_o_1__94_, fifo_data_o_1__93_, fifo_data_o_1__92_, fifo_data_o_1__91_, fifo_data_o_1__90_, fifo_data_o_1__89_, fifo_data_o_1__88_, fifo_data_o_1__87_, fifo_data_o_1__86_, fifo_data_o_1__85_, fifo_data_o_1__84_, fifo_data_o_1__83_, fifo_data_o_1__82_, fifo_data_o_1__81_, fifo_data_o_1__80_, fifo_data_o_1__79_, fifo_data_o_1__78_, fifo_data_o_1__77_, fifo_data_o_1__76_, fifo_data_o_1__75_, fifo_data_o_1__74_, fifo_data_o_1__73_, fifo_data_o_1__72_, fifo_data_o_1__71_, fifo_data_o_1__70_, fifo_data_o_1__69_, fifo_data_o_1__68_, fifo_data_o_1__67_, fifo_data_o_1__66_, fifo_data_o_1__65_, fifo_data_o_1__64_, fifo_data_o_1__63_, fifo_data_o_1__62_, fifo_data_o_1__61_, fifo_data_o_1__60_, fifo_data_o_1__59_, fifo_data_o_1__58_, fifo_data_o_1__57_, fifo_data_o_1__56_, fifo_data_o_1__55_, fifo_data_o_1__54_, fifo_data_o_1__53_, fifo_data_o_1__52_, fifo_data_o_1__51_, fifo_data_o_1__50_, fifo_data_o_1__49_, fifo_data_o_1__48_, fifo_data_o_1__47_, fifo_data_o_1__46_, fifo_data_o_1__45_, fifo_data_o_1__44_, fifo_data_o_1__43_, fifo_data_o_1__42_, fifo_data_o_1__41_, fifo_data_o_1__40_, fifo_data_o_1__39_, fifo_data_o_1__38_, fifo_data_o_1__37_, fifo_data_o_1__36_, fifo_data_o_1__35_, fifo_data_o_1__34_, fifo_data_o_1__33_, fifo_data_o_1__32_, fifo_data_o_1__31_, fifo_data_o_1__30_, fifo_data_o_1__29_, fifo_data_o_1__28_, fifo_data_o_1__27_, fifo_data_o_1__26_, fifo_data_o_1__25_, fifo_data_o_1__24_, fifo_data_o_1__23_, fifo_data_o_1__22_, fifo_data_o_1__21_, fifo_data_o_1__20_, fifo_data_o_1__19_, fifo_data_o_1__18_, fifo_data_o_1__17_, fifo_data_o_1__16_, fifo_data_o_1__15_, fifo_data_o_1__14_, fifo_data_o_1__13_, fifo_data_o_1__12_, fifo_data_o_1__11_, fifo_data_o_1__10_, fifo_data_o_1__9_, fifo_data_o_1__8_, fifo_data_o_1__7_, fifo_data_o_1__6_, fifo_data_o_1__5_, fifo_data_o_1__4_, fifo_data_o_1__3_, fifo_data_o_1__2_, fifo_data_o_1__1_, fifo_data_o_1__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_0__4_, arb_sel_o_0__3_, arb_sel_o_0__2_, arb_sel_o_0__1_, arb_sel_o_0__0_ }),
    .data_o(data_o[135:0])
  );

  assign N278 = N0 & local_x_cord_i[0];
  assign N0 = ~1'b0;
  assign N279 = 1'b0 & N1;
  assign N1 = ~local_x_cord_i[0];
  assign N283 = N2 & local_y_cord_i[0];
  assign N2 = ~1'b0;
  assign N284 = 1'b0 & N3;
  assign N3 = ~local_y_cord_i[0];
  assign N4 = fifo_data_o_1__1_ ^ local_y_cord_i[0];
  assign N285 = ~N4;
  assign N5 = fifo_data_o_1__0_ ^ local_x_cord_i[0];
  assign N287 = ~N5;
  assign N288 = fifo_data_o_1__0_ & N6;
  assign N6 = ~local_x_cord_i[0];
  assign N291 = N7 & local_y_cord_i[0];
  assign N7 = ~fifo_data_o_1__1_;
  assign N292 = fifo_data_o_1__1_ & N8;
  assign N8 = ~local_y_cord_i[0];
  assign N9 = fifo_data_o_3__1_ ^ local_y_cord_i[0];
  assign N293 = ~N9;
  assign N10 = fifo_data_o_3__0_ ^ local_x_cord_i[0];
  assign N295 = ~N10;
  assign N296 = N11 & local_x_cord_i[0];
  assign N11 = ~fifo_data_o_3__0_;
  assign N297 = fifo_data_o_3__0_ & N12;
  assign N12 = ~local_x_cord_i[0];
  assign N301 = fifo_data_o_3__1_ & N13;
  assign N13 = ~local_y_cord_i[0];
  assign N323 = out_count_r[2] | out_count_r[3];
  assign N324 = ~N323;
  assign N325 = out_count_r[2] | out_count_r[3];
  assign N326 = ~N325;
  assign N327 = out_count_r[2] | out_count_r[3];
  assign N328 = ~N327;
  assign N329 = out_count_r[2] | out_count_r[3];
  assign N330 = ~N329;
  assign N331 = out_count_r[4] | out_count_r[5];
  assign N332 = ~N331;
  assign N333 = out_count_r[4] | out_count_r[5];
  assign N334 = ~N333;
  assign N335 = out_count_r[4] | out_count_r[5];
  assign N336 = ~N335;
  assign N337 = out_count_r[4] | out_count_r[5];
  assign N338 = ~N337;
  assign N339 = out_count_r[6] | out_count_r[7];
  assign N340 = ~N339;
  assign N341 = out_count_r[6] | out_count_r[7];
  assign N342 = ~N341;
  assign N343 = out_count_r[6] | out_count_r[7];
  assign N344 = ~N343;
  assign N345 = out_count_r[6] | out_count_r[7];
  assign N346 = ~N345;
  assign N347 = out_count_r[8] | out_count_r[9];
  assign N348 = ~N347;
  assign N349 = out_count_r[8] | out_count_r[9];
  assign N350 = ~N349;
  assign N351 = out_count_r[8] | out_count_r[9];
  assign N352 = ~N351;
  assign N353 = out_count_r[8] | out_count_r[9];
  assign N354 = ~N353;
  assign N355 = out_count_r[0] | out_count_r[1];
  assign N356 = ~N355;
  assign N357 = out_count_r[0] | out_count_r[1];
  assign N358 = ~N357;
  assign N359 = out_count_r[0] | out_count_r[1];
  assign N360 = ~N359;
  assign N361 = out_count_r[0] | out_count_r[1];
  assign N362 = ~N361;
  assign N363 = out_count_r[0] | out_count_r[1];
  assign N364 = ~N363;
  assign N365 = out_count_r[0] | out_count_r[1];
  assign N366 = out_count_r[2] | out_count_r[3];
  assign N367 = out_count_r[4] | out_count_r[5];
  assign N368 = out_count_r[6] | out_count_r[7];
  assign N369 = out_count_r[8] | out_count_r[9];
  assign N370 = out_count_r[0] | out_count_r[1];
  assign N371 = out_count_r[4] | out_count_r[5];
  assign N372 = out_count_r[6] | out_count_r[7];
  assign N373 = out_count_r[8] | out_count_r[9];
  assign N374 = out_count_r[0] | out_count_r[1];
  assign N375 = out_count_r[2] | out_count_r[3];
  assign N376 = out_count_r[6] | out_count_r[7];
  assign N377 = out_count_r[8] | out_count_r[9];
  assign N378 = out_count_r[0] | out_count_r[1];
  assign N379 = out_count_r[2] | out_count_r[3];
  assign N380 = out_count_r[4] | out_count_r[5];
  assign N381 = out_count_r[8] | out_count_r[9];
  assign N382 = out_count_r[0] | out_count_r[1];
  assign N383 = out_count_r[2] | out_count_r[3];
  assign N384 = out_count_r[4] | out_count_r[5];
  assign N385 = out_count_r[6] | out_count_r[7];
  assign N386 = count_r[8] | count_r[9];
  assign N387 = ~N386;
  assign N388 = count_r[6] | count_r[7];
  assign N389 = ~N388;
  assign N390 = count_r[4] | count_r[5];
  assign N391 = ~N390;
  assign N392 = count_r[2] | count_r[3];
  assign N393 = ~N392;
  assign N394 = count_r[0] | count_r[1];
  assign N395 = ~N394;
  assign N396 = ~local_y_cord_i[0];
  assign N397 = ~local_x_cord_i[0];
  assign N398 = count_r[0] | count_r[1];
  assign N399 = ~N398;
  assign N400 = count_r[2] | count_r[3];
  assign N401 = ~N400;
  assign N402 = count_r[4] | count_r[5];
  assign N403 = ~N402;
  assign N404 = count_r[6] | count_r[7];
  assign N405 = ~N404;
  assign N406 = count_r[8] | count_r[9];
  assign N407 = ~N406;
  assign N408 = out_count_r[0] | out_count_r[1];
  assign N409 = ~N408;
  assign N410 = out_count_r[2] | out_count_r[3];
  assign N411 = ~N410;
  assign N412 = out_count_r[4] | out_count_r[5];
  assign N413 = ~N412;
  assign N414 = out_count_r[6] | out_count_r[7];
  assign N415 = ~N414;
  assign N416 = out_count_r[8] | out_count_r[9];
  assign N417 = ~N416;
  assign { N126, N125 } = count_r[1:0] - 1'b1;
  assign { N140, N139 } = count_r[3:2] - 1'b1;
  assign { N153, N152 } = count_r[5:4] - 1'b1;
  assign { N167, N166 } = count_r[7:6] - 1'b1;
  assign { N180, N179 } = count_r[9:8] - 1'b1;
  assign { N194, N193 } = out_count_r[1:0] - 1'b1;
  assign { N208, N207 } = out_count_r[3:2] - 1'b1;
  assign { N222, N221 } = out_count_r[5:4] - 1'b1;
  assign { N236, N235 } = out_count_r[7:6] - 1'b1;
  assign { N250, N249 } = out_count_r[9:8] - 1'b1;
  assign { N128, N127 } = (N14)? { 1'b0, 1'b0 } :
                          (N15)? { N126, N125 } : 1'b0;
  assign N14 = N399;
  assign N15 = N398;
  assign { N130, N129 } = (N16)? { N128, N127 } :
                          (N123)? count_r[1:0] : 1'b0;
  assign N16 = fifo_yumi_i[0];
  assign { N132, N131 } = (N17)? { 1'b0, 1'b0 } :
                          (N18)? { N130, N129 } : 1'b0;
  assign N17 = N121;
  assign N18 = N120;
  assign { N142, N141 } = (N19)? { fifo_data_o_1__3_, fifo_data_o_1__2_ } :
                          (N20)? { N140, N139 } : 1'b0;
  assign N19 = N401;
  assign N20 = N400;
  assign { N144, N143 } = (N21)? { N142, N141 } :
                          (N137)? count_r[3:2] : 1'b0;
  assign N21 = N136;
  assign { N146, N145 } = (N22)? { 1'b0, 1'b0 } :
                          (N23)? { N144, N143 } : 1'b0;
  assign N22 = N134;
  assign N23 = N133;
  assign { N155, N154 } = (N24)? { 1'b0, 1'b0 } :
                          (N25)? { N153, N152 } : 1'b0;
  assign N24 = N403;
  assign N25 = N402;
  assign { N157, N156 } = (N26)? { N155, N154 } :
                          (N150)? count_r[5:4] : 1'b0;
  assign N26 = fifo_yumi_i[2];
  assign { N159, N158 } = (N27)? { 1'b0, 1'b0 } :
                          (N28)? { N157, N156 } : 1'b0;
  assign N27 = N148;
  assign N28 = N147;
  assign { N169, N168 } = (N29)? { fifo_data_o_3__3_, fifo_data_o_3__2_ } :
                          (N30)? { N167, N166 } : 1'b0;
  assign N29 = N405;
  assign N30 = N404;
  assign { N171, N170 } = (N31)? { N169, N168 } :
                          (N164)? count_r[7:6] : 1'b0;
  assign N31 = N163;
  assign { N173, N172 } = (N32)? { 1'b0, 1'b0 } :
                          (N33)? { N171, N170 } : 1'b0;
  assign N32 = N161;
  assign N33 = N160;
  assign { N182, N181 } = (N34)? { 1'b0, 1'b0 } :
                          (N35)? { N180, N179 } : 1'b0;
  assign N34 = N407;
  assign N35 = N406;
  assign { N184, N183 } = (N36)? { N182, N181 } :
                          (N177)? count_r[9:8] : 1'b0;
  assign N36 = fifo_yumi_i[4];
  assign { N186, N185 } = (N37)? { 1'b0, 1'b0 } :
                          (N38)? { N184, N183 } : 1'b0;
  assign N37 = N175;
  assign N38 = N174;
  assign { N196, N195 } = (N39)? data_o[3:2] :
                          (N40)? { N194, N193 } : 1'b0;
  assign N39 = N409;
  assign N40 = N408;
  assign { N198, N197 } = (N41)? { N196, N195 } :
                          (N191)? out_count_r[1:0] : 1'b0;
  assign N41 = N190;
  assign { N200, N199 } = (N42)? { 1'b0, 1'b0 } :
                          (N43)? { N198, N197 } : 1'b0;
  assign N42 = N188;
  assign N43 = N187;
  assign { N210, N209 } = (N44)? data_o[139:138] :
                          (N45)? { N208, N207 } : 1'b0;
  assign N44 = N411;
  assign N45 = N410;
  assign { N212, N211 } = (N46)? { N210, N209 } :
                          (N205)? out_count_r[3:2] : 1'b0;
  assign N46 = N204;
  assign { N214, N213 } = (N47)? { 1'b0, 1'b0 } :
                          (N48)? { N212, N211 } : 1'b0;
  assign N47 = N202;
  assign N48 = N201;
  assign { N224, N223 } = (N49)? data_o[275:274] :
                          (N50)? { N222, N221 } : 1'b0;
  assign N49 = N413;
  assign N50 = N412;
  assign { N226, N225 } = (N51)? { N224, N223 } :
                          (N219)? out_count_r[5:4] : 1'b0;
  assign N51 = N218;
  assign { N228, N227 } = (N52)? { 1'b0, 1'b0 } :
                          (N53)? { N226, N225 } : 1'b0;
  assign N52 = N216;
  assign N53 = N215;
  assign { N238, N237 } = (N54)? data_o[411:410] :
                          (N55)? { N236, N235 } : 1'b0;
  assign N54 = N415;
  assign N55 = N414;
  assign { N240, N239 } = (N56)? { N238, N237 } :
                          (N233)? out_count_r[7:6] : 1'b0;
  assign N56 = N232;
  assign { N242, N241 } = (N57)? { 1'b0, 1'b0 } :
                          (N58)? { N240, N239 } : 1'b0;
  assign N57 = N230;
  assign N58 = N229;
  assign { N252, N251 } = (N59)? data_o[547:546] :
                          (N60)? { N250, N249 } : 1'b0;
  assign N59 = N417;
  assign N60 = N416;
  assign { N254, N253 } = (N61)? { N252, N251 } :
                          (N247)? out_count_r[9:8] : 1'b0;
  assign N61 = N246;
  assign { N256, N255 } = (N62)? { 1'b0, 1'b0 } :
                          (N63)? { N254, N253 } : 1'b0;
  assign N62 = N244;
  assign N63 = N243;
  assign arb_valid_0__0_ = (N64)? new_valid_0__0_ :
                           (N65)? N257 : 1'b0;
  assign N64 = N364;
  assign N65 = N363;
  assign arb_valid_0__1_ = (N66)? new_valid_0__1_ :
                           (N67)? N258 : 1'b0;
  assign N66 = N330;
  assign N67 = N329;
  assign arb_valid_0__2_ = (N68)? new_valid_0__2_ :
                           (N69)? N259 : 1'b0;
  assign N68 = N338;
  assign N69 = N337;
  assign arb_valid_0__3_ = (N70)? new_valid_0__3_ :
                           (N71)? N260 : 1'b0;
  assign N70 = N346;
  assign N71 = N345;
  assign arb_valid_0__4_ = (N72)? new_valid_0__4_ :
                           (N73)? N261 : 1'b0;
  assign N72 = N354;
  assign N73 = N353;
  assign arb_valid_1__0_ = (N74)? new_valid_1__0_ :
                           (N75)? N262 : 1'b0;
  assign N74 = N362;
  assign N75 = N361;
  assign arb_valid_1__2_ = (N76)? new_valid_1__2_ :
                           (N77)? N263 : 1'b0;
  assign N76 = N336;
  assign N77 = N335;
  assign arb_valid_1__3_ = (N78)? new_valid_1__3_ :
                           (N79)? N264 : 1'b0;
  assign N78 = N344;
  assign N79 = N343;
  assign arb_valid_1__4_ = (N80)? new_valid_1__4_ :
                           (N81)? N265 : 1'b0;
  assign N80 = N352;
  assign N81 = N351;
  assign arb_valid_2__0_ = (N82)? new_valid_2__0_ :
                           (N83)? N266 : 1'b0;
  assign N82 = N360;
  assign N83 = N359;
  assign arb_valid_2__1_ = (N84)? new_valid_2__1_ :
                           (N85)? N267 : 1'b0;
  assign N84 = N328;
  assign N85 = N327;
  assign arb_valid_2__3_ = (N86)? new_valid_2__3_ :
                           (N87)? N268 : 1'b0;
  assign N86 = N342;
  assign N87 = N341;
  assign arb_valid_2__4_ = (N88)? new_valid_2__4_ :
                           (N89)? N269 : 1'b0;
  assign N88 = N350;
  assign N89 = N349;
  assign arb_valid_3__0_ = (N90)? new_valid_3__0_ :
                           (N91)? N270 : 1'b0;
  assign N90 = N358;
  assign N91 = N357;
  assign arb_valid_3__1_ = (N92)? new_valid_3__1_ :
                           (N93)? N271 : 1'b0;
  assign N92 = N326;
  assign N93 = N325;
  assign arb_valid_3__2_ = (N94)? new_valid_3__2_ :
                           (N95)? N272 : 1'b0;
  assign N94 = N334;
  assign N95 = N333;
  assign arb_valid_3__4_ = (N96)? new_valid_3__4_ :
                           (N97)? N273 : 1'b0;
  assign N96 = N348;
  assign N97 = N347;
  assign arb_valid_4__0_ = (N98)? new_valid_4__0_ :
                           (N99)? N274 : 1'b0;
  assign N98 = N356;
  assign N99 = N355;
  assign arb_valid_4__1_ = (N100)? new_valid_4__1_ :
                           (N101)? N275 : 1'b0;
  assign N100 = N324;
  assign N101 = N323;
  assign arb_valid_4__2_ = (N102)? new_valid_4__2_ :
                           (N103)? N276 : 1'b0;
  assign N102 = N332;
  assign N103 = N331;
  assign arb_valid_4__3_ = (N104)? new_valid_4__3_ :
                           (N105)? N277 : 1'b0;
  assign N104 = N340;
  assign N105 = N339;
  assign { N282, N281, N280 } = (N106)? { N279, N278, N397 } :
                                (N107)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N106 = N396;
  assign N107 = local_y_cord_i[0];
  assign { dest_n_0__4_, dest_n_0__3_, dest_n_0__2_, dest_n_0__1_, dest_n_0__0_ } = (N108)? { N284, N283, N282, N281, N280 } :
                                                                                    (N109)? { dest_r_0__4_, dest_r_0__3_, dest_r_0__2_, dest_r_0__1_, dest_r_0__0_ } : 1'b0;
  assign N108 = N395;
  assign N109 = N394;
  assign { N290, N289 } = (N110)? { N288, N287 } :
                          (N286)? { 1'b0, 1'b0 } : 1'b0;
  assign N110 = N285;
  assign { dest_n_1__4_, dest_n_1__3_, dest_n_1__2_, dest_n_1__0_ } = (N111)? { N292, N291, N290, N289 } :
                                                                      (N112)? { dest_r_1__4_, dest_r_1__3_, dest_r_1__2_, dest_r_1__0_ } : 1'b0;
  assign N111 = N393;
  assign N112 = N392;
  assign { dest_n_2__4_, dest_n_2__3_, dest_n_2__1_, dest_n_2__0_ } = (N113)? { N284, N283, N281, N280 } :
                                                                      (N114)? { dest_r_2__4_, dest_r_2__3_, dest_r_2__1_, dest_r_2__0_ } : 1'b0;
  assign N113 = N391;
  assign N114 = N390;
  assign { N300, N299, N298 } = (N115)? { N297, N296, N295 } :
                                (N294)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N115 = N293;
  assign { dest_n_3__4_, dest_n_3__2_, dest_n_3__1_, dest_n_3__0_ } = (N116)? { N301, N300, N299, N298 } :
                                                                      (N117)? { dest_r_3__4_, dest_r_3__2_, dest_r_3__1_, dest_r_3__0_ } : 1'b0;
  assign N116 = N389;
  assign N117 = N388;
  assign { dest_n_4__3_, dest_n_4__2_, dest_n_4__1_, dest_n_4__0_ } = (N118)? { N283, N282, N281, N280 } :
                                                                      (N119)? { dest_r_4__3_, dest_r_4__2_, dest_r_4__1_, dest_r_4__0_ } : 1'b0;
  assign N118 = N387;
  assign N119 = N386;
  assign N120 = ~reset_i;
  assign N121 = reset_i;
  assign N122 = N120;
  assign N123 = ~fifo_yumi_i[0];
  assign N124 = N122 & fifo_yumi_i[0];
  assign N133 = ~reset_i;
  assign N134 = reset_i;
  assign N135 = N133;
  assign N136 = fifo_yumi_i[1];
  assign N137 = ~N136;
  assign N138 = N135 & N136;
  assign N147 = ~reset_i;
  assign N148 = reset_i;
  assign N149 = N147;
  assign N150 = ~fifo_yumi_i[2];
  assign N151 = N149 & fifo_yumi_i[2];
  assign N160 = ~reset_i;
  assign N161 = reset_i;
  assign N162 = N160;
  assign N163 = fifo_yumi_i[3];
  assign N164 = ~N163;
  assign N165 = N162 & N163;
  assign N174 = ~reset_i;
  assign N175 = reset_i;
  assign N176 = N174;
  assign N177 = ~fifo_yumi_i[4];
  assign N178 = N176 & fifo_yumi_i[4];
  assign new_valid_0__0_ = 1'b0 & dest_n_0__0_;
  assign new_valid_0__1_ = 1'b0 & dest_n_0__1_;
  assign new_valid_0__2_ = 1'b0 & dest_n_0__2_;
  assign new_valid_0__3_ = 1'b0 & dest_n_0__3_;
  assign new_valid_0__4_ = 1'b0 & dest_n_0__4_;
  assign new_valid_1__0_ = fifo_valid_o_1 & dest_n_1__0_;
  assign new_valid_1__2_ = fifo_valid_o_1 & dest_n_1__2_;
  assign new_valid_1__3_ = fifo_valid_o_1 & dest_n_1__3_;
  assign new_valid_1__4_ = fifo_valid_o_1 & dest_n_1__4_;
  assign new_valid_2__0_ = 1'b0 & dest_n_2__0_;
  assign new_valid_2__1_ = 1'b0 & dest_n_2__1_;
  assign new_valid_2__3_ = 1'b0 & dest_n_2__3_;
  assign new_valid_2__4_ = 1'b0 & dest_n_2__4_;
  assign new_valid_3__0_ = fifo_valid_o[3] & dest_n_3__0_;
  assign new_valid_3__1_ = fifo_valid_o[3] & dest_n_3__1_;
  assign new_valid_3__2_ = fifo_valid_o[3] & dest_n_3__2_;
  assign new_valid_3__4_ = fifo_valid_o[3] & dest_n_3__4_;
  assign new_valid_4__0_ = 1'b0 & dest_n_4__0_;
  assign new_valid_4__1_ = 1'b0 & dest_n_4__1_;
  assign new_valid_4__2_ = 1'b0 & dest_n_4__2_;
  assign new_valid_4__3_ = 1'b0 & dest_n_4__3_;
  assign fifo_yumi_i[0] = N420 | arb_grants_o_0__0_;
  assign N420 = N419 | arb_grants_o_0__1_;
  assign N419 = N418 | arb_grants_o_0__2_;
  assign N418 = arb_grants_o_0__4_ | arb_grants_o_0__3_;
  assign fifo_yumi_i[1] = N423 | arb_grants_o_1__0_;
  assign N423 = N422 | 1'b0;
  assign N422 = N421 | arb_grants_o_1__2_;
  assign N421 = arb_grants_o_1__4_ | arb_grants_o_1__3_;
  assign fifo_yumi_i[2] = N426 | arb_grants_o_2__0_;
  assign N426 = N425 | arb_grants_o_2__1_;
  assign N425 = N424 | 1'b0;
  assign N424 = arb_grants_o_2__4_ | arb_grants_o_2__3_;
  assign fifo_yumi_i[3] = N429 | arb_grants_o_3__0_;
  assign N429 = N428 | arb_grants_o_3__1_;
  assign N428 = N427 | arb_grants_o_3__2_;
  assign N427 = arb_grants_o_3__4_ | 1'b0;
  assign fifo_yumi_i[4] = N432 | arb_grants_o_4__0_;
  assign N432 = N431 | arb_grants_o_4__1_;
  assign N431 = N430 | arb_grants_o_4__2_;
  assign N430 = 1'b0 | arb_grants_o_4__3_;
  assign N187 = ~reset_i;
  assign N188 = reset_i;
  assign N189 = N187;
  assign N190 = valid_o[0] & ready_i[0];
  assign N191 = ~N190;
  assign N192 = N189 & N190;
  assign N201 = ~reset_i;
  assign N202 = reset_i;
  assign N203 = N201;
  assign N204 = valid_o[1] & ready_i[1];
  assign N205 = ~N204;
  assign N206 = N203 & N204;
  assign N215 = ~reset_i;
  assign N216 = reset_i;
  assign N217 = N215;
  assign N218 = valid_o[2] & 1'b1;
  assign N219 = ~N218;
  assign N220 = N217 & N218;
  assign N229 = ~reset_i;
  assign N230 = reset_i;
  assign N231 = N229;
  assign N232 = valid_o[3] & 1'b1;
  assign N233 = ~N232;
  assign N234 = N231 & N232;
  assign N243 = ~reset_i;
  assign N244 = reset_i;
  assign N245 = N243;
  assign N246 = valid_o[4] & 1'b1;
  assign N247 = ~N246;
  assign N248 = N245 & N246;
  assign N257 = new_valid_0__0_ & arb_grants_r_0__0_;
  assign N258 = new_valid_0__1_ & arb_grants_r_0__1_;
  assign N259 = new_valid_0__2_ & arb_grants_r_0__2_;
  assign N260 = new_valid_0__3_ & arb_grants_r_0__3_;
  assign N261 = new_valid_0__4_ & arb_grants_r_0__4_;
  assign N262 = new_valid_1__0_ & arb_grants_r_1__0_;
  assign N263 = new_valid_1__2_ & arb_grants_r_1__2_;
  assign N264 = new_valid_1__3_ & arb_grants_r_1__3_;
  assign N265 = new_valid_1__4_ & arb_grants_r_1__4_;
  assign N266 = new_valid_2__0_ & arb_grants_r_2__0_;
  assign N267 = new_valid_2__1_ & arb_grants_r_2__1_;
  assign N268 = new_valid_2__3_ & arb_grants_r_2__3_;
  assign N269 = new_valid_2__4_ & arb_grants_r_2__4_;
  assign N270 = new_valid_3__0_ & arb_grants_r_3__0_;
  assign N271 = new_valid_3__1_ & arb_grants_r_3__1_;
  assign N272 = new_valid_3__2_ & arb_grants_r_3__2_;
  assign N273 = new_valid_3__4_ & arb_grants_r_3__4_;
  assign N274 = new_valid_4__0_ & arb_grants_r_4__0_;
  assign N275 = new_valid_4__1_ & arb_grants_r_4__1_;
  assign N276 = new_valid_4__2_ & arb_grants_r_4__2_;
  assign N277 = new_valid_4__3_ & arb_grants_r_4__3_;
  assign n_3_net_ = valid_o[1] & ready_i[1];
  assign n_9_net_ = valid_o[2] & 1'b1;
  assign n_15_net_ = valid_o[3] & 1'b1;
  assign n_21_net_ = valid_o[4] & 1'b1;
  assign n_27_net_ = valid_o[0] & ready_i[0];
  assign N286 = ~N285;
  assign N294 = ~N293;
  assign N302 = ~N365;
  assign N303 = ~N366;
  assign N304 = ~N367;
  assign N305 = ~N368;
  assign N306 = ~N369;
  assign N307 = ~N370;
  assign N308 = ~N371;
  assign N309 = ~N372;
  assign N310 = ~N373;
  assign N311 = ~N374;
  assign N312 = ~N375;
  assign N313 = ~N376;
  assign N314 = ~N377;
  assign N315 = ~N378;
  assign N316 = ~N379;
  assign N317 = ~N380;
  assign N318 = ~N381;
  assign N319 = ~N382;
  assign N320 = ~N383;
  assign N321 = ~N384;
  assign N322 = ~N385;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { count_r[9:0] } <= { N186, N185, N173, N172, N159, N158, N146, N145, N132, N131 };
      dest_r_0__4_ <= dest_n_0__4_;
      dest_r_0__3_ <= dest_n_0__3_;
      dest_r_0__2_ <= dest_n_0__2_;
      dest_r_0__1_ <= dest_n_0__1_;
      dest_r_0__0_ <= dest_n_0__0_;
      dest_r_1__4_ <= dest_n_1__4_;
      dest_r_1__3_ <= dest_n_1__3_;
      dest_r_1__2_ <= dest_n_1__2_;
      dest_r_1__0_ <= dest_n_1__0_;
      dest_r_2__4_ <= dest_n_2__4_;
      dest_r_2__3_ <= dest_n_2__3_;
      dest_r_2__1_ <= dest_n_2__1_;
      dest_r_2__0_ <= dest_n_2__0_;
      dest_r_3__4_ <= dest_n_3__4_;
      dest_r_3__2_ <= dest_n_3__2_;
      dest_r_3__1_ <= dest_n_3__1_;
      dest_r_3__0_ <= dest_n_3__0_;
      dest_r_4__3_ <= dest_n_4__3_;
      dest_r_4__2_ <= dest_n_4__2_;
      dest_r_4__1_ <= dest_n_4__1_;
      dest_r_4__0_ <= dest_n_4__0_;
      { out_count_r[9:0] } <= { N256, N255, N242, N241, N228, N227, N214, N213, N200, N199 };
    end
    if(N302) begin
      arb_grants_r_0__0_ <= arb_grants_o_0__0_;
    end
    if(N303) begin
      arb_grants_r_0__1_ <= arb_grants_o_0__1_;
    end
    if(N304) begin
      arb_grants_r_0__2_ <= arb_grants_o_0__2_;
    end
    if(N305) begin
      arb_grants_r_0__3_ <= arb_grants_o_0__3_;
    end
    if(N306) begin
      arb_grants_r_0__4_ <= arb_grants_o_0__4_;
    end
    if(N307) begin
      arb_grants_r_1__0_ <= arb_grants_o_1__0_;
    end
    if(N308) begin
      arb_grants_r_1__2_ <= arb_grants_o_1__2_;
    end
    if(N309) begin
      arb_grants_r_1__3_ <= arb_grants_o_1__3_;
    end
    if(N310) begin
      arb_grants_r_1__4_ <= arb_grants_o_1__4_;
    end
    if(N311) begin
      arb_grants_r_2__0_ <= arb_grants_o_2__0_;
    end
    if(N312) begin
      arb_grants_r_2__1_ <= arb_grants_o_2__1_;
    end
    if(N313) begin
      arb_grants_r_2__3_ <= arb_grants_o_2__3_;
    end
    if(N314) begin
      arb_grants_r_2__4_ <= arb_grants_o_2__4_;
    end
    if(N315) begin
      arb_grants_r_3__0_ <= arb_grants_o_3__0_;
    end
    if(N316) begin
      arb_grants_r_3__1_ <= arb_grants_o_3__1_;
    end
    if(N317) begin
      arb_grants_r_3__2_ <= arb_grants_o_3__2_;
    end
    if(N318) begin
      arb_grants_r_3__4_ <= arb_grants_o_3__4_;
    end
    if(N319) begin
      arb_grants_r_4__0_ <= arb_grants_o_4__0_;
    end
    if(N320) begin
      arb_grants_r_4__1_ <= arb_grants_o_4__1_;
    end
    if(N321) begin
      arb_grants_r_4__2_ <= arb_grants_o_4__2_;
    end
    if(N322) begin
      arb_grants_r_4__3_ <= arb_grants_o_4__3_;
    end
  end


endmodule



module bp_me_network_pkt_encode_data_resp_num_lce_p2_num_cce_p1_paddr_width_p22_block_size_in_bits_p512_max_num_flit_p4_x_cord_width_p1_y_cord_width_p1
(
  payload_i,
  packet_o
);

  input [536:0] payload_i;
  output [540:0] packet_o;
  wire [540:0] packet_o;
  wire N0;
  assign packet_o[1] = 1'b0;
  assign packet_o[2] = packet_o[3];
  assign packet_o[540] = payload_i[536];
  assign packet_o[539] = payload_i[535];
  assign packet_o[538] = payload_i[534];
  assign packet_o[537] = payload_i[533];
  assign packet_o[536] = payload_i[532];
  assign packet_o[535] = payload_i[531];
  assign packet_o[534] = payload_i[530];
  assign packet_o[533] = payload_i[529];
  assign packet_o[532] = payload_i[528];
  assign packet_o[531] = payload_i[527];
  assign packet_o[530] = payload_i[526];
  assign packet_o[529] = payload_i[525];
  assign packet_o[528] = payload_i[524];
  assign packet_o[527] = payload_i[523];
  assign packet_o[526] = payload_i[522];
  assign packet_o[525] = payload_i[521];
  assign packet_o[524] = payload_i[520];
  assign packet_o[523] = payload_i[519];
  assign packet_o[522] = payload_i[518];
  assign packet_o[521] = payload_i[517];
  assign packet_o[520] = payload_i[516];
  assign packet_o[519] = payload_i[515];
  assign packet_o[518] = payload_i[514];
  assign packet_o[517] = payload_i[513];
  assign packet_o[516] = payload_i[512];
  assign packet_o[515] = payload_i[511];
  assign packet_o[514] = payload_i[510];
  assign packet_o[513] = payload_i[509];
  assign packet_o[512] = payload_i[508];
  assign packet_o[511] = payload_i[507];
  assign packet_o[510] = payload_i[506];
  assign packet_o[509] = payload_i[505];
  assign packet_o[508] = payload_i[504];
  assign packet_o[507] = payload_i[503];
  assign packet_o[506] = payload_i[502];
  assign packet_o[505] = payload_i[501];
  assign packet_o[504] = payload_i[500];
  assign packet_o[503] = payload_i[499];
  assign packet_o[502] = payload_i[498];
  assign packet_o[501] = payload_i[497];
  assign packet_o[500] = payload_i[496];
  assign packet_o[499] = payload_i[495];
  assign packet_o[498] = payload_i[494];
  assign packet_o[497] = payload_i[493];
  assign packet_o[496] = payload_i[492];
  assign packet_o[495] = payload_i[491];
  assign packet_o[494] = payload_i[490];
  assign packet_o[493] = payload_i[489];
  assign packet_o[492] = payload_i[488];
  assign packet_o[491] = payload_i[487];
  assign packet_o[490] = payload_i[486];
  assign packet_o[489] = payload_i[485];
  assign packet_o[488] = payload_i[484];
  assign packet_o[487] = payload_i[483];
  assign packet_o[486] = payload_i[482];
  assign packet_o[485] = payload_i[481];
  assign packet_o[484] = payload_i[480];
  assign packet_o[483] = payload_i[479];
  assign packet_o[482] = payload_i[478];
  assign packet_o[481] = payload_i[477];
  assign packet_o[480] = payload_i[476];
  assign packet_o[479] = payload_i[475];
  assign packet_o[478] = payload_i[474];
  assign packet_o[477] = payload_i[473];
  assign packet_o[476] = payload_i[472];
  assign packet_o[475] = payload_i[471];
  assign packet_o[474] = payload_i[470];
  assign packet_o[473] = payload_i[469];
  assign packet_o[472] = payload_i[468];
  assign packet_o[471] = payload_i[467];
  assign packet_o[470] = payload_i[466];
  assign packet_o[469] = payload_i[465];
  assign packet_o[468] = payload_i[464];
  assign packet_o[467] = payload_i[463];
  assign packet_o[466] = payload_i[462];
  assign packet_o[465] = payload_i[461];
  assign packet_o[464] = payload_i[460];
  assign packet_o[463] = payload_i[459];
  assign packet_o[462] = payload_i[458];
  assign packet_o[461] = payload_i[457];
  assign packet_o[460] = payload_i[456];
  assign packet_o[459] = payload_i[455];
  assign packet_o[458] = payload_i[454];
  assign packet_o[457] = payload_i[453];
  assign packet_o[456] = payload_i[452];
  assign packet_o[455] = payload_i[451];
  assign packet_o[454] = payload_i[450];
  assign packet_o[453] = payload_i[449];
  assign packet_o[452] = payload_i[448];
  assign packet_o[451] = payload_i[447];
  assign packet_o[450] = payload_i[446];
  assign packet_o[449] = payload_i[445];
  assign packet_o[448] = payload_i[444];
  assign packet_o[447] = payload_i[443];
  assign packet_o[446] = payload_i[442];
  assign packet_o[445] = payload_i[441];
  assign packet_o[444] = payload_i[440];
  assign packet_o[443] = payload_i[439];
  assign packet_o[442] = payload_i[438];
  assign packet_o[441] = payload_i[437];
  assign packet_o[440] = payload_i[436];
  assign packet_o[439] = payload_i[435];
  assign packet_o[438] = payload_i[434];
  assign packet_o[437] = payload_i[433];
  assign packet_o[436] = payload_i[432];
  assign packet_o[435] = payload_i[431];
  assign packet_o[434] = payload_i[430];
  assign packet_o[433] = payload_i[429];
  assign packet_o[432] = payload_i[428];
  assign packet_o[431] = payload_i[427];
  assign packet_o[430] = payload_i[426];
  assign packet_o[429] = payload_i[425];
  assign packet_o[428] = payload_i[424];
  assign packet_o[427] = payload_i[423];
  assign packet_o[426] = payload_i[422];
  assign packet_o[425] = payload_i[421];
  assign packet_o[424] = payload_i[420];
  assign packet_o[423] = payload_i[419];
  assign packet_o[422] = payload_i[418];
  assign packet_o[421] = payload_i[417];
  assign packet_o[420] = payload_i[416];
  assign packet_o[419] = payload_i[415];
  assign packet_o[418] = payload_i[414];
  assign packet_o[417] = payload_i[413];
  assign packet_o[416] = payload_i[412];
  assign packet_o[415] = payload_i[411];
  assign packet_o[414] = payload_i[410];
  assign packet_o[413] = payload_i[409];
  assign packet_o[412] = payload_i[408];
  assign packet_o[411] = payload_i[407];
  assign packet_o[410] = payload_i[406];
  assign packet_o[409] = payload_i[405];
  assign packet_o[408] = payload_i[404];
  assign packet_o[407] = payload_i[403];
  assign packet_o[406] = payload_i[402];
  assign packet_o[405] = payload_i[401];
  assign packet_o[404] = payload_i[400];
  assign packet_o[403] = payload_i[399];
  assign packet_o[402] = payload_i[398];
  assign packet_o[401] = payload_i[397];
  assign packet_o[400] = payload_i[396];
  assign packet_o[399] = payload_i[395];
  assign packet_o[398] = payload_i[394];
  assign packet_o[397] = payload_i[393];
  assign packet_o[396] = payload_i[392];
  assign packet_o[395] = payload_i[391];
  assign packet_o[394] = payload_i[390];
  assign packet_o[393] = payload_i[389];
  assign packet_o[392] = payload_i[388];
  assign packet_o[391] = payload_i[387];
  assign packet_o[390] = payload_i[386];
  assign packet_o[389] = payload_i[385];
  assign packet_o[388] = payload_i[384];
  assign packet_o[387] = payload_i[383];
  assign packet_o[386] = payload_i[382];
  assign packet_o[385] = payload_i[381];
  assign packet_o[384] = payload_i[380];
  assign packet_o[383] = payload_i[379];
  assign packet_o[382] = payload_i[378];
  assign packet_o[381] = payload_i[377];
  assign packet_o[380] = payload_i[376];
  assign packet_o[379] = payload_i[375];
  assign packet_o[378] = payload_i[374];
  assign packet_o[377] = payload_i[373];
  assign packet_o[376] = payload_i[372];
  assign packet_o[375] = payload_i[371];
  assign packet_o[374] = payload_i[370];
  assign packet_o[373] = payload_i[369];
  assign packet_o[372] = payload_i[368];
  assign packet_o[371] = payload_i[367];
  assign packet_o[370] = payload_i[366];
  assign packet_o[369] = payload_i[365];
  assign packet_o[368] = payload_i[364];
  assign packet_o[367] = payload_i[363];
  assign packet_o[366] = payload_i[362];
  assign packet_o[365] = payload_i[361];
  assign packet_o[364] = payload_i[360];
  assign packet_o[363] = payload_i[359];
  assign packet_o[362] = payload_i[358];
  assign packet_o[361] = payload_i[357];
  assign packet_o[360] = payload_i[356];
  assign packet_o[359] = payload_i[355];
  assign packet_o[358] = payload_i[354];
  assign packet_o[357] = payload_i[353];
  assign packet_o[356] = payload_i[352];
  assign packet_o[355] = payload_i[351];
  assign packet_o[354] = payload_i[350];
  assign packet_o[353] = payload_i[349];
  assign packet_o[352] = payload_i[348];
  assign packet_o[351] = payload_i[347];
  assign packet_o[350] = payload_i[346];
  assign packet_o[349] = payload_i[345];
  assign packet_o[348] = payload_i[344];
  assign packet_o[347] = payload_i[343];
  assign packet_o[346] = payload_i[342];
  assign packet_o[345] = payload_i[341];
  assign packet_o[344] = payload_i[340];
  assign packet_o[343] = payload_i[339];
  assign packet_o[342] = payload_i[338];
  assign packet_o[341] = payload_i[337];
  assign packet_o[340] = payload_i[336];
  assign packet_o[339] = payload_i[335];
  assign packet_o[338] = payload_i[334];
  assign packet_o[337] = payload_i[333];
  assign packet_o[336] = payload_i[332];
  assign packet_o[335] = payload_i[331];
  assign packet_o[334] = payload_i[330];
  assign packet_o[333] = payload_i[329];
  assign packet_o[332] = payload_i[328];
  assign packet_o[331] = payload_i[327];
  assign packet_o[330] = payload_i[326];
  assign packet_o[329] = payload_i[325];
  assign packet_o[328] = payload_i[324];
  assign packet_o[327] = payload_i[323];
  assign packet_o[326] = payload_i[322];
  assign packet_o[325] = payload_i[321];
  assign packet_o[324] = payload_i[320];
  assign packet_o[323] = payload_i[319];
  assign packet_o[322] = payload_i[318];
  assign packet_o[321] = payload_i[317];
  assign packet_o[320] = payload_i[316];
  assign packet_o[319] = payload_i[315];
  assign packet_o[318] = payload_i[314];
  assign packet_o[317] = payload_i[313];
  assign packet_o[316] = payload_i[312];
  assign packet_o[315] = payload_i[311];
  assign packet_o[314] = payload_i[310];
  assign packet_o[313] = payload_i[309];
  assign packet_o[312] = payload_i[308];
  assign packet_o[311] = payload_i[307];
  assign packet_o[310] = payload_i[306];
  assign packet_o[309] = payload_i[305];
  assign packet_o[308] = payload_i[304];
  assign packet_o[307] = payload_i[303];
  assign packet_o[306] = payload_i[302];
  assign packet_o[305] = payload_i[301];
  assign packet_o[304] = payload_i[300];
  assign packet_o[303] = payload_i[299];
  assign packet_o[302] = payload_i[298];
  assign packet_o[301] = payload_i[297];
  assign packet_o[300] = payload_i[296];
  assign packet_o[299] = payload_i[295];
  assign packet_o[298] = payload_i[294];
  assign packet_o[297] = payload_i[293];
  assign packet_o[296] = payload_i[292];
  assign packet_o[295] = payload_i[291];
  assign packet_o[294] = payload_i[290];
  assign packet_o[293] = payload_i[289];
  assign packet_o[292] = payload_i[288];
  assign packet_o[291] = payload_i[287];
  assign packet_o[290] = payload_i[286];
  assign packet_o[289] = payload_i[285];
  assign packet_o[288] = payload_i[284];
  assign packet_o[287] = payload_i[283];
  assign packet_o[286] = payload_i[282];
  assign packet_o[285] = payload_i[281];
  assign packet_o[284] = payload_i[280];
  assign packet_o[283] = payload_i[279];
  assign packet_o[282] = payload_i[278];
  assign packet_o[281] = payload_i[277];
  assign packet_o[280] = payload_i[276];
  assign packet_o[279] = payload_i[275];
  assign packet_o[278] = payload_i[274];
  assign packet_o[277] = payload_i[273];
  assign packet_o[276] = payload_i[272];
  assign packet_o[275] = payload_i[271];
  assign packet_o[274] = payload_i[270];
  assign packet_o[273] = payload_i[269];
  assign packet_o[272] = payload_i[268];
  assign packet_o[271] = payload_i[267];
  assign packet_o[270] = payload_i[266];
  assign packet_o[269] = payload_i[265];
  assign packet_o[268] = payload_i[264];
  assign packet_o[267] = payload_i[263];
  assign packet_o[266] = payload_i[262];
  assign packet_o[265] = payload_i[261];
  assign packet_o[264] = payload_i[260];
  assign packet_o[263] = payload_i[259];
  assign packet_o[262] = payload_i[258];
  assign packet_o[261] = payload_i[257];
  assign packet_o[260] = payload_i[256];
  assign packet_o[259] = payload_i[255];
  assign packet_o[258] = payload_i[254];
  assign packet_o[257] = payload_i[253];
  assign packet_o[256] = payload_i[252];
  assign packet_o[255] = payload_i[251];
  assign packet_o[254] = payload_i[250];
  assign packet_o[253] = payload_i[249];
  assign packet_o[252] = payload_i[248];
  assign packet_o[251] = payload_i[247];
  assign packet_o[250] = payload_i[246];
  assign packet_o[249] = payload_i[245];
  assign packet_o[248] = payload_i[244];
  assign packet_o[247] = payload_i[243];
  assign packet_o[246] = payload_i[242];
  assign packet_o[245] = payload_i[241];
  assign packet_o[244] = payload_i[240];
  assign packet_o[243] = payload_i[239];
  assign packet_o[242] = payload_i[238];
  assign packet_o[241] = payload_i[237];
  assign packet_o[240] = payload_i[236];
  assign packet_o[239] = payload_i[235];
  assign packet_o[238] = payload_i[234];
  assign packet_o[237] = payload_i[233];
  assign packet_o[236] = payload_i[232];
  assign packet_o[235] = payload_i[231];
  assign packet_o[234] = payload_i[230];
  assign packet_o[233] = payload_i[229];
  assign packet_o[232] = payload_i[228];
  assign packet_o[231] = payload_i[227];
  assign packet_o[230] = payload_i[226];
  assign packet_o[229] = payload_i[225];
  assign packet_o[228] = payload_i[224];
  assign packet_o[227] = payload_i[223];
  assign packet_o[226] = payload_i[222];
  assign packet_o[225] = payload_i[221];
  assign packet_o[224] = payload_i[220];
  assign packet_o[223] = payload_i[219];
  assign packet_o[222] = payload_i[218];
  assign packet_o[221] = payload_i[217];
  assign packet_o[220] = payload_i[216];
  assign packet_o[219] = payload_i[215];
  assign packet_o[218] = payload_i[214];
  assign packet_o[217] = payload_i[213];
  assign packet_o[216] = payload_i[212];
  assign packet_o[215] = payload_i[211];
  assign packet_o[214] = payload_i[210];
  assign packet_o[213] = payload_i[209];
  assign packet_o[212] = payload_i[208];
  assign packet_o[211] = payload_i[207];
  assign packet_o[210] = payload_i[206];
  assign packet_o[209] = payload_i[205];
  assign packet_o[208] = payload_i[204];
  assign packet_o[207] = payload_i[203];
  assign packet_o[206] = payload_i[202];
  assign packet_o[205] = payload_i[201];
  assign packet_o[204] = payload_i[200];
  assign packet_o[203] = payload_i[199];
  assign packet_o[202] = payload_i[198];
  assign packet_o[201] = payload_i[197];
  assign packet_o[200] = payload_i[196];
  assign packet_o[199] = payload_i[195];
  assign packet_o[198] = payload_i[194];
  assign packet_o[197] = payload_i[193];
  assign packet_o[196] = payload_i[192];
  assign packet_o[195] = payload_i[191];
  assign packet_o[194] = payload_i[190];
  assign packet_o[193] = payload_i[189];
  assign packet_o[192] = payload_i[188];
  assign packet_o[191] = payload_i[187];
  assign packet_o[190] = payload_i[186];
  assign packet_o[189] = payload_i[185];
  assign packet_o[188] = payload_i[184];
  assign packet_o[187] = payload_i[183];
  assign packet_o[186] = payload_i[182];
  assign packet_o[185] = payload_i[181];
  assign packet_o[184] = payload_i[180];
  assign packet_o[183] = payload_i[179];
  assign packet_o[182] = payload_i[178];
  assign packet_o[181] = payload_i[177];
  assign packet_o[180] = payload_i[176];
  assign packet_o[179] = payload_i[175];
  assign packet_o[178] = payload_i[174];
  assign packet_o[177] = payload_i[173];
  assign packet_o[176] = payload_i[172];
  assign packet_o[175] = payload_i[171];
  assign packet_o[174] = payload_i[170];
  assign packet_o[173] = payload_i[169];
  assign packet_o[172] = payload_i[168];
  assign packet_o[171] = payload_i[167];
  assign packet_o[170] = payload_i[166];
  assign packet_o[169] = payload_i[165];
  assign packet_o[168] = payload_i[164];
  assign packet_o[167] = payload_i[163];
  assign packet_o[166] = payload_i[162];
  assign packet_o[165] = payload_i[161];
  assign packet_o[164] = payload_i[160];
  assign packet_o[163] = payload_i[159];
  assign packet_o[162] = payload_i[158];
  assign packet_o[161] = payload_i[157];
  assign packet_o[160] = payload_i[156];
  assign packet_o[159] = payload_i[155];
  assign packet_o[158] = payload_i[154];
  assign packet_o[157] = payload_i[153];
  assign packet_o[156] = payload_i[152];
  assign packet_o[155] = payload_i[151];
  assign packet_o[154] = payload_i[150];
  assign packet_o[153] = payload_i[149];
  assign packet_o[152] = payload_i[148];
  assign packet_o[151] = payload_i[147];
  assign packet_o[150] = payload_i[146];
  assign packet_o[149] = payload_i[145];
  assign packet_o[148] = payload_i[144];
  assign packet_o[147] = payload_i[143];
  assign packet_o[146] = payload_i[142];
  assign packet_o[145] = payload_i[141];
  assign packet_o[144] = payload_i[140];
  assign packet_o[143] = payload_i[139];
  assign packet_o[142] = payload_i[138];
  assign packet_o[141] = payload_i[137];
  assign packet_o[140] = payload_i[136];
  assign packet_o[139] = payload_i[135];
  assign packet_o[138] = payload_i[134];
  assign packet_o[137] = payload_i[133];
  assign packet_o[136] = payload_i[132];
  assign packet_o[135] = payload_i[131];
  assign packet_o[134] = payload_i[130];
  assign packet_o[133] = payload_i[129];
  assign packet_o[132] = payload_i[128];
  assign packet_o[131] = payload_i[127];
  assign packet_o[130] = payload_i[126];
  assign packet_o[129] = payload_i[125];
  assign packet_o[128] = payload_i[124];
  assign packet_o[127] = payload_i[123];
  assign packet_o[126] = payload_i[122];
  assign packet_o[125] = payload_i[121];
  assign packet_o[124] = payload_i[120];
  assign packet_o[123] = payload_i[119];
  assign packet_o[122] = payload_i[118];
  assign packet_o[121] = payload_i[117];
  assign packet_o[120] = payload_i[116];
  assign packet_o[119] = payload_i[115];
  assign packet_o[118] = payload_i[114];
  assign packet_o[117] = payload_i[113];
  assign packet_o[116] = payload_i[112];
  assign packet_o[115] = payload_i[111];
  assign packet_o[114] = payload_i[110];
  assign packet_o[113] = payload_i[109];
  assign packet_o[112] = payload_i[108];
  assign packet_o[111] = payload_i[107];
  assign packet_o[110] = payload_i[106];
  assign packet_o[109] = payload_i[105];
  assign packet_o[108] = payload_i[104];
  assign packet_o[107] = payload_i[103];
  assign packet_o[106] = payload_i[102];
  assign packet_o[105] = payload_i[101];
  assign packet_o[104] = payload_i[100];
  assign packet_o[103] = payload_i[99];
  assign packet_o[102] = payload_i[98];
  assign packet_o[101] = payload_i[97];
  assign packet_o[100] = payload_i[96];
  assign packet_o[99] = payload_i[95];
  assign packet_o[98] = payload_i[94];
  assign packet_o[97] = payload_i[93];
  assign packet_o[96] = payload_i[92];
  assign packet_o[95] = payload_i[91];
  assign packet_o[94] = payload_i[90];
  assign packet_o[93] = payload_i[89];
  assign packet_o[92] = payload_i[88];
  assign packet_o[91] = payload_i[87];
  assign packet_o[90] = payload_i[86];
  assign packet_o[89] = payload_i[85];
  assign packet_o[88] = payload_i[84];
  assign packet_o[87] = payload_i[83];
  assign packet_o[86] = payload_i[82];
  assign packet_o[85] = payload_i[81];
  assign packet_o[84] = payload_i[80];
  assign packet_o[83] = payload_i[79];
  assign packet_o[82] = payload_i[78];
  assign packet_o[81] = payload_i[77];
  assign packet_o[80] = payload_i[76];
  assign packet_o[79] = payload_i[75];
  assign packet_o[78] = payload_i[74];
  assign packet_o[77] = payload_i[73];
  assign packet_o[76] = payload_i[72];
  assign packet_o[75] = payload_i[71];
  assign packet_o[74] = payload_i[70];
  assign packet_o[73] = payload_i[69];
  assign packet_o[72] = payload_i[68];
  assign packet_o[71] = payload_i[67];
  assign packet_o[70] = payload_i[66];
  assign packet_o[69] = payload_i[65];
  assign packet_o[68] = payload_i[64];
  assign packet_o[67] = payload_i[63];
  assign packet_o[66] = payload_i[62];
  assign packet_o[65] = payload_i[61];
  assign packet_o[64] = payload_i[60];
  assign packet_o[63] = payload_i[59];
  assign packet_o[62] = payload_i[58];
  assign packet_o[61] = payload_i[57];
  assign packet_o[60] = payload_i[56];
  assign packet_o[59] = payload_i[55];
  assign packet_o[58] = payload_i[54];
  assign packet_o[57] = payload_i[53];
  assign packet_o[56] = payload_i[52];
  assign packet_o[55] = payload_i[51];
  assign packet_o[54] = payload_i[50];
  assign packet_o[53] = payload_i[49];
  assign packet_o[52] = payload_i[48];
  assign packet_o[51] = payload_i[47];
  assign packet_o[50] = payload_i[46];
  assign packet_o[49] = payload_i[45];
  assign packet_o[48] = payload_i[44];
  assign packet_o[47] = payload_i[43];
  assign packet_o[46] = payload_i[42];
  assign packet_o[45] = payload_i[41];
  assign packet_o[44] = payload_i[40];
  assign packet_o[43] = payload_i[39];
  assign packet_o[42] = payload_i[38];
  assign packet_o[41] = payload_i[37];
  assign packet_o[40] = payload_i[36];
  assign packet_o[39] = payload_i[35];
  assign packet_o[38] = payload_i[34];
  assign packet_o[37] = payload_i[33];
  assign packet_o[36] = payload_i[32];
  assign packet_o[35] = payload_i[31];
  assign packet_o[34] = payload_i[30];
  assign packet_o[33] = payload_i[29];
  assign packet_o[32] = payload_i[28];
  assign packet_o[31] = payload_i[27];
  assign packet_o[30] = payload_i[26];
  assign packet_o[29] = payload_i[25];
  assign packet_o[0] = payload_i[24];
  assign packet_o[28] = payload_i[24];
  assign packet_o[27] = payload_i[23];
  assign packet_o[26] = payload_i[22];
  assign packet_o[25] = payload_i[21];
  assign packet_o[24] = payload_i[20];
  assign packet_o[23] = payload_i[19];
  assign packet_o[22] = payload_i[18];
  assign packet_o[21] = payload_i[17];
  assign packet_o[20] = payload_i[16];
  assign packet_o[19] = payload_i[15];
  assign packet_o[18] = payload_i[14];
  assign packet_o[17] = payload_i[13];
  assign packet_o[16] = payload_i[12];
  assign packet_o[15] = payload_i[11];
  assign packet_o[14] = payload_i[10];
  assign packet_o[13] = payload_i[9];
  assign packet_o[12] = payload_i[8];
  assign packet_o[11] = payload_i[7];
  assign packet_o[10] = payload_i[6];
  assign packet_o[9] = payload_i[5];
  assign packet_o[8] = payload_i[4];
  assign packet_o[7] = payload_i[3];
  assign packet_o[6] = payload_i[2];
  assign packet_o[5] = payload_i[1];
  assign packet_o[4] = payload_i[0];
  assign N0 = ~payload_i[22];
  assign packet_o[3] = N0;

endmodule



module bsg_mux_width_p136_els_p4
(
  data_i,
  sel_i,
  data_o
);

  input [543:0] data_i;
  input [1:0] sel_i;
  output [135:0] data_o;
  wire [135:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[135] = (N2)? data_i[135] :
                       (N4)? data_i[271] :
                       (N3)? data_i[407] :
                       (N5)? data_i[543] : 1'b0;
  assign data_o[134] = (N2)? data_i[134] :
                       (N4)? data_i[270] :
                       (N3)? data_i[406] :
                       (N5)? data_i[542] : 1'b0;
  assign data_o[133] = (N2)? data_i[133] :
                       (N4)? data_i[269] :
                       (N3)? data_i[405] :
                       (N5)? data_i[541] : 1'b0;
  assign data_o[132] = (N2)? data_i[132] :
                       (N4)? data_i[268] :
                       (N3)? data_i[404] :
                       (N5)? data_i[540] : 1'b0;
  assign data_o[131] = (N2)? data_i[131] :
                       (N4)? data_i[267] :
                       (N3)? data_i[403] :
                       (N5)? data_i[539] : 1'b0;
  assign data_o[130] = (N2)? data_i[130] :
                       (N4)? data_i[266] :
                       (N3)? data_i[402] :
                       (N5)? data_i[538] : 1'b0;
  assign data_o[129] = (N2)? data_i[129] :
                       (N4)? data_i[265] :
                       (N3)? data_i[401] :
                       (N5)? data_i[537] : 1'b0;
  assign data_o[128] = (N2)? data_i[128] :
                       (N4)? data_i[264] :
                       (N3)? data_i[400] :
                       (N5)? data_i[536] : 1'b0;
  assign data_o[127] = (N2)? data_i[127] :
                       (N4)? data_i[263] :
                       (N3)? data_i[399] :
                       (N5)? data_i[535] : 1'b0;
  assign data_o[126] = (N2)? data_i[126] :
                       (N4)? data_i[262] :
                       (N3)? data_i[398] :
                       (N5)? data_i[534] : 1'b0;
  assign data_o[125] = (N2)? data_i[125] :
                       (N4)? data_i[261] :
                       (N3)? data_i[397] :
                       (N5)? data_i[533] : 1'b0;
  assign data_o[124] = (N2)? data_i[124] :
                       (N4)? data_i[260] :
                       (N3)? data_i[396] :
                       (N5)? data_i[532] : 1'b0;
  assign data_o[123] = (N2)? data_i[123] :
                       (N4)? data_i[259] :
                       (N3)? data_i[395] :
                       (N5)? data_i[531] : 1'b0;
  assign data_o[122] = (N2)? data_i[122] :
                       (N4)? data_i[258] :
                       (N3)? data_i[394] :
                       (N5)? data_i[530] : 1'b0;
  assign data_o[121] = (N2)? data_i[121] :
                       (N4)? data_i[257] :
                       (N3)? data_i[393] :
                       (N5)? data_i[529] : 1'b0;
  assign data_o[120] = (N2)? data_i[120] :
                       (N4)? data_i[256] :
                       (N3)? data_i[392] :
                       (N5)? data_i[528] : 1'b0;
  assign data_o[119] = (N2)? data_i[119] :
                       (N4)? data_i[255] :
                       (N3)? data_i[391] :
                       (N5)? data_i[527] : 1'b0;
  assign data_o[118] = (N2)? data_i[118] :
                       (N4)? data_i[254] :
                       (N3)? data_i[390] :
                       (N5)? data_i[526] : 1'b0;
  assign data_o[117] = (N2)? data_i[117] :
                       (N4)? data_i[253] :
                       (N3)? data_i[389] :
                       (N5)? data_i[525] : 1'b0;
  assign data_o[116] = (N2)? data_i[116] :
                       (N4)? data_i[252] :
                       (N3)? data_i[388] :
                       (N5)? data_i[524] : 1'b0;
  assign data_o[115] = (N2)? data_i[115] :
                       (N4)? data_i[251] :
                       (N3)? data_i[387] :
                       (N5)? data_i[523] : 1'b0;
  assign data_o[114] = (N2)? data_i[114] :
                       (N4)? data_i[250] :
                       (N3)? data_i[386] :
                       (N5)? data_i[522] : 1'b0;
  assign data_o[113] = (N2)? data_i[113] :
                       (N4)? data_i[249] :
                       (N3)? data_i[385] :
                       (N5)? data_i[521] : 1'b0;
  assign data_o[112] = (N2)? data_i[112] :
                       (N4)? data_i[248] :
                       (N3)? data_i[384] :
                       (N5)? data_i[520] : 1'b0;
  assign data_o[111] = (N2)? data_i[111] :
                       (N4)? data_i[247] :
                       (N3)? data_i[383] :
                       (N5)? data_i[519] : 1'b0;
  assign data_o[110] = (N2)? data_i[110] :
                       (N4)? data_i[246] :
                       (N3)? data_i[382] :
                       (N5)? data_i[518] : 1'b0;
  assign data_o[109] = (N2)? data_i[109] :
                       (N4)? data_i[245] :
                       (N3)? data_i[381] :
                       (N5)? data_i[517] : 1'b0;
  assign data_o[108] = (N2)? data_i[108] :
                       (N4)? data_i[244] :
                       (N3)? data_i[380] :
                       (N5)? data_i[516] : 1'b0;
  assign data_o[107] = (N2)? data_i[107] :
                       (N4)? data_i[243] :
                       (N3)? data_i[379] :
                       (N5)? data_i[515] : 1'b0;
  assign data_o[106] = (N2)? data_i[106] :
                       (N4)? data_i[242] :
                       (N3)? data_i[378] :
                       (N5)? data_i[514] : 1'b0;
  assign data_o[105] = (N2)? data_i[105] :
                       (N4)? data_i[241] :
                       (N3)? data_i[377] :
                       (N5)? data_i[513] : 1'b0;
  assign data_o[104] = (N2)? data_i[104] :
                       (N4)? data_i[240] :
                       (N3)? data_i[376] :
                       (N5)? data_i[512] : 1'b0;
  assign data_o[103] = (N2)? data_i[103] :
                       (N4)? data_i[239] :
                       (N3)? data_i[375] :
                       (N5)? data_i[511] : 1'b0;
  assign data_o[102] = (N2)? data_i[102] :
                       (N4)? data_i[238] :
                       (N3)? data_i[374] :
                       (N5)? data_i[510] : 1'b0;
  assign data_o[101] = (N2)? data_i[101] :
                       (N4)? data_i[237] :
                       (N3)? data_i[373] :
                       (N5)? data_i[509] : 1'b0;
  assign data_o[100] = (N2)? data_i[100] :
                       (N4)? data_i[236] :
                       (N3)? data_i[372] :
                       (N5)? data_i[508] : 1'b0;
  assign data_o[99] = (N2)? data_i[99] :
                      (N4)? data_i[235] :
                      (N3)? data_i[371] :
                      (N5)? data_i[507] : 1'b0;
  assign data_o[98] = (N2)? data_i[98] :
                      (N4)? data_i[234] :
                      (N3)? data_i[370] :
                      (N5)? data_i[506] : 1'b0;
  assign data_o[97] = (N2)? data_i[97] :
                      (N4)? data_i[233] :
                      (N3)? data_i[369] :
                      (N5)? data_i[505] : 1'b0;
  assign data_o[96] = (N2)? data_i[96] :
                      (N4)? data_i[232] :
                      (N3)? data_i[368] :
                      (N5)? data_i[504] : 1'b0;
  assign data_o[95] = (N2)? data_i[95] :
                      (N4)? data_i[231] :
                      (N3)? data_i[367] :
                      (N5)? data_i[503] : 1'b0;
  assign data_o[94] = (N2)? data_i[94] :
                      (N4)? data_i[230] :
                      (N3)? data_i[366] :
                      (N5)? data_i[502] : 1'b0;
  assign data_o[93] = (N2)? data_i[93] :
                      (N4)? data_i[229] :
                      (N3)? data_i[365] :
                      (N5)? data_i[501] : 1'b0;
  assign data_o[92] = (N2)? data_i[92] :
                      (N4)? data_i[228] :
                      (N3)? data_i[364] :
                      (N5)? data_i[500] : 1'b0;
  assign data_o[91] = (N2)? data_i[91] :
                      (N4)? data_i[227] :
                      (N3)? data_i[363] :
                      (N5)? data_i[499] : 1'b0;
  assign data_o[90] = (N2)? data_i[90] :
                      (N4)? data_i[226] :
                      (N3)? data_i[362] :
                      (N5)? data_i[498] : 1'b0;
  assign data_o[89] = (N2)? data_i[89] :
                      (N4)? data_i[225] :
                      (N3)? data_i[361] :
                      (N5)? data_i[497] : 1'b0;
  assign data_o[88] = (N2)? data_i[88] :
                      (N4)? data_i[224] :
                      (N3)? data_i[360] :
                      (N5)? data_i[496] : 1'b0;
  assign data_o[87] = (N2)? data_i[87] :
                      (N4)? data_i[223] :
                      (N3)? data_i[359] :
                      (N5)? data_i[495] : 1'b0;
  assign data_o[86] = (N2)? data_i[86] :
                      (N4)? data_i[222] :
                      (N3)? data_i[358] :
                      (N5)? data_i[494] : 1'b0;
  assign data_o[85] = (N2)? data_i[85] :
                      (N4)? data_i[221] :
                      (N3)? data_i[357] :
                      (N5)? data_i[493] : 1'b0;
  assign data_o[84] = (N2)? data_i[84] :
                      (N4)? data_i[220] :
                      (N3)? data_i[356] :
                      (N5)? data_i[492] : 1'b0;
  assign data_o[83] = (N2)? data_i[83] :
                      (N4)? data_i[219] :
                      (N3)? data_i[355] :
                      (N5)? data_i[491] : 1'b0;
  assign data_o[82] = (N2)? data_i[82] :
                      (N4)? data_i[218] :
                      (N3)? data_i[354] :
                      (N5)? data_i[490] : 1'b0;
  assign data_o[81] = (N2)? data_i[81] :
                      (N4)? data_i[217] :
                      (N3)? data_i[353] :
                      (N5)? data_i[489] : 1'b0;
  assign data_o[80] = (N2)? data_i[80] :
                      (N4)? data_i[216] :
                      (N3)? data_i[352] :
                      (N5)? data_i[488] : 1'b0;
  assign data_o[79] = (N2)? data_i[79] :
                      (N4)? data_i[215] :
                      (N3)? data_i[351] :
                      (N5)? data_i[487] : 1'b0;
  assign data_o[78] = (N2)? data_i[78] :
                      (N4)? data_i[214] :
                      (N3)? data_i[350] :
                      (N5)? data_i[486] : 1'b0;
  assign data_o[77] = (N2)? data_i[77] :
                      (N4)? data_i[213] :
                      (N3)? data_i[349] :
                      (N5)? data_i[485] : 1'b0;
  assign data_o[76] = (N2)? data_i[76] :
                      (N4)? data_i[212] :
                      (N3)? data_i[348] :
                      (N5)? data_i[484] : 1'b0;
  assign data_o[75] = (N2)? data_i[75] :
                      (N4)? data_i[211] :
                      (N3)? data_i[347] :
                      (N5)? data_i[483] : 1'b0;
  assign data_o[74] = (N2)? data_i[74] :
                      (N4)? data_i[210] :
                      (N3)? data_i[346] :
                      (N5)? data_i[482] : 1'b0;
  assign data_o[73] = (N2)? data_i[73] :
                      (N4)? data_i[209] :
                      (N3)? data_i[345] :
                      (N5)? data_i[481] : 1'b0;
  assign data_o[72] = (N2)? data_i[72] :
                      (N4)? data_i[208] :
                      (N3)? data_i[344] :
                      (N5)? data_i[480] : 1'b0;
  assign data_o[71] = (N2)? data_i[71] :
                      (N4)? data_i[207] :
                      (N3)? data_i[343] :
                      (N5)? data_i[479] : 1'b0;
  assign data_o[70] = (N2)? data_i[70] :
                      (N4)? data_i[206] :
                      (N3)? data_i[342] :
                      (N5)? data_i[478] : 1'b0;
  assign data_o[69] = (N2)? data_i[69] :
                      (N4)? data_i[205] :
                      (N3)? data_i[341] :
                      (N5)? data_i[477] : 1'b0;
  assign data_o[68] = (N2)? data_i[68] :
                      (N4)? data_i[204] :
                      (N3)? data_i[340] :
                      (N5)? data_i[476] : 1'b0;
  assign data_o[67] = (N2)? data_i[67] :
                      (N4)? data_i[203] :
                      (N3)? data_i[339] :
                      (N5)? data_i[475] : 1'b0;
  assign data_o[66] = (N2)? data_i[66] :
                      (N4)? data_i[202] :
                      (N3)? data_i[338] :
                      (N5)? data_i[474] : 1'b0;
  assign data_o[65] = (N2)? data_i[65] :
                      (N4)? data_i[201] :
                      (N3)? data_i[337] :
                      (N5)? data_i[473] : 1'b0;
  assign data_o[64] = (N2)? data_i[64] :
                      (N4)? data_i[200] :
                      (N3)? data_i[336] :
                      (N5)? data_i[472] : 1'b0;
  assign data_o[63] = (N2)? data_i[63] :
                      (N4)? data_i[199] :
                      (N3)? data_i[335] :
                      (N5)? data_i[471] : 1'b0;
  assign data_o[62] = (N2)? data_i[62] :
                      (N4)? data_i[198] :
                      (N3)? data_i[334] :
                      (N5)? data_i[470] : 1'b0;
  assign data_o[61] = (N2)? data_i[61] :
                      (N4)? data_i[197] :
                      (N3)? data_i[333] :
                      (N5)? data_i[469] : 1'b0;
  assign data_o[60] = (N2)? data_i[60] :
                      (N4)? data_i[196] :
                      (N3)? data_i[332] :
                      (N5)? data_i[468] : 1'b0;
  assign data_o[59] = (N2)? data_i[59] :
                      (N4)? data_i[195] :
                      (N3)? data_i[331] :
                      (N5)? data_i[467] : 1'b0;
  assign data_o[58] = (N2)? data_i[58] :
                      (N4)? data_i[194] :
                      (N3)? data_i[330] :
                      (N5)? data_i[466] : 1'b0;
  assign data_o[57] = (N2)? data_i[57] :
                      (N4)? data_i[193] :
                      (N3)? data_i[329] :
                      (N5)? data_i[465] : 1'b0;
  assign data_o[56] = (N2)? data_i[56] :
                      (N4)? data_i[192] :
                      (N3)? data_i[328] :
                      (N5)? data_i[464] : 1'b0;
  assign data_o[55] = (N2)? data_i[55] :
                      (N4)? data_i[191] :
                      (N3)? data_i[327] :
                      (N5)? data_i[463] : 1'b0;
  assign data_o[54] = (N2)? data_i[54] :
                      (N4)? data_i[190] :
                      (N3)? data_i[326] :
                      (N5)? data_i[462] : 1'b0;
  assign data_o[53] = (N2)? data_i[53] :
                      (N4)? data_i[189] :
                      (N3)? data_i[325] :
                      (N5)? data_i[461] : 1'b0;
  assign data_o[52] = (N2)? data_i[52] :
                      (N4)? data_i[188] :
                      (N3)? data_i[324] :
                      (N5)? data_i[460] : 1'b0;
  assign data_o[51] = (N2)? data_i[51] :
                      (N4)? data_i[187] :
                      (N3)? data_i[323] :
                      (N5)? data_i[459] : 1'b0;
  assign data_o[50] = (N2)? data_i[50] :
                      (N4)? data_i[186] :
                      (N3)? data_i[322] :
                      (N5)? data_i[458] : 1'b0;
  assign data_o[49] = (N2)? data_i[49] :
                      (N4)? data_i[185] :
                      (N3)? data_i[321] :
                      (N5)? data_i[457] : 1'b0;
  assign data_o[48] = (N2)? data_i[48] :
                      (N4)? data_i[184] :
                      (N3)? data_i[320] :
                      (N5)? data_i[456] : 1'b0;
  assign data_o[47] = (N2)? data_i[47] :
                      (N4)? data_i[183] :
                      (N3)? data_i[319] :
                      (N5)? data_i[455] : 1'b0;
  assign data_o[46] = (N2)? data_i[46] :
                      (N4)? data_i[182] :
                      (N3)? data_i[318] :
                      (N5)? data_i[454] : 1'b0;
  assign data_o[45] = (N2)? data_i[45] :
                      (N4)? data_i[181] :
                      (N3)? data_i[317] :
                      (N5)? data_i[453] : 1'b0;
  assign data_o[44] = (N2)? data_i[44] :
                      (N4)? data_i[180] :
                      (N3)? data_i[316] :
                      (N5)? data_i[452] : 1'b0;
  assign data_o[43] = (N2)? data_i[43] :
                      (N4)? data_i[179] :
                      (N3)? data_i[315] :
                      (N5)? data_i[451] : 1'b0;
  assign data_o[42] = (N2)? data_i[42] :
                      (N4)? data_i[178] :
                      (N3)? data_i[314] :
                      (N5)? data_i[450] : 1'b0;
  assign data_o[41] = (N2)? data_i[41] :
                      (N4)? data_i[177] :
                      (N3)? data_i[313] :
                      (N5)? data_i[449] : 1'b0;
  assign data_o[40] = (N2)? data_i[40] :
                      (N4)? data_i[176] :
                      (N3)? data_i[312] :
                      (N5)? data_i[448] : 1'b0;
  assign data_o[39] = (N2)? data_i[39] :
                      (N4)? data_i[175] :
                      (N3)? data_i[311] :
                      (N5)? data_i[447] : 1'b0;
  assign data_o[38] = (N2)? data_i[38] :
                      (N4)? data_i[174] :
                      (N3)? data_i[310] :
                      (N5)? data_i[446] : 1'b0;
  assign data_o[37] = (N2)? data_i[37] :
                      (N4)? data_i[173] :
                      (N3)? data_i[309] :
                      (N5)? data_i[445] : 1'b0;
  assign data_o[36] = (N2)? data_i[36] :
                      (N4)? data_i[172] :
                      (N3)? data_i[308] :
                      (N5)? data_i[444] : 1'b0;
  assign data_o[35] = (N2)? data_i[35] :
                      (N4)? data_i[171] :
                      (N3)? data_i[307] :
                      (N5)? data_i[443] : 1'b0;
  assign data_o[34] = (N2)? data_i[34] :
                      (N4)? data_i[170] :
                      (N3)? data_i[306] :
                      (N5)? data_i[442] : 1'b0;
  assign data_o[33] = (N2)? data_i[33] :
                      (N4)? data_i[169] :
                      (N3)? data_i[305] :
                      (N5)? data_i[441] : 1'b0;
  assign data_o[32] = (N2)? data_i[32] :
                      (N4)? data_i[168] :
                      (N3)? data_i[304] :
                      (N5)? data_i[440] : 1'b0;
  assign data_o[31] = (N2)? data_i[31] :
                      (N4)? data_i[167] :
                      (N3)? data_i[303] :
                      (N5)? data_i[439] : 1'b0;
  assign data_o[30] = (N2)? data_i[30] :
                      (N4)? data_i[166] :
                      (N3)? data_i[302] :
                      (N5)? data_i[438] : 1'b0;
  assign data_o[29] = (N2)? data_i[29] :
                      (N4)? data_i[165] :
                      (N3)? data_i[301] :
                      (N5)? data_i[437] : 1'b0;
  assign data_o[28] = (N2)? data_i[28] :
                      (N4)? data_i[164] :
                      (N3)? data_i[300] :
                      (N5)? data_i[436] : 1'b0;
  assign data_o[27] = (N2)? data_i[27] :
                      (N4)? data_i[163] :
                      (N3)? data_i[299] :
                      (N5)? data_i[435] : 1'b0;
  assign data_o[26] = (N2)? data_i[26] :
                      (N4)? data_i[162] :
                      (N3)? data_i[298] :
                      (N5)? data_i[434] : 1'b0;
  assign data_o[25] = (N2)? data_i[25] :
                      (N4)? data_i[161] :
                      (N3)? data_i[297] :
                      (N5)? data_i[433] : 1'b0;
  assign data_o[24] = (N2)? data_i[24] :
                      (N4)? data_i[160] :
                      (N3)? data_i[296] :
                      (N5)? data_i[432] : 1'b0;
  assign data_o[23] = (N2)? data_i[23] :
                      (N4)? data_i[159] :
                      (N3)? data_i[295] :
                      (N5)? data_i[431] : 1'b0;
  assign data_o[22] = (N2)? data_i[22] :
                      (N4)? data_i[158] :
                      (N3)? data_i[294] :
                      (N5)? data_i[430] : 1'b0;
  assign data_o[21] = (N2)? data_i[21] :
                      (N4)? data_i[157] :
                      (N3)? data_i[293] :
                      (N5)? data_i[429] : 1'b0;
  assign data_o[20] = (N2)? data_i[20] :
                      (N4)? data_i[156] :
                      (N3)? data_i[292] :
                      (N5)? data_i[428] : 1'b0;
  assign data_o[19] = (N2)? data_i[19] :
                      (N4)? data_i[155] :
                      (N3)? data_i[291] :
                      (N5)? data_i[427] : 1'b0;
  assign data_o[18] = (N2)? data_i[18] :
                      (N4)? data_i[154] :
                      (N3)? data_i[290] :
                      (N5)? data_i[426] : 1'b0;
  assign data_o[17] = (N2)? data_i[17] :
                      (N4)? data_i[153] :
                      (N3)? data_i[289] :
                      (N5)? data_i[425] : 1'b0;
  assign data_o[16] = (N2)? data_i[16] :
                      (N4)? data_i[152] :
                      (N3)? data_i[288] :
                      (N5)? data_i[424] : 1'b0;
  assign data_o[15] = (N2)? data_i[15] :
                      (N4)? data_i[151] :
                      (N3)? data_i[287] :
                      (N5)? data_i[423] : 1'b0;
  assign data_o[14] = (N2)? data_i[14] :
                      (N4)? data_i[150] :
                      (N3)? data_i[286] :
                      (N5)? data_i[422] : 1'b0;
  assign data_o[13] = (N2)? data_i[13] :
                      (N4)? data_i[149] :
                      (N3)? data_i[285] :
                      (N5)? data_i[421] : 1'b0;
  assign data_o[12] = (N2)? data_i[12] :
                      (N4)? data_i[148] :
                      (N3)? data_i[284] :
                      (N5)? data_i[420] : 1'b0;
  assign data_o[11] = (N2)? data_i[11] :
                      (N4)? data_i[147] :
                      (N3)? data_i[283] :
                      (N5)? data_i[419] : 1'b0;
  assign data_o[10] = (N2)? data_i[10] :
                      (N4)? data_i[146] :
                      (N3)? data_i[282] :
                      (N5)? data_i[418] : 1'b0;
  assign data_o[9] = (N2)? data_i[9] :
                     (N4)? data_i[145] :
                     (N3)? data_i[281] :
                     (N5)? data_i[417] : 1'b0;
  assign data_o[8] = (N2)? data_i[8] :
                     (N4)? data_i[144] :
                     (N3)? data_i[280] :
                     (N5)? data_i[416] : 1'b0;
  assign data_o[7] = (N2)? data_i[7] :
                     (N4)? data_i[143] :
                     (N3)? data_i[279] :
                     (N5)? data_i[415] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] :
                     (N4)? data_i[142] :
                     (N3)? data_i[278] :
                     (N5)? data_i[414] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] :
                     (N4)? data_i[141] :
                     (N3)? data_i[277] :
                     (N5)? data_i[413] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] :
                     (N4)? data_i[140] :
                     (N3)? data_i[276] :
                     (N5)? data_i[412] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] :
                     (N4)? data_i[139] :
                     (N3)? data_i[275] :
                     (N5)? data_i[411] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] :
                     (N4)? data_i[138] :
                     (N3)? data_i[274] :
                     (N5)? data_i[410] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] :
                     (N4)? data_i[137] :
                     (N3)? data_i[273] :
                     (N5)? data_i[409] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] :
                     (N4)? data_i[136] :
                     (N3)? data_i[272] :
                     (N5)? data_i[408] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_wormhole_router_adapter_in_max_num_flit_p4_max_payload_width_p537_x_cord_width_p1_y_cord_width_p1
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  ready_o,
  data_o,
  v_o,
  ready_i
);

  input [540:0] data_i;
  output [135:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input ready_i;
  output ready_o;
  output v_o;
  wire [135:0] data_o;
  wire ready_o,v_o,N0,N1,N2,N3,state_n,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24,N25;
  wire [1:0] count_n;
  reg [1:0] count_r;
  reg state_r;

  bsg_mux_width_p136_els_p4
  mux
  (
    .data_i({ 1'b0, 1'b0, 1'b0, data_i }),
    .sel_i(count_r),
    .data_o(data_o)
  );

  assign N10 = count_r == data_i[3:2];
  assign N12 = count_r == data_i[3:2];
  assign { N9, N8 } = count_r + 1'b1;
  assign N14 = ~N13;
  assign count_n = (N0)? { 1'b0, 1'b0 } :
                   (N1)? { N9, N8 } : 1'b0;
  assign N0 = N4;
  assign N1 = v_o;
  assign state_n = (N0)? 1'b1 :
                   (N1)? N14 : 1'b0;
  assign ready_o = (N0)? 1'b0 :
                   (N1)? N11 : 1'b0;
  assign N16 = (N2)? 1'b0 :
               (N3)? state_n : 1'b0;
  assign N2 = reset_i;
  assign N3 = N15;
  assign { N18, N17 } = (N2)? { 1'b0, 1'b0 } :
                        (N3)? count_n : 1'b0;
  assign N4 = ~state_r;
  assign v_o = state_r;
  assign N5 = ~v_i;
  assign N6 = v_o;
  assign N7 = ~ready_i;
  assign N11 = ready_i & N10;
  assign N13 = ready_i & N12;
  assign N15 = ~reset_i;
  assign N19 = N4 & N15;
  assign N20 = N5 & N19;
  assign N21 = v_o & N15;
  assign N22 = N7 & N21;
  assign N23 = N20 | N22;
  assign N24 = ~N23;
  assign N25 = ~N20;

  always @(posedge clk_i) begin
    if(N24) begin
      { count_r[1:0] } <= { N18, N17 };
    end
    if(N25) begin
      state_r <= N16;
    end
  end


endmodule



module bsg_wormhole_router_adapter_out_max_num_flit_p4_max_payload_width_p537_x_cord_width_p1_y_cord_width_p1
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  ready_o,
  data_o,
  v_o,
  ready_i
);

  input [135:0] data_i;
  output [540:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input ready_i;
  output ready_o;
  output v_o;
  wire ready_o,v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,we,clear,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,
  N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,
  N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,
  N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,
  N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,
  N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,
  N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,
  N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,
  N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211,N212,N213,N214,N215,N216;
  wire [1:0] state_n,count_n;
  reg [540:0] data_o;
  reg [1:0] state_r,count_r;
  assign N16 = N14 & N15;
  assign N17 = state_r[1] | N15;
  assign N19 = N14 | state_r[0];
  assign N21 = state_r[1] & state_r[0];
  assign N29 = data_o[3:2] == count_r;
  assign N215 = data_i[2] | data_i[3];
  assign N216 = ~N215;
  assign { N25, N24 } = count_r + 1'b1;
  assign { N28, N27 } = count_r + 1'b1;
  assign N38 = count_r[0] & count_r[1];
  assign N37 = N0 & count_r[1];
  assign N0 = ~count_r[0];
  assign N36 = count_r[0] & N1;
  assign N1 = ~count_r[1];
  assign N35 = N2 & N3;
  assign N2 = ~count_r[0];
  assign N3 = ~count_r[1];
  assign N30 = ~N29;
  assign ready_o = (N4)? 1'b1 :
                   (N5)? 1'b1 :
                   (N6)? 1'b0 :
                   (N7)? 1'b0 : 1'b0;
  assign N4 = N16;
  assign N5 = N18;
  assign N6 = N20;
  assign N7 = N21;
  assign state_n = (N4)? { N216, N215 } :
                   (N5)? { N29, N30 } :
                   (N6)? { 1'b0, 1'b0 } :
                   (N7)? { 1'b0, 1'b0 } : 1'b0;
  assign we = (N4)? v_i :
              (N5)? v_i :
              (N6)? ready_i :
              (N7)? 1'b0 : 1'b0;
  assign count_n = (N4)? { N25, N24 } :
                   (N5)? { N28, N27 } :
                   (N6)? { 1'b0, 1'b0 } : 1'b0;
  assign v_o = (N4)? 1'b0 :
               (N5)? 1'b0 :
               (N6)? 1'b1 :
               (N7)? 1'b0 : 1'b0;
  assign clear = (N4)? 1'b0 :
                 (N5)? 1'b0 :
                 (N6)? ready_i :
                 (N7)? 1'b0 : 1'b0;
  assign { N182, N181, N180, N179, N178, N177, N41, N39 } = (N8)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } :
                                                            (N9)? { N38, N38, N37, N37, N36, N36, N35, N35 } : 1'b0;
  assign N8 = clear;
  assign N9 = N34;
  assign { N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N40 } = (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   (N9)? data_i : 1'b0;
  assign { N190, N189, N188, N187, N186, N185, N184, N183 } = (N10)? { N182, N181, N180, N179, N178, N177, N41, N39 } :
                                                              (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = we;
  assign N11 = N33;
  assign { N192, N191 } = (N12)? { 1'b0, 1'b0 } :
                          (N13)? state_n : 1'b0;
  assign N12 = reset_i;
  assign N13 = N32;
  assign { N194, N193 } = (N12)? { 1'b0, 1'b0 } :
                          (N13)? count_n : 1'b0;
  assign { N202, N201, N200, N199, N198, N197, N196, N195 } = (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                              (N13)? { N190, N189, N188, N187, N186, N185, N184, N183 } : 1'b0;
  assign N14 = ~state_r[1];
  assign N15 = ~state_r[0];
  assign N18 = ~N17;
  assign N20 = ~N19;
  assign N22 = N16;
  assign N23 = ~v_i;
  assign N26 = N18;
  assign N31 = ~ready_i;
  assign N32 = ~reset_i;
  assign N33 = ~we;
  assign N34 = ~clear;
  assign N203 = N16 & N32;
  assign N204 = N23 & N203;
  assign N205 = N18 & N32;
  assign N206 = N23 & N205;
  assign N207 = N204 | N206;
  assign N208 = N20 & N32;
  assign N209 = N31 & N208;
  assign N210 = N207 | N209;
  assign N211 = ~N210;
  assign N212 = N21 & N32;
  assign N213 = N210 | N212;
  assign N214 = ~N213;

  always @(posedge clk_i) begin
    if(N201) begin
      { data_o[540:442], data_o[408:408] } <= { N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N40 };
    end
    if(N202) begin
      { data_o[441:409] } <= { N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42 };
    end
    if(N199) begin
      { data_o[407:309], data_o[272:272] } <= { N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N40 };
    end
    if(N200) begin
      { data_o[308:273] } <= { N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42 };
    end
    if(N197) begin
      { data_o[271:173], data_o[136:136] } <= { N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N40 };
    end
    if(N198) begin
      { data_o[172:137] } <= { N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42 };
    end
    if(N195) begin
      { data_o[135:37], data_o[0:0] } <= { N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N40 };
    end
    if(N196) begin
      { data_o[36:1] } <= { N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42 };
    end
    if(N211) begin
      { state_r[1:0] } <= { N192, N191 };
    end
    if(N214) begin
      { count_r[1:0] } <= { N194, N193 };
    end
  end


endmodule



module bp_me_network_channel_data_resp_num_lce_p2_num_cce_p1_paddr_width_p22_block_size_in_bits_p512_max_num_flit_p4
(
  clk_i,
  reset_i,
  lce_data_resp_i,
  lce_data_resp_v_i,
  lce_data_resp_ready_o,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i
);

  input [1073:0] lce_data_resp_i;
  input [1:0] lce_data_resp_v_i;
  output [1:0] lce_data_resp_ready_o;
  output [536:0] lce_data_resp_o;
  output [0:0] lce_data_resp_v_o;
  input [0:0] lce_data_resp_ready_i;
  input clk_i;
  input reset_i;
  wire [1:0] lce_data_resp_ready_o;
  wire [536:0] lce_data_resp_o;
  wire [0:0] lce_data_resp_v_o;
  wire valid_li_1__4_,valid_li_1__3_,valid_li_1__2_,valid_li_1__0_,valid_li_0__4_,
  valid_li_0__3_,valid_li_0__1_,valid_li_0__0_,data_li_1__0__135_,data_li_1__0__134_,
  data_li_1__0__133_,data_li_1__0__132_,data_li_1__0__131_,data_li_1__0__130_,
  data_li_1__0__129_,data_li_1__0__128_,data_li_1__0__127_,data_li_1__0__126_,
  data_li_1__0__125_,data_li_1__0__124_,data_li_1__0__123_,data_li_1__0__122_,
  data_li_1__0__121_,data_li_1__0__120_,data_li_1__0__119_,data_li_1__0__118_,
  data_li_1__0__117_,data_li_1__0__116_,data_li_1__0__115_,data_li_1__0__114_,data_li_1__0__113_,
  data_li_1__0__112_,data_li_1__0__111_,data_li_1__0__110_,data_li_1__0__109_,
  data_li_1__0__108_,data_li_1__0__107_,data_li_1__0__106_,data_li_1__0__105_,
  data_li_1__0__104_,data_li_1__0__103_,data_li_1__0__102_,data_li_1__0__101_,
  data_li_1__0__100_,data_li_1__0__99_,data_li_1__0__98_,data_li_1__0__97_,data_li_1__0__96_,
  data_li_1__0__95_,data_li_1__0__94_,data_li_1__0__93_,data_li_1__0__92_,
  data_li_1__0__91_,data_li_1__0__90_,data_li_1__0__89_,data_li_1__0__88_,data_li_1__0__87_,
  data_li_1__0__86_,data_li_1__0__85_,data_li_1__0__84_,data_li_1__0__83_,
  data_li_1__0__82_,data_li_1__0__81_,data_li_1__0__80_,data_li_1__0__79_,data_li_1__0__78_,
  data_li_1__0__77_,data_li_1__0__76_,data_li_1__0__75_,data_li_1__0__74_,
  data_li_1__0__73_,data_li_1__0__72_,data_li_1__0__71_,data_li_1__0__70_,
  data_li_1__0__69_,data_li_1__0__68_,data_li_1__0__67_,data_li_1__0__66_,data_li_1__0__65_,
  data_li_1__0__64_,data_li_1__0__63_,data_li_1__0__62_,data_li_1__0__61_,
  data_li_1__0__60_,data_li_1__0__59_,data_li_1__0__58_,data_li_1__0__57_,data_li_1__0__56_,
  data_li_1__0__55_,data_li_1__0__54_,data_li_1__0__53_,data_li_1__0__52_,
  data_li_1__0__51_,data_li_1__0__50_,data_li_1__0__49_,data_li_1__0__48_,data_li_1__0__47_,
  data_li_1__0__46_,data_li_1__0__45_,data_li_1__0__44_,data_li_1__0__43_,
  data_li_1__0__42_,data_li_1__0__41_,data_li_1__0__40_,data_li_1__0__39_,data_li_1__0__38_,
  data_li_1__0__37_,data_li_1__0__36_,data_li_1__0__35_,data_li_1__0__34_,
  data_li_1__0__33_,data_li_1__0__32_,data_li_1__0__31_,data_li_1__0__30_,
  data_li_1__0__29_,data_li_1__0__28_,data_li_1__0__27_,data_li_1__0__26_,data_li_1__0__25_,
  data_li_1__0__24_,data_li_1__0__23_,data_li_1__0__22_,data_li_1__0__21_,
  data_li_1__0__20_,data_li_1__0__19_,data_li_1__0__18_,data_li_1__0__17_,data_li_1__0__16_,
  data_li_1__0__15_,data_li_1__0__14_,data_li_1__0__13_,data_li_1__0__12_,
  data_li_1__0__11_,data_li_1__0__10_,data_li_1__0__9_,data_li_1__0__8_,data_li_1__0__7_,
  data_li_1__0__6_,data_li_1__0__5_,data_li_1__0__4_,data_li_1__0__3_,data_li_1__0__2_,
  data_li_1__0__1_,data_li_1__0__0_,data_li_0__4__135_,data_li_0__4__134_,
  data_li_0__4__133_,data_li_0__4__132_,data_li_0__4__131_,data_li_0__4__130_,
  data_li_0__4__129_,data_li_0__4__128_,data_li_0__4__127_,data_li_0__4__126_,
  data_li_0__4__125_,data_li_0__4__124_,data_li_0__4__123_,data_li_0__4__122_,data_li_0__4__121_,
  data_li_0__4__120_,data_li_0__4__119_,data_li_0__4__118_,data_li_0__4__117_,
  data_li_0__4__116_,data_li_0__4__115_,data_li_0__4__114_,data_li_0__4__113_,
  data_li_0__4__112_,data_li_0__4__111_,data_li_0__4__110_,data_li_0__4__109_,
  data_li_0__4__108_,data_li_0__4__107_,data_li_0__4__106_,data_li_0__4__105_,
  data_li_0__4__104_,data_li_0__4__103_,data_li_0__4__102_,data_li_0__4__101_,data_li_0__4__100_,
  data_li_0__4__99_,data_li_0__4__98_,data_li_0__4__97_,data_li_0__4__96_,
  data_li_0__4__95_,data_li_0__4__94_,data_li_0__4__93_,data_li_0__4__92_,data_li_0__4__91_,
  data_li_0__4__90_,data_li_0__4__89_,data_li_0__4__88_,data_li_0__4__87_,
  data_li_0__4__86_,data_li_0__4__85_,data_li_0__4__84_,data_li_0__4__83_,
  data_li_0__4__82_,data_li_0__4__81_,data_li_0__4__80_,data_li_0__4__79_,data_li_0__4__78_,
  data_li_0__4__77_,data_li_0__4__76_,data_li_0__4__75_,data_li_0__4__74_,
  data_li_0__4__73_,data_li_0__4__72_,data_li_0__4__71_,data_li_0__4__70_,data_li_0__4__69_,
  data_li_0__4__68_,data_li_0__4__67_,data_li_0__4__66_,data_li_0__4__65_,
  data_li_0__4__64_,data_li_0__4__63_,data_li_0__4__62_,data_li_0__4__61_,data_li_0__4__60_,
  data_li_0__4__59_,data_li_0__4__58_,data_li_0__4__57_,data_li_0__4__56_,
  data_li_0__4__55_,data_li_0__4__54_,data_li_0__4__53_,data_li_0__4__52_,data_li_0__4__51_,
  data_li_0__4__50_,data_li_0__4__49_,data_li_0__4__48_,data_li_0__4__47_,
  data_li_0__4__46_,data_li_0__4__45_,data_li_0__4__44_,data_li_0__4__43_,
  data_li_0__4__42_,data_li_0__4__41_,data_li_0__4__40_,data_li_0__4__39_,data_li_0__4__38_,
  data_li_0__4__37_,data_li_0__4__36_,data_li_0__4__35_,data_li_0__4__34_,
  data_li_0__4__33_,data_li_0__4__32_,data_li_0__4__31_,data_li_0__4__30_,data_li_0__4__29_,
  data_li_0__4__28_,data_li_0__4__27_,data_li_0__4__26_,data_li_0__4__25_,
  data_li_0__4__24_,data_li_0__4__23_,data_li_0__4__22_,data_li_0__4__21_,data_li_0__4__20_,
  data_li_0__4__19_,data_li_0__4__18_,data_li_0__4__17_,data_li_0__4__16_,
  data_li_0__4__15_,data_li_0__4__14_,data_li_0__4__13_,data_li_0__4__12_,data_li_0__4__11_,
  data_li_0__4__10_,data_li_0__4__9_,data_li_0__4__8_,data_li_0__4__7_,
  data_li_0__4__6_,data_li_0__4__5_,data_li_0__4__4_,data_li_0__4__3_,data_li_0__4__2_,
  data_li_0__4__1_,data_li_0__4__0_,data_li_0__3__135_,data_li_0__3__134_,
  data_li_0__3__133_,data_li_0__3__132_,data_li_0__3__131_,data_li_0__3__130_,
  data_li_0__3__129_,data_li_0__3__128_,data_li_0__3__127_,data_li_0__3__126_,data_li_0__3__125_,
  data_li_0__3__124_,data_li_0__3__123_,data_li_0__3__122_,data_li_0__3__121_,
  data_li_0__3__120_,data_li_0__3__119_,data_li_0__3__118_,data_li_0__3__117_,
  data_li_0__3__116_,data_li_0__3__115_,data_li_0__3__114_,data_li_0__3__113_,
  data_li_0__3__112_,data_li_0__3__111_,data_li_0__3__110_,data_li_0__3__109_,data_li_0__3__108_,
  data_li_0__3__107_,data_li_0__3__106_,data_li_0__3__105_,data_li_0__3__104_,
  data_li_0__3__103_,data_li_0__3__102_,data_li_0__3__101_,data_li_0__3__100_,
  data_li_0__3__99_,data_li_0__3__98_,data_li_0__3__97_,data_li_0__3__96_,
  data_li_0__3__95_,data_li_0__3__94_,data_li_0__3__93_,data_li_0__3__92_,data_li_0__3__91_,
  data_li_0__3__90_,data_li_0__3__89_,data_li_0__3__88_,data_li_0__3__87_,
  data_li_0__3__86_,data_li_0__3__85_,data_li_0__3__84_,data_li_0__3__83_,data_li_0__3__82_,
  data_li_0__3__81_,data_li_0__3__80_,data_li_0__3__79_,data_li_0__3__78_,
  data_li_0__3__77_,data_li_0__3__76_,data_li_0__3__75_,data_li_0__3__74_,data_li_0__3__73_,
  data_li_0__3__72_,data_li_0__3__71_,data_li_0__3__70_,data_li_0__3__69_,
  data_li_0__3__68_,data_li_0__3__67_,data_li_0__3__66_,data_li_0__3__65_,data_li_0__3__64_,
  data_li_0__3__63_,data_li_0__3__62_,data_li_0__3__61_,data_li_0__3__60_,
  data_li_0__3__59_,data_li_0__3__58_,data_li_0__3__57_,data_li_0__3__56_,
  data_li_0__3__55_,data_li_0__3__54_,data_li_0__3__53_,data_li_0__3__52_,data_li_0__3__51_,
  data_li_0__3__50_,data_li_0__3__49_,data_li_0__3__48_,data_li_0__3__47_,
  data_li_0__3__46_,data_li_0__3__45_,data_li_0__3__44_,data_li_0__3__43_,data_li_0__3__42_,
  data_li_0__3__41_,data_li_0__3__40_,data_li_0__3__39_,data_li_0__3__38_,
  data_li_0__3__37_,data_li_0__3__36_,data_li_0__3__35_,data_li_0__3__34_,data_li_0__3__33_,
  data_li_0__3__32_,data_li_0__3__31_,data_li_0__3__30_,data_li_0__3__29_,
  data_li_0__3__28_,data_li_0__3__27_,data_li_0__3__26_,data_li_0__3__25_,data_li_0__3__24_,
  data_li_0__3__23_,data_li_0__3__22_,data_li_0__3__21_,data_li_0__3__20_,
  data_li_0__3__19_,data_li_0__3__18_,data_li_0__3__17_,data_li_0__3__16_,
  data_li_0__3__15_,data_li_0__3__14_,data_li_0__3__13_,data_li_0__3__12_,data_li_0__3__11_,
  data_li_0__3__10_,data_li_0__3__9_,data_li_0__3__8_,data_li_0__3__7_,data_li_0__3__6_,
  data_li_0__3__5_,data_li_0__3__4_,data_li_0__3__3_,data_li_0__3__2_,
  data_li_0__3__1_,data_li_0__3__0_,data_li_0__1__135_,data_li_0__1__134_,data_li_0__1__133_,
  data_li_0__1__132_,data_li_0__1__131_,data_li_0__1__130_,data_li_0__1__129_,
  data_li_0__1__128_,data_li_0__1__127_,data_li_0__1__126_,data_li_0__1__125_,
  data_li_0__1__124_,data_li_0__1__123_,data_li_0__1__122_,data_li_0__1__121_,
  data_li_0__1__120_,data_li_0__1__119_,data_li_0__1__118_,data_li_0__1__117_,
  data_li_0__1__116_,data_li_0__1__115_,data_li_0__1__114_,data_li_0__1__113_,data_li_0__1__112_,
  data_li_0__1__111_,data_li_0__1__110_,data_li_0__1__109_,data_li_0__1__108_,
  data_li_0__1__107_,data_li_0__1__106_,data_li_0__1__105_,data_li_0__1__104_,
  data_li_0__1__103_,data_li_0__1__102_,data_li_0__1__101_,data_li_0__1__100_,
  data_li_0__1__99_,data_li_0__1__98_,data_li_0__1__97_,data_li_0__1__96_,data_li_0__1__95_,
  data_li_0__1__94_,data_li_0__1__93_,data_li_0__1__92_,data_li_0__1__91_,
  data_li_0__1__90_,data_li_0__1__89_,data_li_0__1__88_,data_li_0__1__87_,data_li_0__1__86_,
  data_li_0__1__85_,data_li_0__1__84_,data_li_0__1__83_,data_li_0__1__82_,
  data_li_0__1__81_,data_li_0__1__80_,data_li_0__1__79_,data_li_0__1__78_,data_li_0__1__77_,
  data_li_0__1__76_,data_li_0__1__75_,data_li_0__1__74_,data_li_0__1__73_,
  data_li_0__1__72_,data_li_0__1__71_,data_li_0__1__70_,data_li_0__1__69_,
  data_li_0__1__68_,data_li_0__1__67_,data_li_0__1__66_,data_li_0__1__65_,data_li_0__1__64_,
  data_li_0__1__63_,data_li_0__1__62_,data_li_0__1__61_,data_li_0__1__60_,
  data_li_0__1__59_,data_li_0__1__58_,data_li_0__1__57_,data_li_0__1__56_,data_li_0__1__55_,
  data_li_0__1__54_,data_li_0__1__53_,data_li_0__1__52_,data_li_0__1__51_,
  data_li_0__1__50_,data_li_0__1__49_,data_li_0__1__48_,data_li_0__1__47_,data_li_0__1__46_,
  data_li_0__1__45_,data_li_0__1__44_,data_li_0__1__43_,data_li_0__1__42_,
  data_li_0__1__41_,data_li_0__1__40_,data_li_0__1__39_,data_li_0__1__38_,data_li_0__1__37_,
  data_li_0__1__36_,data_li_0__1__35_,data_li_0__1__34_,data_li_0__1__33_,
  data_li_0__1__32_,data_li_0__1__31_,data_li_0__1__30_,data_li_0__1__29_,
  data_li_0__1__28_,data_li_0__1__27_,data_li_0__1__26_,data_li_0__1__25_,data_li_0__1__24_,
  data_li_0__1__23_,data_li_0__1__22_,data_li_0__1__21_,data_li_0__1__20_,
  data_li_0__1__19_,data_li_0__1__18_,data_li_0__1__17_,data_li_0__1__16_,data_li_0__1__15_,
  data_li_0__1__14_,data_li_0__1__13_,data_li_0__1__12_,data_li_0__1__11_,
  data_li_0__1__10_,data_li_0__1__9_,data_li_0__1__8_,data_li_0__1__7_,data_li_0__1__6_,
  data_li_0__1__5_,data_li_0__1__4_,data_li_0__1__3_,data_li_0__1__2_,data_li_0__1__1_,
  data_li_0__1__0_,data_li_0__0__135_,data_li_0__0__134_,data_li_0__0__133_,
  data_li_0__0__132_,data_li_0__0__131_,data_li_0__0__130_,data_li_0__0__129_,
  data_li_0__0__128_,data_li_0__0__127_,data_li_0__0__126_,data_li_0__0__125_,
  data_li_0__0__124_,data_li_0__0__123_,data_li_0__0__122_,data_li_0__0__121_,data_li_0__0__120_,
  data_li_0__0__119_,data_li_0__0__118_,data_li_0__0__117_,data_li_0__0__116_,
  data_li_0__0__115_,data_li_0__0__114_,data_li_0__0__113_,data_li_0__0__112_,
  data_li_0__0__111_,data_li_0__0__110_,data_li_0__0__109_,data_li_0__0__108_,
  data_li_0__0__107_,data_li_0__0__106_,data_li_0__0__105_,data_li_0__0__104_,
  data_li_0__0__103_,data_li_0__0__102_,data_li_0__0__101_,data_li_0__0__100_,data_li_0__0__99_,
  data_li_0__0__98_,data_li_0__0__97_,data_li_0__0__96_,data_li_0__0__95_,
  data_li_0__0__94_,data_li_0__0__93_,data_li_0__0__92_,data_li_0__0__91_,data_li_0__0__90_,
  data_li_0__0__89_,data_li_0__0__88_,data_li_0__0__87_,data_li_0__0__86_,
  data_li_0__0__85_,data_li_0__0__84_,data_li_0__0__83_,data_li_0__0__82_,
  data_li_0__0__81_,data_li_0__0__80_,data_li_0__0__79_,data_li_0__0__78_,data_li_0__0__77_,
  data_li_0__0__76_,data_li_0__0__75_,data_li_0__0__74_,data_li_0__0__73_,
  data_li_0__0__72_,data_li_0__0__71_,data_li_0__0__70_,data_li_0__0__69_,data_li_0__0__68_,
  data_li_0__0__67_,data_li_0__0__66_,data_li_0__0__65_,data_li_0__0__64_,
  data_li_0__0__63_,data_li_0__0__62_,data_li_0__0__61_,data_li_0__0__60_,data_li_0__0__59_,
  data_li_0__0__58_,data_li_0__0__57_,data_li_0__0__56_,data_li_0__0__55_,
  data_li_0__0__54_,data_li_0__0__53_,data_li_0__0__52_,data_li_0__0__51_,data_li_0__0__50_,
  data_li_0__0__49_,data_li_0__0__48_,data_li_0__0__47_,data_li_0__0__46_,
  data_li_0__0__45_,data_li_0__0__44_,data_li_0__0__43_,data_li_0__0__42_,
  data_li_0__0__41_,data_li_0__0__40_,data_li_0__0__39_,data_li_0__0__38_,data_li_0__0__37_,
  data_li_0__0__36_,data_li_0__0__35_,data_li_0__0__34_,data_li_0__0__33_,
  data_li_0__0__32_,data_li_0__0__31_,data_li_0__0__30_,data_li_0__0__29_,data_li_0__0__28_,
  data_li_0__0__27_,data_li_0__0__26_,data_li_0__0__25_,data_li_0__0__24_,
  data_li_0__0__23_,data_li_0__0__22_,data_li_0__0__21_,data_li_0__0__20_,data_li_0__0__19_,
  data_li_0__0__18_,data_li_0__0__17_,data_li_0__0__16_,data_li_0__0__15_,
  data_li_0__0__14_,data_li_0__0__13_,data_li_0__0__12_,data_li_0__0__11_,data_li_0__0__10_,
  data_li_0__0__9_,data_li_0__0__8_,data_li_0__0__7_,data_li_0__0__6_,
  data_li_0__0__5_,data_li_0__0__4_,data_li_0__0__3_,data_li_0__0__2_,data_li_0__0__1_,
  data_li_0__0__0_,ready_li_1__4_,ready_li_1__3_,ready_li_1__2_,ready_li_1__0_,
  ready_li_0__4_,ready_li_0__3_,ready_li_0__1_,ready_li_0__0_,data_li_1__4__135_,
  data_li_1__4__134_,data_li_1__4__133_,data_li_1__4__132_,data_li_1__4__131_,
  data_li_1__4__130_,data_li_1__4__129_,data_li_1__4__128_,data_li_1__4__127_,data_li_1__4__126_,
  data_li_1__4__125_,data_li_1__4__124_,data_li_1__4__123_,data_li_1__4__122_,
  data_li_1__4__121_,data_li_1__4__120_,data_li_1__4__119_,data_li_1__4__118_,
  data_li_1__4__117_,data_li_1__4__116_,data_li_1__4__115_,data_li_1__4__114_,
  data_li_1__4__113_,data_li_1__4__112_,data_li_1__4__111_,data_li_1__4__110_,
  data_li_1__4__109_,data_li_1__4__108_,data_li_1__4__107_,data_li_1__4__106_,data_li_1__4__105_,
  data_li_1__4__104_,data_li_1__4__103_,data_li_1__4__102_,data_li_1__4__101_,
  data_li_1__4__100_,data_li_1__4__99_,data_li_1__4__98_,data_li_1__4__97_,
  data_li_1__4__96_,data_li_1__4__95_,data_li_1__4__94_,data_li_1__4__93_,data_li_1__4__92_,
  data_li_1__4__91_,data_li_1__4__90_,data_li_1__4__89_,data_li_1__4__88_,
  data_li_1__4__87_,data_li_1__4__86_,data_li_1__4__85_,data_li_1__4__84_,data_li_1__4__83_,
  data_li_1__4__82_,data_li_1__4__81_,data_li_1__4__80_,data_li_1__4__79_,
  data_li_1__4__78_,data_li_1__4__77_,data_li_1__4__76_,data_li_1__4__75_,
  data_li_1__4__74_,data_li_1__4__73_,data_li_1__4__72_,data_li_1__4__71_,data_li_1__4__70_,
  data_li_1__4__69_,data_li_1__4__68_,data_li_1__4__67_,data_li_1__4__66_,
  data_li_1__4__65_,data_li_1__4__64_,data_li_1__4__63_,data_li_1__4__62_,data_li_1__4__61_,
  data_li_1__4__60_,data_li_1__4__59_,data_li_1__4__58_,data_li_1__4__57_,
  data_li_1__4__56_,data_li_1__4__55_,data_li_1__4__54_,data_li_1__4__53_,data_li_1__4__52_,
  data_li_1__4__51_,data_li_1__4__50_,data_li_1__4__49_,data_li_1__4__48_,
  data_li_1__4__47_,data_li_1__4__46_,data_li_1__4__45_,data_li_1__4__44_,data_li_1__4__43_,
  data_li_1__4__42_,data_li_1__4__41_,data_li_1__4__40_,data_li_1__4__39_,
  data_li_1__4__38_,data_li_1__4__37_,data_li_1__4__36_,data_li_1__4__35_,
  data_li_1__4__34_,data_li_1__4__33_,data_li_1__4__32_,data_li_1__4__31_,data_li_1__4__30_,
  data_li_1__4__29_,data_li_1__4__28_,data_li_1__4__27_,data_li_1__4__26_,
  data_li_1__4__25_,data_li_1__4__24_,data_li_1__4__23_,data_li_1__4__22_,data_li_1__4__21_,
  data_li_1__4__20_,data_li_1__4__19_,data_li_1__4__18_,data_li_1__4__17_,
  data_li_1__4__16_,data_li_1__4__15_,data_li_1__4__14_,data_li_1__4__13_,data_li_1__4__12_,
  data_li_1__4__11_,data_li_1__4__10_,data_li_1__4__9_,data_li_1__4__8_,
  data_li_1__4__7_,data_li_1__4__6_,data_li_1__4__5_,data_li_1__4__4_,data_li_1__4__3_,
  data_li_1__4__2_,data_li_1__4__1_,data_li_1__4__0_,data_li_1__3__135_,
  data_li_1__3__134_,data_li_1__3__133_,data_li_1__3__132_,data_li_1__3__131_,data_li_1__3__130_,
  data_li_1__3__129_,data_li_1__3__128_,data_li_1__3__127_,data_li_1__3__126_,
  data_li_1__3__125_,data_li_1__3__124_,data_li_1__3__123_,data_li_1__3__122_,
  data_li_1__3__121_,data_li_1__3__120_,data_li_1__3__119_,data_li_1__3__118_,
  data_li_1__3__117_,data_li_1__3__116_,data_li_1__3__115_,data_li_1__3__114_,
  data_li_1__3__113_,data_li_1__3__112_,data_li_1__3__111_,data_li_1__3__110_,data_li_1__3__109_,
  data_li_1__3__108_,data_li_1__3__107_,data_li_1__3__106_,data_li_1__3__105_,
  data_li_1__3__104_,data_li_1__3__103_,data_li_1__3__102_,data_li_1__3__101_,
  data_li_1__3__100_,data_li_1__3__99_,data_li_1__3__98_,data_li_1__3__97_,data_li_1__3__96_,
  data_li_1__3__95_,data_li_1__3__94_,data_li_1__3__93_,data_li_1__3__92_,
  data_li_1__3__91_,data_li_1__3__90_,data_li_1__3__89_,data_li_1__3__88_,
  data_li_1__3__87_,data_li_1__3__86_,data_li_1__3__85_,data_li_1__3__84_,data_li_1__3__83_,
  data_li_1__3__82_,data_li_1__3__81_,data_li_1__3__80_,data_li_1__3__79_,
  data_li_1__3__78_,data_li_1__3__77_,data_li_1__3__76_,data_li_1__3__75_,data_li_1__3__74_,
  data_li_1__3__73_,data_li_1__3__72_,data_li_1__3__71_,data_li_1__3__70_,
  data_li_1__3__69_,data_li_1__3__68_,data_li_1__3__67_,data_li_1__3__66_,data_li_1__3__65_,
  data_li_1__3__64_,data_li_1__3__63_,data_li_1__3__62_,data_li_1__3__61_,
  data_li_1__3__60_,data_li_1__3__59_,data_li_1__3__58_,data_li_1__3__57_,data_li_1__3__56_,
  data_li_1__3__55_,data_li_1__3__54_,data_li_1__3__53_,data_li_1__3__52_,
  data_li_1__3__51_,data_li_1__3__50_,data_li_1__3__49_,data_li_1__3__48_,
  data_li_1__3__47_,data_li_1__3__46_,data_li_1__3__45_,data_li_1__3__44_,data_li_1__3__43_,
  data_li_1__3__42_,data_li_1__3__41_,data_li_1__3__40_,data_li_1__3__39_,
  data_li_1__3__38_,data_li_1__3__37_,data_li_1__3__36_,data_li_1__3__35_,data_li_1__3__34_,
  data_li_1__3__33_,data_li_1__3__32_,data_li_1__3__31_,data_li_1__3__30_,
  data_li_1__3__29_,data_li_1__3__28_,data_li_1__3__27_,data_li_1__3__26_,data_li_1__3__25_,
  data_li_1__3__24_,data_li_1__3__23_,data_li_1__3__22_,data_li_1__3__21_,
  data_li_1__3__20_,data_li_1__3__19_,data_li_1__3__18_,data_li_1__3__17_,data_li_1__3__16_,
  data_li_1__3__15_,data_li_1__3__14_,data_li_1__3__13_,data_li_1__3__12_,
  data_li_1__3__11_,data_li_1__3__10_,data_li_1__3__9_,data_li_1__3__8_,data_li_1__3__7_,
  data_li_1__3__6_,data_li_1__3__5_,data_li_1__3__4_,data_li_1__3__3_,
  data_li_1__3__2_,data_li_1__3__1_,data_li_1__3__0_,data_li_1__2__135_,data_li_1__2__134_,
  data_li_1__2__133_,data_li_1__2__132_,data_li_1__2__131_,data_li_1__2__130_,
  data_li_1__2__129_,data_li_1__2__128_,data_li_1__2__127_,data_li_1__2__126_,
  data_li_1__2__125_,data_li_1__2__124_,data_li_1__2__123_,data_li_1__2__122_,
  data_li_1__2__121_,data_li_1__2__120_,data_li_1__2__119_,data_li_1__2__118_,data_li_1__2__117_,
  data_li_1__2__116_,data_li_1__2__115_,data_li_1__2__114_,data_li_1__2__113_,
  data_li_1__2__112_,data_li_1__2__111_,data_li_1__2__110_,data_li_1__2__109_,
  data_li_1__2__108_,data_li_1__2__107_,data_li_1__2__106_,data_li_1__2__105_,
  data_li_1__2__104_,data_li_1__2__103_,data_li_1__2__102_,data_li_1__2__101_,
  data_li_1__2__100_,data_li_1__2__99_,data_li_1__2__98_,data_li_1__2__97_,data_li_1__2__96_,
  data_li_1__2__95_,data_li_1__2__94_,data_li_1__2__93_,data_li_1__2__92_,
  data_li_1__2__91_,data_li_1__2__90_,data_li_1__2__89_,data_li_1__2__88_,data_li_1__2__87_,
  data_li_1__2__86_,data_li_1__2__85_,data_li_1__2__84_,data_li_1__2__83_,
  data_li_1__2__82_,data_li_1__2__81_,data_li_1__2__80_,data_li_1__2__79_,data_li_1__2__78_,
  data_li_1__2__77_,data_li_1__2__76_,data_li_1__2__75_,data_li_1__2__74_,
  data_li_1__2__73_,data_li_1__2__72_,data_li_1__2__71_,data_li_1__2__70_,data_li_1__2__69_,
  data_li_1__2__68_,data_li_1__2__67_,data_li_1__2__66_,data_li_1__2__65_,
  data_li_1__2__64_,data_li_1__2__63_,data_li_1__2__62_,data_li_1__2__61_,
  data_li_1__2__60_,data_li_1__2__59_,data_li_1__2__58_,data_li_1__2__57_,data_li_1__2__56_,
  data_li_1__2__55_,data_li_1__2__54_,data_li_1__2__53_,data_li_1__2__52_,
  data_li_1__2__51_,data_li_1__2__50_,data_li_1__2__49_,data_li_1__2__48_,data_li_1__2__47_,
  data_li_1__2__46_,data_li_1__2__45_,data_li_1__2__44_,data_li_1__2__43_,
  data_li_1__2__42_,data_li_1__2__41_,data_li_1__2__40_,data_li_1__2__39_,data_li_1__2__38_,
  data_li_1__2__37_,data_li_1__2__36_,data_li_1__2__35_,data_li_1__2__34_,
  data_li_1__2__33_,data_li_1__2__32_,data_li_1__2__31_,data_li_1__2__30_,data_li_1__2__29_,
  data_li_1__2__28_,data_li_1__2__27_,data_li_1__2__26_,data_li_1__2__25_,
  data_li_1__2__24_,data_li_1__2__23_,data_li_1__2__22_,data_li_1__2__21_,
  data_li_1__2__20_,data_li_1__2__19_,data_li_1__2__18_,data_li_1__2__17_,data_li_1__2__16_,
  data_li_1__2__15_,data_li_1__2__14_,data_li_1__2__13_,data_li_1__2__12_,
  data_li_1__2__11_,data_li_1__2__10_,data_li_1__2__9_,data_li_1__2__8_,data_li_1__2__7_,
  data_li_1__2__6_,data_li_1__2__5_,data_li_1__2__4_,data_li_1__2__3_,data_li_1__2__2_,
  data_li_1__2__1_,data_li_1__2__0_,cce_packet_0__3_,cce_packet_0__2_,
  cce_packet_0__1_,cce_packet_0__0_;
  wire [9:0] ready_lo,valid_lo;
  wire [1359:0] data_lo;
  wire [1081:0] lce_packet;

  bsg_wormhole_router_136_1_1_2_1_1_1_00000013_0000001a
  router_0__router
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .local_x_cord_i(1'b0),
    .local_y_cord_i(1'b0),
    .valid_i({ valid_li_0__4_, valid_li_0__3_, valid_lo[6:6], valid_li_0__1_, valid_li_0__0_ }),
    .data_i({ data_li_0__4__135_, data_li_0__4__134_, data_li_0__4__133_, data_li_0__4__132_, data_li_0__4__131_, data_li_0__4__130_, data_li_0__4__129_, data_li_0__4__128_, data_li_0__4__127_, data_li_0__4__126_, data_li_0__4__125_, data_li_0__4__124_, data_li_0__4__123_, data_li_0__4__122_, data_li_0__4__121_, data_li_0__4__120_, data_li_0__4__119_, data_li_0__4__118_, data_li_0__4__117_, data_li_0__4__116_, data_li_0__4__115_, data_li_0__4__114_, data_li_0__4__113_, data_li_0__4__112_, data_li_0__4__111_, data_li_0__4__110_, data_li_0__4__109_, data_li_0__4__108_, data_li_0__4__107_, data_li_0__4__106_, data_li_0__4__105_, data_li_0__4__104_, data_li_0__4__103_, data_li_0__4__102_, data_li_0__4__101_, data_li_0__4__100_, data_li_0__4__99_, data_li_0__4__98_, data_li_0__4__97_, data_li_0__4__96_, data_li_0__4__95_, data_li_0__4__94_, data_li_0__4__93_, data_li_0__4__92_, data_li_0__4__91_, data_li_0__4__90_, data_li_0__4__89_, data_li_0__4__88_, data_li_0__4__87_, data_li_0__4__86_, data_li_0__4__85_, data_li_0__4__84_, data_li_0__4__83_, data_li_0__4__82_, data_li_0__4__81_, data_li_0__4__80_, data_li_0__4__79_, data_li_0__4__78_, data_li_0__4__77_, data_li_0__4__76_, data_li_0__4__75_, data_li_0__4__74_, data_li_0__4__73_, data_li_0__4__72_, data_li_0__4__71_, data_li_0__4__70_, data_li_0__4__69_, data_li_0__4__68_, data_li_0__4__67_, data_li_0__4__66_, data_li_0__4__65_, data_li_0__4__64_, data_li_0__4__63_, data_li_0__4__62_, data_li_0__4__61_, data_li_0__4__60_, data_li_0__4__59_, data_li_0__4__58_, data_li_0__4__57_, data_li_0__4__56_, data_li_0__4__55_, data_li_0__4__54_, data_li_0__4__53_, data_li_0__4__52_, data_li_0__4__51_, data_li_0__4__50_, data_li_0__4__49_, data_li_0__4__48_, data_li_0__4__47_, data_li_0__4__46_, data_li_0__4__45_, data_li_0__4__44_, data_li_0__4__43_, data_li_0__4__42_, data_li_0__4__41_, data_li_0__4__40_, data_li_0__4__39_, data_li_0__4__38_, data_li_0__4__37_, data_li_0__4__36_, data_li_0__4__35_, data_li_0__4__34_, data_li_0__4__33_, data_li_0__4__32_, data_li_0__4__31_, data_li_0__4__30_, data_li_0__4__29_, data_li_0__4__28_, data_li_0__4__27_, data_li_0__4__26_, data_li_0__4__25_, data_li_0__4__24_, data_li_0__4__23_, data_li_0__4__22_, data_li_0__4__21_, data_li_0__4__20_, data_li_0__4__19_, data_li_0__4__18_, data_li_0__4__17_, data_li_0__4__16_, data_li_0__4__15_, data_li_0__4__14_, data_li_0__4__13_, data_li_0__4__12_, data_li_0__4__11_, data_li_0__4__10_, data_li_0__4__9_, data_li_0__4__8_, data_li_0__4__7_, data_li_0__4__6_, data_li_0__4__5_, data_li_0__4__4_, data_li_0__4__3_, data_li_0__4__2_, data_li_0__4__1_, data_li_0__4__0_, data_li_0__3__135_, data_li_0__3__134_, data_li_0__3__133_, data_li_0__3__132_, data_li_0__3__131_, data_li_0__3__130_, data_li_0__3__129_, data_li_0__3__128_, data_li_0__3__127_, data_li_0__3__126_, data_li_0__3__125_, data_li_0__3__124_, data_li_0__3__123_, data_li_0__3__122_, data_li_0__3__121_, data_li_0__3__120_, data_li_0__3__119_, data_li_0__3__118_, data_li_0__3__117_, data_li_0__3__116_, data_li_0__3__115_, data_li_0__3__114_, data_li_0__3__113_, data_li_0__3__112_, data_li_0__3__111_, data_li_0__3__110_, data_li_0__3__109_, data_li_0__3__108_, data_li_0__3__107_, data_li_0__3__106_, data_li_0__3__105_, data_li_0__3__104_, data_li_0__3__103_, data_li_0__3__102_, data_li_0__3__101_, data_li_0__3__100_, data_li_0__3__99_, data_li_0__3__98_, data_li_0__3__97_, data_li_0__3__96_, data_li_0__3__95_, data_li_0__3__94_, data_li_0__3__93_, data_li_0__3__92_, data_li_0__3__91_, data_li_0__3__90_, data_li_0__3__89_, data_li_0__3__88_, data_li_0__3__87_, data_li_0__3__86_, data_li_0__3__85_, data_li_0__3__84_, data_li_0__3__83_, data_li_0__3__82_, data_li_0__3__81_, data_li_0__3__80_, data_li_0__3__79_, data_li_0__3__78_, data_li_0__3__77_, data_li_0__3__76_, data_li_0__3__75_, data_li_0__3__74_, data_li_0__3__73_, data_li_0__3__72_, data_li_0__3__71_, data_li_0__3__70_, data_li_0__3__69_, data_li_0__3__68_, data_li_0__3__67_, data_li_0__3__66_, data_li_0__3__65_, data_li_0__3__64_, data_li_0__3__63_, data_li_0__3__62_, data_li_0__3__61_, data_li_0__3__60_, data_li_0__3__59_, data_li_0__3__58_, data_li_0__3__57_, data_li_0__3__56_, data_li_0__3__55_, data_li_0__3__54_, data_li_0__3__53_, data_li_0__3__52_, data_li_0__3__51_, data_li_0__3__50_, data_li_0__3__49_, data_li_0__3__48_, data_li_0__3__47_, data_li_0__3__46_, data_li_0__3__45_, data_li_0__3__44_, data_li_0__3__43_, data_li_0__3__42_, data_li_0__3__41_, data_li_0__3__40_, data_li_0__3__39_, data_li_0__3__38_, data_li_0__3__37_, data_li_0__3__36_, data_li_0__3__35_, data_li_0__3__34_, data_li_0__3__33_, data_li_0__3__32_, data_li_0__3__31_, data_li_0__3__30_, data_li_0__3__29_, data_li_0__3__28_, data_li_0__3__27_, data_li_0__3__26_, data_li_0__3__25_, data_li_0__3__24_, data_li_0__3__23_, data_li_0__3__22_, data_li_0__3__21_, data_li_0__3__20_, data_li_0__3__19_, data_li_0__3__18_, data_li_0__3__17_, data_li_0__3__16_, data_li_0__3__15_, data_li_0__3__14_, data_li_0__3__13_, data_li_0__3__12_, data_li_0__3__11_, data_li_0__3__10_, data_li_0__3__9_, data_li_0__3__8_, data_li_0__3__7_, data_li_0__3__6_, data_li_0__3__5_, data_li_0__3__4_, data_li_0__3__3_, data_li_0__3__2_, data_li_0__3__1_, data_li_0__3__0_, data_lo[951:816], data_li_0__1__135_, data_li_0__1__134_, data_li_0__1__133_, data_li_0__1__132_, data_li_0__1__131_, data_li_0__1__130_, data_li_0__1__129_, data_li_0__1__128_, data_li_0__1__127_, data_li_0__1__126_, data_li_0__1__125_, data_li_0__1__124_, data_li_0__1__123_, data_li_0__1__122_, data_li_0__1__121_, data_li_0__1__120_, data_li_0__1__119_, data_li_0__1__118_, data_li_0__1__117_, data_li_0__1__116_, data_li_0__1__115_, data_li_0__1__114_, data_li_0__1__113_, data_li_0__1__112_, data_li_0__1__111_, data_li_0__1__110_, data_li_0__1__109_, data_li_0__1__108_, data_li_0__1__107_, data_li_0__1__106_, data_li_0__1__105_, data_li_0__1__104_, data_li_0__1__103_, data_li_0__1__102_, data_li_0__1__101_, data_li_0__1__100_, data_li_0__1__99_, data_li_0__1__98_, data_li_0__1__97_, data_li_0__1__96_, data_li_0__1__95_, data_li_0__1__94_, data_li_0__1__93_, data_li_0__1__92_, data_li_0__1__91_, data_li_0__1__90_, data_li_0__1__89_, data_li_0__1__88_, data_li_0__1__87_, data_li_0__1__86_, data_li_0__1__85_, data_li_0__1__84_, data_li_0__1__83_, data_li_0__1__82_, data_li_0__1__81_, data_li_0__1__80_, data_li_0__1__79_, data_li_0__1__78_, data_li_0__1__77_, data_li_0__1__76_, data_li_0__1__75_, data_li_0__1__74_, data_li_0__1__73_, data_li_0__1__72_, data_li_0__1__71_, data_li_0__1__70_, data_li_0__1__69_, data_li_0__1__68_, data_li_0__1__67_, data_li_0__1__66_, data_li_0__1__65_, data_li_0__1__64_, data_li_0__1__63_, data_li_0__1__62_, data_li_0__1__61_, data_li_0__1__60_, data_li_0__1__59_, data_li_0__1__58_, data_li_0__1__57_, data_li_0__1__56_, data_li_0__1__55_, data_li_0__1__54_, data_li_0__1__53_, data_li_0__1__52_, data_li_0__1__51_, data_li_0__1__50_, data_li_0__1__49_, data_li_0__1__48_, data_li_0__1__47_, data_li_0__1__46_, data_li_0__1__45_, data_li_0__1__44_, data_li_0__1__43_, data_li_0__1__42_, data_li_0__1__41_, data_li_0__1__40_, data_li_0__1__39_, data_li_0__1__38_, data_li_0__1__37_, data_li_0__1__36_, data_li_0__1__35_, data_li_0__1__34_, data_li_0__1__33_, data_li_0__1__32_, data_li_0__1__31_, data_li_0__1__30_, data_li_0__1__29_, data_li_0__1__28_, data_li_0__1__27_, data_li_0__1__26_, data_li_0__1__25_, data_li_0__1__24_, data_li_0__1__23_, data_li_0__1__22_, data_li_0__1__21_, data_li_0__1__20_, data_li_0__1__19_, data_li_0__1__18_, data_li_0__1__17_, data_li_0__1__16_, data_li_0__1__15_, data_li_0__1__14_, data_li_0__1__13_, data_li_0__1__12_, data_li_0__1__11_, data_li_0__1__10_, data_li_0__1__9_, data_li_0__1__8_, data_li_0__1__7_, data_li_0__1__6_, data_li_0__1__5_, data_li_0__1__4_, data_li_0__1__3_, data_li_0__1__2_, data_li_0__1__1_, data_li_0__1__0_, data_li_0__0__135_, data_li_0__0__134_, data_li_0__0__133_, data_li_0__0__132_, data_li_0__0__131_, data_li_0__0__130_, data_li_0__0__129_, data_li_0__0__128_, data_li_0__0__127_, data_li_0__0__126_, data_li_0__0__125_, data_li_0__0__124_, data_li_0__0__123_, data_li_0__0__122_, data_li_0__0__121_, data_li_0__0__120_, data_li_0__0__119_, data_li_0__0__118_, data_li_0__0__117_, data_li_0__0__116_, data_li_0__0__115_, data_li_0__0__114_, data_li_0__0__113_, data_li_0__0__112_, data_li_0__0__111_, data_li_0__0__110_, data_li_0__0__109_, data_li_0__0__108_, data_li_0__0__107_, data_li_0__0__106_, data_li_0__0__105_, data_li_0__0__104_, data_li_0__0__103_, data_li_0__0__102_, data_li_0__0__101_, data_li_0__0__100_, data_li_0__0__99_, data_li_0__0__98_, data_li_0__0__97_, data_li_0__0__96_, data_li_0__0__95_, data_li_0__0__94_, data_li_0__0__93_, data_li_0__0__92_, data_li_0__0__91_, data_li_0__0__90_, data_li_0__0__89_, data_li_0__0__88_, data_li_0__0__87_, data_li_0__0__86_, data_li_0__0__85_, data_li_0__0__84_, data_li_0__0__83_, data_li_0__0__82_, data_li_0__0__81_, data_li_0__0__80_, data_li_0__0__79_, data_li_0__0__78_, data_li_0__0__77_, data_li_0__0__76_, data_li_0__0__75_, data_li_0__0__74_, data_li_0__0__73_, data_li_0__0__72_, data_li_0__0__71_, data_li_0__0__70_, data_li_0__0__69_, data_li_0__0__68_, data_li_0__0__67_, data_li_0__0__66_, data_li_0__0__65_, data_li_0__0__64_, data_li_0__0__63_, data_li_0__0__62_, data_li_0__0__61_, data_li_0__0__60_, data_li_0__0__59_, data_li_0__0__58_, data_li_0__0__57_, data_li_0__0__56_, data_li_0__0__55_, data_li_0__0__54_, data_li_0__0__53_, data_li_0__0__52_, data_li_0__0__51_, data_li_0__0__50_, data_li_0__0__49_, data_li_0__0__48_, data_li_0__0__47_, data_li_0__0__46_, data_li_0__0__45_, data_li_0__0__44_, data_li_0__0__43_, data_li_0__0__42_, data_li_0__0__41_, data_li_0__0__40_, data_li_0__0__39_, data_li_0__0__38_, data_li_0__0__37_, data_li_0__0__36_, data_li_0__0__35_, data_li_0__0__34_, data_li_0__0__33_, data_li_0__0__32_, data_li_0__0__31_, data_li_0__0__30_, data_li_0__0__29_, data_li_0__0__28_, data_li_0__0__27_, data_li_0__0__26_, data_li_0__0__25_, data_li_0__0__24_, data_li_0__0__23_, data_li_0__0__22_, data_li_0__0__21_, data_li_0__0__20_, data_li_0__0__19_, data_li_0__0__18_, data_li_0__0__17_, data_li_0__0__16_, data_li_0__0__15_, data_li_0__0__14_, data_li_0__0__13_, data_li_0__0__12_, data_li_0__0__11_, data_li_0__0__10_, data_li_0__0__9_, data_li_0__0__8_, data_li_0__0__7_, data_li_0__0__6_, data_li_0__0__5_, data_li_0__0__4_, data_li_0__0__3_, data_li_0__0__2_, data_li_0__0__1_, data_li_0__0__0_ }),
    .ready_o(ready_lo[4:0]),
    .valid_o(valid_lo[4:0]),
    .data_o(data_lo[679:0]),
    .ready_i({ ready_li_0__4_, ready_li_0__3_, ready_lo[6:6], ready_li_0__1_, ready_li_0__0_ })
  );


  bsg_wormhole_router_136_1_1_2_1_1_1_00000015_0000001c
  router_1__router
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .local_x_cord_i(1'b1),
    .local_y_cord_i(1'b0),
    .valid_i({ valid_li_1__4_, valid_li_1__3_, valid_li_1__2_, valid_lo[2:2], valid_li_1__0_ }),
    .data_i({ data_li_1__4__135_, data_li_1__4__134_, data_li_1__4__133_, data_li_1__4__132_, data_li_1__4__131_, data_li_1__4__130_, data_li_1__4__129_, data_li_1__4__128_, data_li_1__4__127_, data_li_1__4__126_, data_li_1__4__125_, data_li_1__4__124_, data_li_1__4__123_, data_li_1__4__122_, data_li_1__4__121_, data_li_1__4__120_, data_li_1__4__119_, data_li_1__4__118_, data_li_1__4__117_, data_li_1__4__116_, data_li_1__4__115_, data_li_1__4__114_, data_li_1__4__113_, data_li_1__4__112_, data_li_1__4__111_, data_li_1__4__110_, data_li_1__4__109_, data_li_1__4__108_, data_li_1__4__107_, data_li_1__4__106_, data_li_1__4__105_, data_li_1__4__104_, data_li_1__4__103_, data_li_1__4__102_, data_li_1__4__101_, data_li_1__4__100_, data_li_1__4__99_, data_li_1__4__98_, data_li_1__4__97_, data_li_1__4__96_, data_li_1__4__95_, data_li_1__4__94_, data_li_1__4__93_, data_li_1__4__92_, data_li_1__4__91_, data_li_1__4__90_, data_li_1__4__89_, data_li_1__4__88_, data_li_1__4__87_, data_li_1__4__86_, data_li_1__4__85_, data_li_1__4__84_, data_li_1__4__83_, data_li_1__4__82_, data_li_1__4__81_, data_li_1__4__80_, data_li_1__4__79_, data_li_1__4__78_, data_li_1__4__77_, data_li_1__4__76_, data_li_1__4__75_, data_li_1__4__74_, data_li_1__4__73_, data_li_1__4__72_, data_li_1__4__71_, data_li_1__4__70_, data_li_1__4__69_, data_li_1__4__68_, data_li_1__4__67_, data_li_1__4__66_, data_li_1__4__65_, data_li_1__4__64_, data_li_1__4__63_, data_li_1__4__62_, data_li_1__4__61_, data_li_1__4__60_, data_li_1__4__59_, data_li_1__4__58_, data_li_1__4__57_, data_li_1__4__56_, data_li_1__4__55_, data_li_1__4__54_, data_li_1__4__53_, data_li_1__4__52_, data_li_1__4__51_, data_li_1__4__50_, data_li_1__4__49_, data_li_1__4__48_, data_li_1__4__47_, data_li_1__4__46_, data_li_1__4__45_, data_li_1__4__44_, data_li_1__4__43_, data_li_1__4__42_, data_li_1__4__41_, data_li_1__4__40_, data_li_1__4__39_, data_li_1__4__38_, data_li_1__4__37_, data_li_1__4__36_, data_li_1__4__35_, data_li_1__4__34_, data_li_1__4__33_, data_li_1__4__32_, data_li_1__4__31_, data_li_1__4__30_, data_li_1__4__29_, data_li_1__4__28_, data_li_1__4__27_, data_li_1__4__26_, data_li_1__4__25_, data_li_1__4__24_, data_li_1__4__23_, data_li_1__4__22_, data_li_1__4__21_, data_li_1__4__20_, data_li_1__4__19_, data_li_1__4__18_, data_li_1__4__17_, data_li_1__4__16_, data_li_1__4__15_, data_li_1__4__14_, data_li_1__4__13_, data_li_1__4__12_, data_li_1__4__11_, data_li_1__4__10_, data_li_1__4__9_, data_li_1__4__8_, data_li_1__4__7_, data_li_1__4__6_, data_li_1__4__5_, data_li_1__4__4_, data_li_1__4__3_, data_li_1__4__2_, data_li_1__4__1_, data_li_1__4__0_, data_li_1__3__135_, data_li_1__3__134_, data_li_1__3__133_, data_li_1__3__132_, data_li_1__3__131_, data_li_1__3__130_, data_li_1__3__129_, data_li_1__3__128_, data_li_1__3__127_, data_li_1__3__126_, data_li_1__3__125_, data_li_1__3__124_, data_li_1__3__123_, data_li_1__3__122_, data_li_1__3__121_, data_li_1__3__120_, data_li_1__3__119_, data_li_1__3__118_, data_li_1__3__117_, data_li_1__3__116_, data_li_1__3__115_, data_li_1__3__114_, data_li_1__3__113_, data_li_1__3__112_, data_li_1__3__111_, data_li_1__3__110_, data_li_1__3__109_, data_li_1__3__108_, data_li_1__3__107_, data_li_1__3__106_, data_li_1__3__105_, data_li_1__3__104_, data_li_1__3__103_, data_li_1__3__102_, data_li_1__3__101_, data_li_1__3__100_, data_li_1__3__99_, data_li_1__3__98_, data_li_1__3__97_, data_li_1__3__96_, data_li_1__3__95_, data_li_1__3__94_, data_li_1__3__93_, data_li_1__3__92_, data_li_1__3__91_, data_li_1__3__90_, data_li_1__3__89_, data_li_1__3__88_, data_li_1__3__87_, data_li_1__3__86_, data_li_1__3__85_, data_li_1__3__84_, data_li_1__3__83_, data_li_1__3__82_, data_li_1__3__81_, data_li_1__3__80_, data_li_1__3__79_, data_li_1__3__78_, data_li_1__3__77_, data_li_1__3__76_, data_li_1__3__75_, data_li_1__3__74_, data_li_1__3__73_, data_li_1__3__72_, data_li_1__3__71_, data_li_1__3__70_, data_li_1__3__69_, data_li_1__3__68_, data_li_1__3__67_, data_li_1__3__66_, data_li_1__3__65_, data_li_1__3__64_, data_li_1__3__63_, data_li_1__3__62_, data_li_1__3__61_, data_li_1__3__60_, data_li_1__3__59_, data_li_1__3__58_, data_li_1__3__57_, data_li_1__3__56_, data_li_1__3__55_, data_li_1__3__54_, data_li_1__3__53_, data_li_1__3__52_, data_li_1__3__51_, data_li_1__3__50_, data_li_1__3__49_, data_li_1__3__48_, data_li_1__3__47_, data_li_1__3__46_, data_li_1__3__45_, data_li_1__3__44_, data_li_1__3__43_, data_li_1__3__42_, data_li_1__3__41_, data_li_1__3__40_, data_li_1__3__39_, data_li_1__3__38_, data_li_1__3__37_, data_li_1__3__36_, data_li_1__3__35_, data_li_1__3__34_, data_li_1__3__33_, data_li_1__3__32_, data_li_1__3__31_, data_li_1__3__30_, data_li_1__3__29_, data_li_1__3__28_, data_li_1__3__27_, data_li_1__3__26_, data_li_1__3__25_, data_li_1__3__24_, data_li_1__3__23_, data_li_1__3__22_, data_li_1__3__21_, data_li_1__3__20_, data_li_1__3__19_, data_li_1__3__18_, data_li_1__3__17_, data_li_1__3__16_, data_li_1__3__15_, data_li_1__3__14_, data_li_1__3__13_, data_li_1__3__12_, data_li_1__3__11_, data_li_1__3__10_, data_li_1__3__9_, data_li_1__3__8_, data_li_1__3__7_, data_li_1__3__6_, data_li_1__3__5_, data_li_1__3__4_, data_li_1__3__3_, data_li_1__3__2_, data_li_1__3__1_, data_li_1__3__0_, data_li_1__2__135_, data_li_1__2__134_, data_li_1__2__133_, data_li_1__2__132_, data_li_1__2__131_, data_li_1__2__130_, data_li_1__2__129_, data_li_1__2__128_, data_li_1__2__127_, data_li_1__2__126_, data_li_1__2__125_, data_li_1__2__124_, data_li_1__2__123_, data_li_1__2__122_, data_li_1__2__121_, data_li_1__2__120_, data_li_1__2__119_, data_li_1__2__118_, data_li_1__2__117_, data_li_1__2__116_, data_li_1__2__115_, data_li_1__2__114_, data_li_1__2__113_, data_li_1__2__112_, data_li_1__2__111_, data_li_1__2__110_, data_li_1__2__109_, data_li_1__2__108_, data_li_1__2__107_, data_li_1__2__106_, data_li_1__2__105_, data_li_1__2__104_, data_li_1__2__103_, data_li_1__2__102_, data_li_1__2__101_, data_li_1__2__100_, data_li_1__2__99_, data_li_1__2__98_, data_li_1__2__97_, data_li_1__2__96_, data_li_1__2__95_, data_li_1__2__94_, data_li_1__2__93_, data_li_1__2__92_, data_li_1__2__91_, data_li_1__2__90_, data_li_1__2__89_, data_li_1__2__88_, data_li_1__2__87_, data_li_1__2__86_, data_li_1__2__85_, data_li_1__2__84_, data_li_1__2__83_, data_li_1__2__82_, data_li_1__2__81_, data_li_1__2__80_, data_li_1__2__79_, data_li_1__2__78_, data_li_1__2__77_, data_li_1__2__76_, data_li_1__2__75_, data_li_1__2__74_, data_li_1__2__73_, data_li_1__2__72_, data_li_1__2__71_, data_li_1__2__70_, data_li_1__2__69_, data_li_1__2__68_, data_li_1__2__67_, data_li_1__2__66_, data_li_1__2__65_, data_li_1__2__64_, data_li_1__2__63_, data_li_1__2__62_, data_li_1__2__61_, data_li_1__2__60_, data_li_1__2__59_, data_li_1__2__58_, data_li_1__2__57_, data_li_1__2__56_, data_li_1__2__55_, data_li_1__2__54_, data_li_1__2__53_, data_li_1__2__52_, data_li_1__2__51_, data_li_1__2__50_, data_li_1__2__49_, data_li_1__2__48_, data_li_1__2__47_, data_li_1__2__46_, data_li_1__2__45_, data_li_1__2__44_, data_li_1__2__43_, data_li_1__2__42_, data_li_1__2__41_, data_li_1__2__40_, data_li_1__2__39_, data_li_1__2__38_, data_li_1__2__37_, data_li_1__2__36_, data_li_1__2__35_, data_li_1__2__34_, data_li_1__2__33_, data_li_1__2__32_, data_li_1__2__31_, data_li_1__2__30_, data_li_1__2__29_, data_li_1__2__28_, data_li_1__2__27_, data_li_1__2__26_, data_li_1__2__25_, data_li_1__2__24_, data_li_1__2__23_, data_li_1__2__22_, data_li_1__2__21_, data_li_1__2__20_, data_li_1__2__19_, data_li_1__2__18_, data_li_1__2__17_, data_li_1__2__16_, data_li_1__2__15_, data_li_1__2__14_, data_li_1__2__13_, data_li_1__2__12_, data_li_1__2__11_, data_li_1__2__10_, data_li_1__2__9_, data_li_1__2__8_, data_li_1__2__7_, data_li_1__2__6_, data_li_1__2__5_, data_li_1__2__4_, data_li_1__2__3_, data_li_1__2__2_, data_li_1__2__1_, data_li_1__2__0_, data_lo[407:272], data_li_1__0__135_, data_li_1__0__134_, data_li_1__0__133_, data_li_1__0__132_, data_li_1__0__131_, data_li_1__0__130_, data_li_1__0__129_, data_li_1__0__128_, data_li_1__0__127_, data_li_1__0__126_, data_li_1__0__125_, data_li_1__0__124_, data_li_1__0__123_, data_li_1__0__122_, data_li_1__0__121_, data_li_1__0__120_, data_li_1__0__119_, data_li_1__0__118_, data_li_1__0__117_, data_li_1__0__116_, data_li_1__0__115_, data_li_1__0__114_, data_li_1__0__113_, data_li_1__0__112_, data_li_1__0__111_, data_li_1__0__110_, data_li_1__0__109_, data_li_1__0__108_, data_li_1__0__107_, data_li_1__0__106_, data_li_1__0__105_, data_li_1__0__104_, data_li_1__0__103_, data_li_1__0__102_, data_li_1__0__101_, data_li_1__0__100_, data_li_1__0__99_, data_li_1__0__98_, data_li_1__0__97_, data_li_1__0__96_, data_li_1__0__95_, data_li_1__0__94_, data_li_1__0__93_, data_li_1__0__92_, data_li_1__0__91_, data_li_1__0__90_, data_li_1__0__89_, data_li_1__0__88_, data_li_1__0__87_, data_li_1__0__86_, data_li_1__0__85_, data_li_1__0__84_, data_li_1__0__83_, data_li_1__0__82_, data_li_1__0__81_, data_li_1__0__80_, data_li_1__0__79_, data_li_1__0__78_, data_li_1__0__77_, data_li_1__0__76_, data_li_1__0__75_, data_li_1__0__74_, data_li_1__0__73_, data_li_1__0__72_, data_li_1__0__71_, data_li_1__0__70_, data_li_1__0__69_, data_li_1__0__68_, data_li_1__0__67_, data_li_1__0__66_, data_li_1__0__65_, data_li_1__0__64_, data_li_1__0__63_, data_li_1__0__62_, data_li_1__0__61_, data_li_1__0__60_, data_li_1__0__59_, data_li_1__0__58_, data_li_1__0__57_, data_li_1__0__56_, data_li_1__0__55_, data_li_1__0__54_, data_li_1__0__53_, data_li_1__0__52_, data_li_1__0__51_, data_li_1__0__50_, data_li_1__0__49_, data_li_1__0__48_, data_li_1__0__47_, data_li_1__0__46_, data_li_1__0__45_, data_li_1__0__44_, data_li_1__0__43_, data_li_1__0__42_, data_li_1__0__41_, data_li_1__0__40_, data_li_1__0__39_, data_li_1__0__38_, data_li_1__0__37_, data_li_1__0__36_, data_li_1__0__35_, data_li_1__0__34_, data_li_1__0__33_, data_li_1__0__32_, data_li_1__0__31_, data_li_1__0__30_, data_li_1__0__29_, data_li_1__0__28_, data_li_1__0__27_, data_li_1__0__26_, data_li_1__0__25_, data_li_1__0__24_, data_li_1__0__23_, data_li_1__0__22_, data_li_1__0__21_, data_li_1__0__20_, data_li_1__0__19_, data_li_1__0__18_, data_li_1__0__17_, data_li_1__0__16_, data_li_1__0__15_, data_li_1__0__14_, data_li_1__0__13_, data_li_1__0__12_, data_li_1__0__11_, data_li_1__0__10_, data_li_1__0__9_, data_li_1__0__8_, data_li_1__0__7_, data_li_1__0__6_, data_li_1__0__5_, data_li_1__0__4_, data_li_1__0__3_, data_li_1__0__2_, data_li_1__0__1_, data_li_1__0__0_ }),
    .ready_o(ready_lo[9:5]),
    .valid_o(valid_lo[9:5]),
    .data_o(data_lo[1359:680]),
    .ready_i({ ready_li_1__4_, ready_li_1__3_, ready_li_1__2_, ready_lo[2:2], ready_li_1__0_ })
  );


  bp_me_network_pkt_encode_data_resp_num_lce_p2_num_cce_p1_paddr_width_p22_block_size_in_bits_p512_max_num_flit_p4_x_cord_width_p1_y_cord_width_p1
  genblk3_0__pkt_encode
  (
    .payload_i(lce_data_resp_i[536:0]),
    .packet_o(lce_packet[540:0])
  );


  bp_me_network_pkt_encode_data_resp_num_lce_p2_num_cce_p1_paddr_width_p22_block_size_in_bits_p512_max_num_flit_p4_x_cord_width_p1_y_cord_width_p1
  genblk3_1__pkt_encode
  (
    .payload_i(lce_data_resp_i[1073:537]),
    .packet_o(lce_packet[1081:541])
  );


  bsg_wormhole_router_adapter_in_max_num_flit_p4_max_payload_width_p537_x_cord_width_p1_y_cord_width_p1
  genblk4_0__adapter_in
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(lce_packet[540:0]),
    .v_i(lce_data_resp_v_i[0]),
    .ready_o(lce_data_resp_ready_o[0]),
    .data_o({ data_li_0__3__135_, data_li_0__3__134_, data_li_0__3__133_, data_li_0__3__132_, data_li_0__3__131_, data_li_0__3__130_, data_li_0__3__129_, data_li_0__3__128_, data_li_0__3__127_, data_li_0__3__126_, data_li_0__3__125_, data_li_0__3__124_, data_li_0__3__123_, data_li_0__3__122_, data_li_0__3__121_, data_li_0__3__120_, data_li_0__3__119_, data_li_0__3__118_, data_li_0__3__117_, data_li_0__3__116_, data_li_0__3__115_, data_li_0__3__114_, data_li_0__3__113_, data_li_0__3__112_, data_li_0__3__111_, data_li_0__3__110_, data_li_0__3__109_, data_li_0__3__108_, data_li_0__3__107_, data_li_0__3__106_, data_li_0__3__105_, data_li_0__3__104_, data_li_0__3__103_, data_li_0__3__102_, data_li_0__3__101_, data_li_0__3__100_, data_li_0__3__99_, data_li_0__3__98_, data_li_0__3__97_, data_li_0__3__96_, data_li_0__3__95_, data_li_0__3__94_, data_li_0__3__93_, data_li_0__3__92_, data_li_0__3__91_, data_li_0__3__90_, data_li_0__3__89_, data_li_0__3__88_, data_li_0__3__87_, data_li_0__3__86_, data_li_0__3__85_, data_li_0__3__84_, data_li_0__3__83_, data_li_0__3__82_, data_li_0__3__81_, data_li_0__3__80_, data_li_0__3__79_, data_li_0__3__78_, data_li_0__3__77_, data_li_0__3__76_, data_li_0__3__75_, data_li_0__3__74_, data_li_0__3__73_, data_li_0__3__72_, data_li_0__3__71_, data_li_0__3__70_, data_li_0__3__69_, data_li_0__3__68_, data_li_0__3__67_, data_li_0__3__66_, data_li_0__3__65_, data_li_0__3__64_, data_li_0__3__63_, data_li_0__3__62_, data_li_0__3__61_, data_li_0__3__60_, data_li_0__3__59_, data_li_0__3__58_, data_li_0__3__57_, data_li_0__3__56_, data_li_0__3__55_, data_li_0__3__54_, data_li_0__3__53_, data_li_0__3__52_, data_li_0__3__51_, data_li_0__3__50_, data_li_0__3__49_, data_li_0__3__48_, data_li_0__3__47_, data_li_0__3__46_, data_li_0__3__45_, data_li_0__3__44_, data_li_0__3__43_, data_li_0__3__42_, data_li_0__3__41_, data_li_0__3__40_, data_li_0__3__39_, data_li_0__3__38_, data_li_0__3__37_, data_li_0__3__36_, data_li_0__3__35_, data_li_0__3__34_, data_li_0__3__33_, data_li_0__3__32_, data_li_0__3__31_, data_li_0__3__30_, data_li_0__3__29_, data_li_0__3__28_, data_li_0__3__27_, data_li_0__3__26_, data_li_0__3__25_, data_li_0__3__24_, data_li_0__3__23_, data_li_0__3__22_, data_li_0__3__21_, data_li_0__3__20_, data_li_0__3__19_, data_li_0__3__18_, data_li_0__3__17_, data_li_0__3__16_, data_li_0__3__15_, data_li_0__3__14_, data_li_0__3__13_, data_li_0__3__12_, data_li_0__3__11_, data_li_0__3__10_, data_li_0__3__9_, data_li_0__3__8_, data_li_0__3__7_, data_li_0__3__6_, data_li_0__3__5_, data_li_0__3__4_, data_li_0__3__3_, data_li_0__3__2_, data_li_0__3__1_, data_li_0__3__0_ }),
    .v_o(valid_li_0__3_),
    .ready_i(ready_lo[3])
  );


  bsg_wormhole_router_adapter_in_max_num_flit_p4_max_payload_width_p537_x_cord_width_p1_y_cord_width_p1
  genblk4_1__adapter_in
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(lce_packet[1081:541]),
    .v_i(lce_data_resp_v_i[1]),
    .ready_o(lce_data_resp_ready_o[1]),
    .data_o({ data_li_1__3__135_, data_li_1__3__134_, data_li_1__3__133_, data_li_1__3__132_, data_li_1__3__131_, data_li_1__3__130_, data_li_1__3__129_, data_li_1__3__128_, data_li_1__3__127_, data_li_1__3__126_, data_li_1__3__125_, data_li_1__3__124_, data_li_1__3__123_, data_li_1__3__122_, data_li_1__3__121_, data_li_1__3__120_, data_li_1__3__119_, data_li_1__3__118_, data_li_1__3__117_, data_li_1__3__116_, data_li_1__3__115_, data_li_1__3__114_, data_li_1__3__113_, data_li_1__3__112_, data_li_1__3__111_, data_li_1__3__110_, data_li_1__3__109_, data_li_1__3__108_, data_li_1__3__107_, data_li_1__3__106_, data_li_1__3__105_, data_li_1__3__104_, data_li_1__3__103_, data_li_1__3__102_, data_li_1__3__101_, data_li_1__3__100_, data_li_1__3__99_, data_li_1__3__98_, data_li_1__3__97_, data_li_1__3__96_, data_li_1__3__95_, data_li_1__3__94_, data_li_1__3__93_, data_li_1__3__92_, data_li_1__3__91_, data_li_1__3__90_, data_li_1__3__89_, data_li_1__3__88_, data_li_1__3__87_, data_li_1__3__86_, data_li_1__3__85_, data_li_1__3__84_, data_li_1__3__83_, data_li_1__3__82_, data_li_1__3__81_, data_li_1__3__80_, data_li_1__3__79_, data_li_1__3__78_, data_li_1__3__77_, data_li_1__3__76_, data_li_1__3__75_, data_li_1__3__74_, data_li_1__3__73_, data_li_1__3__72_, data_li_1__3__71_, data_li_1__3__70_, data_li_1__3__69_, data_li_1__3__68_, data_li_1__3__67_, data_li_1__3__66_, data_li_1__3__65_, data_li_1__3__64_, data_li_1__3__63_, data_li_1__3__62_, data_li_1__3__61_, data_li_1__3__60_, data_li_1__3__59_, data_li_1__3__58_, data_li_1__3__57_, data_li_1__3__56_, data_li_1__3__55_, data_li_1__3__54_, data_li_1__3__53_, data_li_1__3__52_, data_li_1__3__51_, data_li_1__3__50_, data_li_1__3__49_, data_li_1__3__48_, data_li_1__3__47_, data_li_1__3__46_, data_li_1__3__45_, data_li_1__3__44_, data_li_1__3__43_, data_li_1__3__42_, data_li_1__3__41_, data_li_1__3__40_, data_li_1__3__39_, data_li_1__3__38_, data_li_1__3__37_, data_li_1__3__36_, data_li_1__3__35_, data_li_1__3__34_, data_li_1__3__33_, data_li_1__3__32_, data_li_1__3__31_, data_li_1__3__30_, data_li_1__3__29_, data_li_1__3__28_, data_li_1__3__27_, data_li_1__3__26_, data_li_1__3__25_, data_li_1__3__24_, data_li_1__3__23_, data_li_1__3__22_, data_li_1__3__21_, data_li_1__3__20_, data_li_1__3__19_, data_li_1__3__18_, data_li_1__3__17_, data_li_1__3__16_, data_li_1__3__15_, data_li_1__3__14_, data_li_1__3__13_, data_li_1__3__12_, data_li_1__3__11_, data_li_1__3__10_, data_li_1__3__9_, data_li_1__3__8_, data_li_1__3__7_, data_li_1__3__6_, data_li_1__3__5_, data_li_1__3__4_, data_li_1__3__3_, data_li_1__3__2_, data_li_1__3__1_, data_li_1__3__0_ }),
    .v_o(valid_li_1__3_),
    .ready_i(ready_lo[8])
  );


  bsg_wormhole_router_adapter_out_max_num_flit_p4_max_payload_width_p537_x_cord_width_p1_y_cord_width_p1
  genblk5_0__adapter_out
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_lo[135:0]),
    .v_i(valid_lo[0]),
    .ready_o(ready_li_0__0_),
    .data_o({ lce_data_resp_o, cce_packet_0__3_, cce_packet_0__2_, cce_packet_0__1_, cce_packet_0__0_ }),
    .v_o(lce_data_resp_v_o[0]),
    .ready_i(lce_data_resp_ready_i[0])
  );


endmodule



module bsg_mem_p131
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [130:0] w_data_i;
  input [0:0] r_addr_i;
  output [130:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [130:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10;
  reg [261:0] mem;
  assign r_data_o[130] = (N3)? mem[130] :
                         (N0)? mem[261] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[129] = (N3)? mem[129] :
                         (N0)? mem[260] : 1'b0;
  assign r_data_o[128] = (N3)? mem[128] :
                         (N0)? mem[259] : 1'b0;
  assign r_data_o[127] = (N3)? mem[127] :
                         (N0)? mem[258] : 1'b0;
  assign r_data_o[126] = (N3)? mem[126] :
                         (N0)? mem[257] : 1'b0;
  assign r_data_o[125] = (N3)? mem[125] :
                         (N0)? mem[256] : 1'b0;
  assign r_data_o[124] = (N3)? mem[124] :
                         (N0)? mem[255] : 1'b0;
  assign r_data_o[123] = (N3)? mem[123] :
                         (N0)? mem[254] : 1'b0;
  assign r_data_o[122] = (N3)? mem[122] :
                         (N0)? mem[253] : 1'b0;
  assign r_data_o[121] = (N3)? mem[121] :
                         (N0)? mem[252] : 1'b0;
  assign r_data_o[120] = (N3)? mem[120] :
                         (N0)? mem[251] : 1'b0;
  assign r_data_o[119] = (N3)? mem[119] :
                         (N0)? mem[250] : 1'b0;
  assign r_data_o[118] = (N3)? mem[118] :
                         (N0)? mem[249] : 1'b0;
  assign r_data_o[117] = (N3)? mem[117] :
                         (N0)? mem[248] : 1'b0;
  assign r_data_o[116] = (N3)? mem[116] :
                         (N0)? mem[247] : 1'b0;
  assign r_data_o[115] = (N3)? mem[115] :
                         (N0)? mem[246] : 1'b0;
  assign r_data_o[114] = (N3)? mem[114] :
                         (N0)? mem[245] : 1'b0;
  assign r_data_o[113] = (N3)? mem[113] :
                         (N0)? mem[244] : 1'b0;
  assign r_data_o[112] = (N3)? mem[112] :
                         (N0)? mem[243] : 1'b0;
  assign r_data_o[111] = (N3)? mem[111] :
                         (N0)? mem[242] : 1'b0;
  assign r_data_o[110] = (N3)? mem[110] :
                         (N0)? mem[241] : 1'b0;
  assign r_data_o[109] = (N3)? mem[109] :
                         (N0)? mem[240] : 1'b0;
  assign r_data_o[108] = (N3)? mem[108] :
                         (N0)? mem[239] : 1'b0;
  assign r_data_o[107] = (N3)? mem[107] :
                         (N0)? mem[238] : 1'b0;
  assign r_data_o[106] = (N3)? mem[106] :
                         (N0)? mem[237] : 1'b0;
  assign r_data_o[105] = (N3)? mem[105] :
                         (N0)? mem[236] : 1'b0;
  assign r_data_o[104] = (N3)? mem[104] :
                         (N0)? mem[235] : 1'b0;
  assign r_data_o[103] = (N3)? mem[103] :
                         (N0)? mem[234] : 1'b0;
  assign r_data_o[102] = (N3)? mem[102] :
                         (N0)? mem[233] : 1'b0;
  assign r_data_o[101] = (N3)? mem[101] :
                         (N0)? mem[232] : 1'b0;
  assign r_data_o[100] = (N3)? mem[100] :
                         (N0)? mem[231] : 1'b0;
  assign r_data_o[99] = (N3)? mem[99] :
                        (N0)? mem[230] : 1'b0;
  assign r_data_o[98] = (N3)? mem[98] :
                        (N0)? mem[229] : 1'b0;
  assign r_data_o[97] = (N3)? mem[97] :
                        (N0)? mem[228] : 1'b0;
  assign r_data_o[96] = (N3)? mem[96] :
                        (N0)? mem[227] : 1'b0;
  assign r_data_o[95] = (N3)? mem[95] :
                        (N0)? mem[226] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] :
                        (N0)? mem[225] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] :
                        (N0)? mem[224] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] :
                        (N0)? mem[223] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] :
                        (N0)? mem[222] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] :
                        (N0)? mem[221] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] :
                        (N0)? mem[220] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] :
                        (N0)? mem[219] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] :
                        (N0)? mem[218] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] :
                        (N0)? mem[217] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] :
                        (N0)? mem[216] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] :
                        (N0)? mem[215] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] :
                        (N0)? mem[214] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] :
                        (N0)? mem[213] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] :
                        (N0)? mem[212] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] :
                        (N0)? mem[211] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] :
                        (N0)? mem[210] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] :
                        (N0)? mem[209] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] :
                        (N0)? mem[208] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] :
                        (N0)? mem[207] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] :
                        (N0)? mem[206] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] :
                        (N0)? mem[205] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] :
                        (N0)? mem[204] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] :
                        (N0)? mem[203] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] :
                        (N0)? mem[202] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] :
                        (N0)? mem[201] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] :
                        (N0)? mem[200] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] :
                        (N0)? mem[199] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] :
                        (N0)? mem[198] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] :
                        (N0)? mem[197] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] :
                        (N0)? mem[196] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] :
                        (N0)? mem[195] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] :
                        (N0)? mem[194] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] :
                        (N0)? mem[193] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] :
                        (N0)? mem[192] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] :
                        (N0)? mem[191] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] :
                        (N0)? mem[190] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] :
                        (N0)? mem[189] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] :
                        (N0)? mem[188] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] :
                        (N0)? mem[187] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] :
                        (N0)? mem[186] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] :
                        (N0)? mem[185] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] :
                        (N0)? mem[184] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] :
                        (N0)? mem[183] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] :
                        (N0)? mem[182] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] :
                        (N0)? mem[181] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] :
                        (N0)? mem[180] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] :
                        (N0)? mem[179] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] :
                        (N0)? mem[178] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] :
                        (N0)? mem[177] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] :
                        (N0)? mem[176] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] :
                        (N0)? mem[175] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] :
                        (N0)? mem[174] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] :
                        (N0)? mem[173] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] :
                        (N0)? mem[172] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] :
                        (N0)? mem[171] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] :
                        (N0)? mem[170] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] :
                        (N0)? mem[169] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] :
                        (N0)? mem[168] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] :
                        (N0)? mem[167] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] :
                        (N0)? mem[166] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] :
                        (N0)? mem[165] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] :
                        (N0)? mem[164] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] :
                        (N0)? mem[163] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] :
                        (N0)? mem[162] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] :
                        (N0)? mem[161] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] :
                        (N0)? mem[160] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] :
                        (N0)? mem[159] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] :
                        (N0)? mem[158] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] :
                        (N0)? mem[157] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] :
                        (N0)? mem[156] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] :
                        (N0)? mem[155] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] :
                        (N0)? mem[154] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] :
                        (N0)? mem[153] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] :
                        (N0)? mem[152] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] :
                        (N0)? mem[151] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] :
                        (N0)? mem[150] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] :
                        (N0)? mem[149] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] :
                        (N0)? mem[148] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] :
                        (N0)? mem[147] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] :
                        (N0)? mem[146] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] :
                        (N0)? mem[145] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] :
                        (N0)? mem[144] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] :
                        (N0)? mem[143] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] :
                        (N0)? mem[142] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] :
                        (N0)? mem[141] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] :
                       (N0)? mem[140] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] :
                       (N0)? mem[139] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] :
                       (N0)? mem[138] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] :
                       (N0)? mem[137] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] :
                       (N0)? mem[136] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] :
                       (N0)? mem[135] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] :
                       (N0)? mem[134] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] :
                       (N0)? mem[133] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] :
                       (N0)? mem[132] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] :
                       (N0)? mem[131] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], N5, N5 } :
                               (N2)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N9) begin
      { mem[261:163], mem[131:131] } <= { w_data_i[130:32], w_data_i[0:0] };
    end
    if(N10) begin
      { mem[162:132] } <= { w_data_i[31:1] };
    end
    if(N7) begin
      { mem[130:32], mem[0:0] } <= { w_data_i[130:32], w_data_i[0:0] };
    end
    if(N8) begin
      { mem[31:1] } <= { w_data_i[31:1] };
    end
  end


endmodule



module bsg_mem_1r1w_width_p131_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [130:0] w_data_i;
  input [0:0] r_addr_i;
  output [130:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [130:0] r_data_o;

  bsg_mem_p131
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p131
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [130:0] data_i;
  output [130:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [130:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p131_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 :
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 :
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 :
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 :
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 :
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 :
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end
    if(N9) begin
      tail_r <= N10;
    end
    if(N11) begin
      head_r <= N12;
    end
  end


endmodule



module bsg_mux_one_hot_width_p131_els_p4
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [523:0] data_i;
  input [3:0] sel_one_hot_i;
  output [130:0] data_o;
  wire [130:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261;
  wire [523:0] data_masked;
  assign data_masked[130] = data_i[130] & sel_one_hot_i[0];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[0];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[0];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[0];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[0];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[0];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[0];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[0];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[0];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[0];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[0];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[0];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[0];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[0];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[0];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[0];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[0];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[0];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[0];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[0];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[0];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[0];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[0];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[0];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[0];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[0];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[0];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[0];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[0];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[0];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[0];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[0];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[0];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[0];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[0];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[0];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[0];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[0];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[0];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[0];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[0];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[0];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[0];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[0];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[0];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[0];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[0];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[0];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[0];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[0];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[0];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[0];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[0];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[0];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[0];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[0];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[0];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[0];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[0];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[0];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[0];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[0];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[0];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[1];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[1];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[1];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[1];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[1];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[1];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[1];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[1];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[1];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[1];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[1];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[1];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[1];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[1];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[1];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[1];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[1];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[1];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[1];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[1];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[1];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[1];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[1];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[1];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[1];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[1];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[1];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[1];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[1];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[1];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[1];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[1];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[1];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[1];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[1];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[1];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[1];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[1];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[1];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[1];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[1];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[1];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[1];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[1];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[1];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[1];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[1];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[1];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[1];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[1];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[1];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[1];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[1];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[1];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[1];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[1];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[1];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[1];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[1];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[1];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[1];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[1];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[1];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[1];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[1];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[1];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[1];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[1];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[1];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[1];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[1];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[1];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[1];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[1];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[1];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[1];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[1];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[1];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[1];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[1];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[1];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[1];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[1];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[1];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[1];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[1];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[1];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[1];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[1];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[1];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[1];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[1];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[1];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[1];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[1];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[1];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[1];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[1];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[1];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[1];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[1];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[1];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[1];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[1];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[1];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[1];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[1];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[1];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[1];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[1];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[1];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[1];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[1];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[1];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[1];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[1];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[1];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[1];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[1];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[1];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[1];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[1];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[1];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[1];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[1];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[1];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[1];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[1];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[1];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[1];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[2];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[2];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[2];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[2];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[2];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[2];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[2];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[2];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[2];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[2];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[2];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[2];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[2];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[2];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[2];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[2];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[2];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[2];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[2];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[2];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[2];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[2];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[2];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[2];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[2];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[2];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[2];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[2];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[2];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[2];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[2];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[2];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[2];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[2];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[2];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[2];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[2];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[2];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[2];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[2];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[2];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[2];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[2];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[2];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[2];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[2];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[2];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[2];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[2];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[2];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[2];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[2];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[2];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[2];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[2];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[2];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[2];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[2];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[2];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[2];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[2];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[2];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[2];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[2];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[2];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[2];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[2];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[2];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[2];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[2];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[2];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[2];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[2];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[2];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[2];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[2];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[2];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[2];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[2];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[2];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[2];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[2];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[2];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[2];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[2];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[2];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[2];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[2];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[2];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[2];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[2];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[2];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[2];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[2];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[2];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[2];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[2];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[2];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[2];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[2];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[2];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[2];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[2];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[2];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[2];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[2];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[2];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[2];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[2];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[2];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[2];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[2];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[2];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[2];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[2];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[2];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[2];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[2];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[2];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[2];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[2];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[2];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[2];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[2];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[2];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[2];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[2];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[2];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[2];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[2];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[2];
  assign data_masked[523] = data_i[523] & sel_one_hot_i[3];
  assign data_masked[522] = data_i[522] & sel_one_hot_i[3];
  assign data_masked[521] = data_i[521] & sel_one_hot_i[3];
  assign data_masked[520] = data_i[520] & sel_one_hot_i[3];
  assign data_masked[519] = data_i[519] & sel_one_hot_i[3];
  assign data_masked[518] = data_i[518] & sel_one_hot_i[3];
  assign data_masked[517] = data_i[517] & sel_one_hot_i[3];
  assign data_masked[516] = data_i[516] & sel_one_hot_i[3];
  assign data_masked[515] = data_i[515] & sel_one_hot_i[3];
  assign data_masked[514] = data_i[514] & sel_one_hot_i[3];
  assign data_masked[513] = data_i[513] & sel_one_hot_i[3];
  assign data_masked[512] = data_i[512] & sel_one_hot_i[3];
  assign data_masked[511] = data_i[511] & sel_one_hot_i[3];
  assign data_masked[510] = data_i[510] & sel_one_hot_i[3];
  assign data_masked[509] = data_i[509] & sel_one_hot_i[3];
  assign data_masked[508] = data_i[508] & sel_one_hot_i[3];
  assign data_masked[507] = data_i[507] & sel_one_hot_i[3];
  assign data_masked[506] = data_i[506] & sel_one_hot_i[3];
  assign data_masked[505] = data_i[505] & sel_one_hot_i[3];
  assign data_masked[504] = data_i[504] & sel_one_hot_i[3];
  assign data_masked[503] = data_i[503] & sel_one_hot_i[3];
  assign data_masked[502] = data_i[502] & sel_one_hot_i[3];
  assign data_masked[501] = data_i[501] & sel_one_hot_i[3];
  assign data_masked[500] = data_i[500] & sel_one_hot_i[3];
  assign data_masked[499] = data_i[499] & sel_one_hot_i[3];
  assign data_masked[498] = data_i[498] & sel_one_hot_i[3];
  assign data_masked[497] = data_i[497] & sel_one_hot_i[3];
  assign data_masked[496] = data_i[496] & sel_one_hot_i[3];
  assign data_masked[495] = data_i[495] & sel_one_hot_i[3];
  assign data_masked[494] = data_i[494] & sel_one_hot_i[3];
  assign data_masked[493] = data_i[493] & sel_one_hot_i[3];
  assign data_masked[492] = data_i[492] & sel_one_hot_i[3];
  assign data_masked[491] = data_i[491] & sel_one_hot_i[3];
  assign data_masked[490] = data_i[490] & sel_one_hot_i[3];
  assign data_masked[489] = data_i[489] & sel_one_hot_i[3];
  assign data_masked[488] = data_i[488] & sel_one_hot_i[3];
  assign data_masked[487] = data_i[487] & sel_one_hot_i[3];
  assign data_masked[486] = data_i[486] & sel_one_hot_i[3];
  assign data_masked[485] = data_i[485] & sel_one_hot_i[3];
  assign data_masked[484] = data_i[484] & sel_one_hot_i[3];
  assign data_masked[483] = data_i[483] & sel_one_hot_i[3];
  assign data_masked[482] = data_i[482] & sel_one_hot_i[3];
  assign data_masked[481] = data_i[481] & sel_one_hot_i[3];
  assign data_masked[480] = data_i[480] & sel_one_hot_i[3];
  assign data_masked[479] = data_i[479] & sel_one_hot_i[3];
  assign data_masked[478] = data_i[478] & sel_one_hot_i[3];
  assign data_masked[477] = data_i[477] & sel_one_hot_i[3];
  assign data_masked[476] = data_i[476] & sel_one_hot_i[3];
  assign data_masked[475] = data_i[475] & sel_one_hot_i[3];
  assign data_masked[474] = data_i[474] & sel_one_hot_i[3];
  assign data_masked[473] = data_i[473] & sel_one_hot_i[3];
  assign data_masked[472] = data_i[472] & sel_one_hot_i[3];
  assign data_masked[471] = data_i[471] & sel_one_hot_i[3];
  assign data_masked[470] = data_i[470] & sel_one_hot_i[3];
  assign data_masked[469] = data_i[469] & sel_one_hot_i[3];
  assign data_masked[468] = data_i[468] & sel_one_hot_i[3];
  assign data_masked[467] = data_i[467] & sel_one_hot_i[3];
  assign data_masked[466] = data_i[466] & sel_one_hot_i[3];
  assign data_masked[465] = data_i[465] & sel_one_hot_i[3];
  assign data_masked[464] = data_i[464] & sel_one_hot_i[3];
  assign data_masked[463] = data_i[463] & sel_one_hot_i[3];
  assign data_masked[462] = data_i[462] & sel_one_hot_i[3];
  assign data_masked[461] = data_i[461] & sel_one_hot_i[3];
  assign data_masked[460] = data_i[460] & sel_one_hot_i[3];
  assign data_masked[459] = data_i[459] & sel_one_hot_i[3];
  assign data_masked[458] = data_i[458] & sel_one_hot_i[3];
  assign data_masked[457] = data_i[457] & sel_one_hot_i[3];
  assign data_masked[456] = data_i[456] & sel_one_hot_i[3];
  assign data_masked[455] = data_i[455] & sel_one_hot_i[3];
  assign data_masked[454] = data_i[454] & sel_one_hot_i[3];
  assign data_masked[453] = data_i[453] & sel_one_hot_i[3];
  assign data_masked[452] = data_i[452] & sel_one_hot_i[3];
  assign data_masked[451] = data_i[451] & sel_one_hot_i[3];
  assign data_masked[450] = data_i[450] & sel_one_hot_i[3];
  assign data_masked[449] = data_i[449] & sel_one_hot_i[3];
  assign data_masked[448] = data_i[448] & sel_one_hot_i[3];
  assign data_masked[447] = data_i[447] & sel_one_hot_i[3];
  assign data_masked[446] = data_i[446] & sel_one_hot_i[3];
  assign data_masked[445] = data_i[445] & sel_one_hot_i[3];
  assign data_masked[444] = data_i[444] & sel_one_hot_i[3];
  assign data_masked[443] = data_i[443] & sel_one_hot_i[3];
  assign data_masked[442] = data_i[442] & sel_one_hot_i[3];
  assign data_masked[441] = data_i[441] & sel_one_hot_i[3];
  assign data_masked[440] = data_i[440] & sel_one_hot_i[3];
  assign data_masked[439] = data_i[439] & sel_one_hot_i[3];
  assign data_masked[438] = data_i[438] & sel_one_hot_i[3];
  assign data_masked[437] = data_i[437] & sel_one_hot_i[3];
  assign data_masked[436] = data_i[436] & sel_one_hot_i[3];
  assign data_masked[435] = data_i[435] & sel_one_hot_i[3];
  assign data_masked[434] = data_i[434] & sel_one_hot_i[3];
  assign data_masked[433] = data_i[433] & sel_one_hot_i[3];
  assign data_masked[432] = data_i[432] & sel_one_hot_i[3];
  assign data_masked[431] = data_i[431] & sel_one_hot_i[3];
  assign data_masked[430] = data_i[430] & sel_one_hot_i[3];
  assign data_masked[429] = data_i[429] & sel_one_hot_i[3];
  assign data_masked[428] = data_i[428] & sel_one_hot_i[3];
  assign data_masked[427] = data_i[427] & sel_one_hot_i[3];
  assign data_masked[426] = data_i[426] & sel_one_hot_i[3];
  assign data_masked[425] = data_i[425] & sel_one_hot_i[3];
  assign data_masked[424] = data_i[424] & sel_one_hot_i[3];
  assign data_masked[423] = data_i[423] & sel_one_hot_i[3];
  assign data_masked[422] = data_i[422] & sel_one_hot_i[3];
  assign data_masked[421] = data_i[421] & sel_one_hot_i[3];
  assign data_masked[420] = data_i[420] & sel_one_hot_i[3];
  assign data_masked[419] = data_i[419] & sel_one_hot_i[3];
  assign data_masked[418] = data_i[418] & sel_one_hot_i[3];
  assign data_masked[417] = data_i[417] & sel_one_hot_i[3];
  assign data_masked[416] = data_i[416] & sel_one_hot_i[3];
  assign data_masked[415] = data_i[415] & sel_one_hot_i[3];
  assign data_masked[414] = data_i[414] & sel_one_hot_i[3];
  assign data_masked[413] = data_i[413] & sel_one_hot_i[3];
  assign data_masked[412] = data_i[412] & sel_one_hot_i[3];
  assign data_masked[411] = data_i[411] & sel_one_hot_i[3];
  assign data_masked[410] = data_i[410] & sel_one_hot_i[3];
  assign data_masked[409] = data_i[409] & sel_one_hot_i[3];
  assign data_masked[408] = data_i[408] & sel_one_hot_i[3];
  assign data_masked[407] = data_i[407] & sel_one_hot_i[3];
  assign data_masked[406] = data_i[406] & sel_one_hot_i[3];
  assign data_masked[405] = data_i[405] & sel_one_hot_i[3];
  assign data_masked[404] = data_i[404] & sel_one_hot_i[3];
  assign data_masked[403] = data_i[403] & sel_one_hot_i[3];
  assign data_masked[402] = data_i[402] & sel_one_hot_i[3];
  assign data_masked[401] = data_i[401] & sel_one_hot_i[3];
  assign data_masked[400] = data_i[400] & sel_one_hot_i[3];
  assign data_masked[399] = data_i[399] & sel_one_hot_i[3];
  assign data_masked[398] = data_i[398] & sel_one_hot_i[3];
  assign data_masked[397] = data_i[397] & sel_one_hot_i[3];
  assign data_masked[396] = data_i[396] & sel_one_hot_i[3];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[3];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[3];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[3];
  assign data_o[0] = N1 | data_masked[0];
  assign N1 = N0 | data_masked[131];
  assign N0 = data_masked[393] | data_masked[262];
  assign data_o[1] = N3 | data_masked[1];
  assign N3 = N2 | data_masked[132];
  assign N2 = data_masked[394] | data_masked[263];
  assign data_o[2] = N5 | data_masked[2];
  assign N5 = N4 | data_masked[133];
  assign N4 = data_masked[395] | data_masked[264];
  assign data_o[3] = N7 | data_masked[3];
  assign N7 = N6 | data_masked[134];
  assign N6 = data_masked[396] | data_masked[265];
  assign data_o[4] = N9 | data_masked[4];
  assign N9 = N8 | data_masked[135];
  assign N8 = data_masked[397] | data_masked[266];
  assign data_o[5] = N11 | data_masked[5];
  assign N11 = N10 | data_masked[136];
  assign N10 = data_masked[398] | data_masked[267];
  assign data_o[6] = N13 | data_masked[6];
  assign N13 = N12 | data_masked[137];
  assign N12 = data_masked[399] | data_masked[268];
  assign data_o[7] = N15 | data_masked[7];
  assign N15 = N14 | data_masked[138];
  assign N14 = data_masked[400] | data_masked[269];
  assign data_o[8] = N17 | data_masked[8];
  assign N17 = N16 | data_masked[139];
  assign N16 = data_masked[401] | data_masked[270];
  assign data_o[9] = N19 | data_masked[9];
  assign N19 = N18 | data_masked[140];
  assign N18 = data_masked[402] | data_masked[271];
  assign data_o[10] = N21 | data_masked[10];
  assign N21 = N20 | data_masked[141];
  assign N20 = data_masked[403] | data_masked[272];
  assign data_o[11] = N23 | data_masked[11];
  assign N23 = N22 | data_masked[142];
  assign N22 = data_masked[404] | data_masked[273];
  assign data_o[12] = N25 | data_masked[12];
  assign N25 = N24 | data_masked[143];
  assign N24 = data_masked[405] | data_masked[274];
  assign data_o[13] = N27 | data_masked[13];
  assign N27 = N26 | data_masked[144];
  assign N26 = data_masked[406] | data_masked[275];
  assign data_o[14] = N29 | data_masked[14];
  assign N29 = N28 | data_masked[145];
  assign N28 = data_masked[407] | data_masked[276];
  assign data_o[15] = N31 | data_masked[15];
  assign N31 = N30 | data_masked[146];
  assign N30 = data_masked[408] | data_masked[277];
  assign data_o[16] = N33 | data_masked[16];
  assign N33 = N32 | data_masked[147];
  assign N32 = data_masked[409] | data_masked[278];
  assign data_o[17] = N35 | data_masked[17];
  assign N35 = N34 | data_masked[148];
  assign N34 = data_masked[410] | data_masked[279];
  assign data_o[18] = N37 | data_masked[18];
  assign N37 = N36 | data_masked[149];
  assign N36 = data_masked[411] | data_masked[280];
  assign data_o[19] = N39 | data_masked[19];
  assign N39 = N38 | data_masked[150];
  assign N38 = data_masked[412] | data_masked[281];
  assign data_o[20] = N41 | data_masked[20];
  assign N41 = N40 | data_masked[151];
  assign N40 = data_masked[413] | data_masked[282];
  assign data_o[21] = N43 | data_masked[21];
  assign N43 = N42 | data_masked[152];
  assign N42 = data_masked[414] | data_masked[283];
  assign data_o[22] = N45 | data_masked[22];
  assign N45 = N44 | data_masked[153];
  assign N44 = data_masked[415] | data_masked[284];
  assign data_o[23] = N47 | data_masked[23];
  assign N47 = N46 | data_masked[154];
  assign N46 = data_masked[416] | data_masked[285];
  assign data_o[24] = N49 | data_masked[24];
  assign N49 = N48 | data_masked[155];
  assign N48 = data_masked[417] | data_masked[286];
  assign data_o[25] = N51 | data_masked[25];
  assign N51 = N50 | data_masked[156];
  assign N50 = data_masked[418] | data_masked[287];
  assign data_o[26] = N53 | data_masked[26];
  assign N53 = N52 | data_masked[157];
  assign N52 = data_masked[419] | data_masked[288];
  assign data_o[27] = N55 | data_masked[27];
  assign N55 = N54 | data_masked[158];
  assign N54 = data_masked[420] | data_masked[289];
  assign data_o[28] = N57 | data_masked[28];
  assign N57 = N56 | data_masked[159];
  assign N56 = data_masked[421] | data_masked[290];
  assign data_o[29] = N59 | data_masked[29];
  assign N59 = N58 | data_masked[160];
  assign N58 = data_masked[422] | data_masked[291];
  assign data_o[30] = N61 | data_masked[30];
  assign N61 = N60 | data_masked[161];
  assign N60 = data_masked[423] | data_masked[292];
  assign data_o[31] = N63 | data_masked[31];
  assign N63 = N62 | data_masked[162];
  assign N62 = data_masked[424] | data_masked[293];
  assign data_o[32] = N65 | data_masked[32];
  assign N65 = N64 | data_masked[163];
  assign N64 = data_masked[425] | data_masked[294];
  assign data_o[33] = N67 | data_masked[33];
  assign N67 = N66 | data_masked[164];
  assign N66 = data_masked[426] | data_masked[295];
  assign data_o[34] = N69 | data_masked[34];
  assign N69 = N68 | data_masked[165];
  assign N68 = data_masked[427] | data_masked[296];
  assign data_o[35] = N71 | data_masked[35];
  assign N71 = N70 | data_masked[166];
  assign N70 = data_masked[428] | data_masked[297];
  assign data_o[36] = N73 | data_masked[36];
  assign N73 = N72 | data_masked[167];
  assign N72 = data_masked[429] | data_masked[298];
  assign data_o[37] = N75 | data_masked[37];
  assign N75 = N74 | data_masked[168];
  assign N74 = data_masked[430] | data_masked[299];
  assign data_o[38] = N77 | data_masked[38];
  assign N77 = N76 | data_masked[169];
  assign N76 = data_masked[431] | data_masked[300];
  assign data_o[39] = N79 | data_masked[39];
  assign N79 = N78 | data_masked[170];
  assign N78 = data_masked[432] | data_masked[301];
  assign data_o[40] = N81 | data_masked[40];
  assign N81 = N80 | data_masked[171];
  assign N80 = data_masked[433] | data_masked[302];
  assign data_o[41] = N83 | data_masked[41];
  assign N83 = N82 | data_masked[172];
  assign N82 = data_masked[434] | data_masked[303];
  assign data_o[42] = N85 | data_masked[42];
  assign N85 = N84 | data_masked[173];
  assign N84 = data_masked[435] | data_masked[304];
  assign data_o[43] = N87 | data_masked[43];
  assign N87 = N86 | data_masked[174];
  assign N86 = data_masked[436] | data_masked[305];
  assign data_o[44] = N89 | data_masked[44];
  assign N89 = N88 | data_masked[175];
  assign N88 = data_masked[437] | data_masked[306];
  assign data_o[45] = N91 | data_masked[45];
  assign N91 = N90 | data_masked[176];
  assign N90 = data_masked[438] | data_masked[307];
  assign data_o[46] = N93 | data_masked[46];
  assign N93 = N92 | data_masked[177];
  assign N92 = data_masked[439] | data_masked[308];
  assign data_o[47] = N95 | data_masked[47];
  assign N95 = N94 | data_masked[178];
  assign N94 = data_masked[440] | data_masked[309];
  assign data_o[48] = N97 | data_masked[48];
  assign N97 = N96 | data_masked[179];
  assign N96 = data_masked[441] | data_masked[310];
  assign data_o[49] = N99 | data_masked[49];
  assign N99 = N98 | data_masked[180];
  assign N98 = data_masked[442] | data_masked[311];
  assign data_o[50] = N101 | data_masked[50];
  assign N101 = N100 | data_masked[181];
  assign N100 = data_masked[443] | data_masked[312];
  assign data_o[51] = N103 | data_masked[51];
  assign N103 = N102 | data_masked[182];
  assign N102 = data_masked[444] | data_masked[313];
  assign data_o[52] = N105 | data_masked[52];
  assign N105 = N104 | data_masked[183];
  assign N104 = data_masked[445] | data_masked[314];
  assign data_o[53] = N107 | data_masked[53];
  assign N107 = N106 | data_masked[184];
  assign N106 = data_masked[446] | data_masked[315];
  assign data_o[54] = N109 | data_masked[54];
  assign N109 = N108 | data_masked[185];
  assign N108 = data_masked[447] | data_masked[316];
  assign data_o[55] = N111 | data_masked[55];
  assign N111 = N110 | data_masked[186];
  assign N110 = data_masked[448] | data_masked[317];
  assign data_o[56] = N113 | data_masked[56];
  assign N113 = N112 | data_masked[187];
  assign N112 = data_masked[449] | data_masked[318];
  assign data_o[57] = N115 | data_masked[57];
  assign N115 = N114 | data_masked[188];
  assign N114 = data_masked[450] | data_masked[319];
  assign data_o[58] = N117 | data_masked[58];
  assign N117 = N116 | data_masked[189];
  assign N116 = data_masked[451] | data_masked[320];
  assign data_o[59] = N119 | data_masked[59];
  assign N119 = N118 | data_masked[190];
  assign N118 = data_masked[452] | data_masked[321];
  assign data_o[60] = N121 | data_masked[60];
  assign N121 = N120 | data_masked[191];
  assign N120 = data_masked[453] | data_masked[322];
  assign data_o[61] = N123 | data_masked[61];
  assign N123 = N122 | data_masked[192];
  assign N122 = data_masked[454] | data_masked[323];
  assign data_o[62] = N125 | data_masked[62];
  assign N125 = N124 | data_masked[193];
  assign N124 = data_masked[455] | data_masked[324];
  assign data_o[63] = N127 | data_masked[63];
  assign N127 = N126 | data_masked[194];
  assign N126 = data_masked[456] | data_masked[325];
  assign data_o[64] = N129 | data_masked[64];
  assign N129 = N128 | data_masked[195];
  assign N128 = data_masked[457] | data_masked[326];
  assign data_o[65] = N131 | data_masked[65];
  assign N131 = N130 | data_masked[196];
  assign N130 = data_masked[458] | data_masked[327];
  assign data_o[66] = N133 | data_masked[66];
  assign N133 = N132 | data_masked[197];
  assign N132 = data_masked[459] | data_masked[328];
  assign data_o[67] = N135 | data_masked[67];
  assign N135 = N134 | data_masked[198];
  assign N134 = data_masked[460] | data_masked[329];
  assign data_o[68] = N137 | data_masked[68];
  assign N137 = N136 | data_masked[199];
  assign N136 = data_masked[461] | data_masked[330];
  assign data_o[69] = N139 | data_masked[69];
  assign N139 = N138 | data_masked[200];
  assign N138 = data_masked[462] | data_masked[331];
  assign data_o[70] = N141 | data_masked[70];
  assign N141 = N140 | data_masked[201];
  assign N140 = data_masked[463] | data_masked[332];
  assign data_o[71] = N143 | data_masked[71];
  assign N143 = N142 | data_masked[202];
  assign N142 = data_masked[464] | data_masked[333];
  assign data_o[72] = N145 | data_masked[72];
  assign N145 = N144 | data_masked[203];
  assign N144 = data_masked[465] | data_masked[334];
  assign data_o[73] = N147 | data_masked[73];
  assign N147 = N146 | data_masked[204];
  assign N146 = data_masked[466] | data_masked[335];
  assign data_o[74] = N149 | data_masked[74];
  assign N149 = N148 | data_masked[205];
  assign N148 = data_masked[467] | data_masked[336];
  assign data_o[75] = N151 | data_masked[75];
  assign N151 = N150 | data_masked[206];
  assign N150 = data_masked[468] | data_masked[337];
  assign data_o[76] = N153 | data_masked[76];
  assign N153 = N152 | data_masked[207];
  assign N152 = data_masked[469] | data_masked[338];
  assign data_o[77] = N155 | data_masked[77];
  assign N155 = N154 | data_masked[208];
  assign N154 = data_masked[470] | data_masked[339];
  assign data_o[78] = N157 | data_masked[78];
  assign N157 = N156 | data_masked[209];
  assign N156 = data_masked[471] | data_masked[340];
  assign data_o[79] = N159 | data_masked[79];
  assign N159 = N158 | data_masked[210];
  assign N158 = data_masked[472] | data_masked[341];
  assign data_o[80] = N161 | data_masked[80];
  assign N161 = N160 | data_masked[211];
  assign N160 = data_masked[473] | data_masked[342];
  assign data_o[81] = N163 | data_masked[81];
  assign N163 = N162 | data_masked[212];
  assign N162 = data_masked[474] | data_masked[343];
  assign data_o[82] = N165 | data_masked[82];
  assign N165 = N164 | data_masked[213];
  assign N164 = data_masked[475] | data_masked[344];
  assign data_o[83] = N167 | data_masked[83];
  assign N167 = N166 | data_masked[214];
  assign N166 = data_masked[476] | data_masked[345];
  assign data_o[84] = N169 | data_masked[84];
  assign N169 = N168 | data_masked[215];
  assign N168 = data_masked[477] | data_masked[346];
  assign data_o[85] = N171 | data_masked[85];
  assign N171 = N170 | data_masked[216];
  assign N170 = data_masked[478] | data_masked[347];
  assign data_o[86] = N173 | data_masked[86];
  assign N173 = N172 | data_masked[217];
  assign N172 = data_masked[479] | data_masked[348];
  assign data_o[87] = N175 | data_masked[87];
  assign N175 = N174 | data_masked[218];
  assign N174 = data_masked[480] | data_masked[349];
  assign data_o[88] = N177 | data_masked[88];
  assign N177 = N176 | data_masked[219];
  assign N176 = data_masked[481] | data_masked[350];
  assign data_o[89] = N179 | data_masked[89];
  assign N179 = N178 | data_masked[220];
  assign N178 = data_masked[482] | data_masked[351];
  assign data_o[90] = N181 | data_masked[90];
  assign N181 = N180 | data_masked[221];
  assign N180 = data_masked[483] | data_masked[352];
  assign data_o[91] = N183 | data_masked[91];
  assign N183 = N182 | data_masked[222];
  assign N182 = data_masked[484] | data_masked[353];
  assign data_o[92] = N185 | data_masked[92];
  assign N185 = N184 | data_masked[223];
  assign N184 = data_masked[485] | data_masked[354];
  assign data_o[93] = N187 | data_masked[93];
  assign N187 = N186 | data_masked[224];
  assign N186 = data_masked[486] | data_masked[355];
  assign data_o[94] = N189 | data_masked[94];
  assign N189 = N188 | data_masked[225];
  assign N188 = data_masked[487] | data_masked[356];
  assign data_o[95] = N191 | data_masked[95];
  assign N191 = N190 | data_masked[226];
  assign N190 = data_masked[488] | data_masked[357];
  assign data_o[96] = N193 | data_masked[96];
  assign N193 = N192 | data_masked[227];
  assign N192 = data_masked[489] | data_masked[358];
  assign data_o[97] = N195 | data_masked[97];
  assign N195 = N194 | data_masked[228];
  assign N194 = data_masked[490] | data_masked[359];
  assign data_o[98] = N197 | data_masked[98];
  assign N197 = N196 | data_masked[229];
  assign N196 = data_masked[491] | data_masked[360];
  assign data_o[99] = N199 | data_masked[99];
  assign N199 = N198 | data_masked[230];
  assign N198 = data_masked[492] | data_masked[361];
  assign data_o[100] = N201 | data_masked[100];
  assign N201 = N200 | data_masked[231];
  assign N200 = data_masked[493] | data_masked[362];
  assign data_o[101] = N203 | data_masked[101];
  assign N203 = N202 | data_masked[232];
  assign N202 = data_masked[494] | data_masked[363];
  assign data_o[102] = N205 | data_masked[102];
  assign N205 = N204 | data_masked[233];
  assign N204 = data_masked[495] | data_masked[364];
  assign data_o[103] = N207 | data_masked[103];
  assign N207 = N206 | data_masked[234];
  assign N206 = data_masked[496] | data_masked[365];
  assign data_o[104] = N209 | data_masked[104];
  assign N209 = N208 | data_masked[235];
  assign N208 = data_masked[497] | data_masked[366];
  assign data_o[105] = N211 | data_masked[105];
  assign N211 = N210 | data_masked[236];
  assign N210 = data_masked[498] | data_masked[367];
  assign data_o[106] = N213 | data_masked[106];
  assign N213 = N212 | data_masked[237];
  assign N212 = data_masked[499] | data_masked[368];
  assign data_o[107] = N215 | data_masked[107];
  assign N215 = N214 | data_masked[238];
  assign N214 = data_masked[500] | data_masked[369];
  assign data_o[108] = N217 | data_masked[108];
  assign N217 = N216 | data_masked[239];
  assign N216 = data_masked[501] | data_masked[370];
  assign data_o[109] = N219 | data_masked[109];
  assign N219 = N218 | data_masked[240];
  assign N218 = data_masked[502] | data_masked[371];
  assign data_o[110] = N221 | data_masked[110];
  assign N221 = N220 | data_masked[241];
  assign N220 = data_masked[503] | data_masked[372];
  assign data_o[111] = N223 | data_masked[111];
  assign N223 = N222 | data_masked[242];
  assign N222 = data_masked[504] | data_masked[373];
  assign data_o[112] = N225 | data_masked[112];
  assign N225 = N224 | data_masked[243];
  assign N224 = data_masked[505] | data_masked[374];
  assign data_o[113] = N227 | data_masked[113];
  assign N227 = N226 | data_masked[244];
  assign N226 = data_masked[506] | data_masked[375];
  assign data_o[114] = N229 | data_masked[114];
  assign N229 = N228 | data_masked[245];
  assign N228 = data_masked[507] | data_masked[376];
  assign data_o[115] = N231 | data_masked[115];
  assign N231 = N230 | data_masked[246];
  assign N230 = data_masked[508] | data_masked[377];
  assign data_o[116] = N233 | data_masked[116];
  assign N233 = N232 | data_masked[247];
  assign N232 = data_masked[509] | data_masked[378];
  assign data_o[117] = N235 | data_masked[117];
  assign N235 = N234 | data_masked[248];
  assign N234 = data_masked[510] | data_masked[379];
  assign data_o[118] = N237 | data_masked[118];
  assign N237 = N236 | data_masked[249];
  assign N236 = data_masked[511] | data_masked[380];
  assign data_o[119] = N239 | data_masked[119];
  assign N239 = N238 | data_masked[250];
  assign N238 = data_masked[512] | data_masked[381];
  assign data_o[120] = N241 | data_masked[120];
  assign N241 = N240 | data_masked[251];
  assign N240 = data_masked[513] | data_masked[382];
  assign data_o[121] = N243 | data_masked[121];
  assign N243 = N242 | data_masked[252];
  assign N242 = data_masked[514] | data_masked[383];
  assign data_o[122] = N245 | data_masked[122];
  assign N245 = N244 | data_masked[253];
  assign N244 = data_masked[515] | data_masked[384];
  assign data_o[123] = N247 | data_masked[123];
  assign N247 = N246 | data_masked[254];
  assign N246 = data_masked[516] | data_masked[385];
  assign data_o[124] = N249 | data_masked[124];
  assign N249 = N248 | data_masked[255];
  assign N248 = data_masked[517] | data_masked[386];
  assign data_o[125] = N251 | data_masked[125];
  assign N251 = N250 | data_masked[256];
  assign N250 = data_masked[518] | data_masked[387];
  assign data_o[126] = N253 | data_masked[126];
  assign N253 = N252 | data_masked[257];
  assign N252 = data_masked[519] | data_masked[388];
  assign data_o[127] = N255 | data_masked[127];
  assign N255 = N254 | data_masked[258];
  assign N254 = data_masked[520] | data_masked[389];
  assign data_o[128] = N257 | data_masked[128];
  assign N257 = N256 | data_masked[259];
  assign N256 = data_masked[521] | data_masked[390];
  assign data_o[129] = N259 | data_masked[129];
  assign N259 = N258 | data_masked[260];
  assign N258 = data_masked[522] | data_masked[391];
  assign data_o[130] = N261 | data_masked[130];
  assign N261 = N260 | data_masked[261];
  assign N260 = data_masked[523] | data_masked[392];

endmodule



module bsg_mux_one_hot_width_p131_els_p5
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [654:0] data_i;
  input [4:0] sel_one_hot_i;
  output [130:0] data_o;
  wire [130:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392;
  wire [654:0] data_masked;
  assign data_masked[130] = data_i[130] & sel_one_hot_i[0];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[0];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[0];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[0];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[0];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[0];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[0];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[0];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[0];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[0];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[0];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[0];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[0];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[0];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[0];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[0];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[0];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[0];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[0];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[0];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[0];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[0];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[0];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[0];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[0];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[0];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[0];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[0];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[0];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[0];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[0];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[0];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[0];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[0];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[0];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[0];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[0];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[0];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[0];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[0];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[0];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[0];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[0];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[0];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[0];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[0];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[0];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[0];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[0];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[0];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[0];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[0];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[0];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[0];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[0];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[0];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[0];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[0];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[0];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[0];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[0];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[0];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[0];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[1];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[1];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[1];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[1];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[1];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[1];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[1];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[1];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[1];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[1];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[1];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[1];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[1];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[1];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[1];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[1];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[1];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[1];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[1];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[1];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[1];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[1];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[1];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[1];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[1];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[1];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[1];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[1];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[1];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[1];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[1];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[1];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[1];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[1];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[1];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[1];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[1];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[1];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[1];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[1];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[1];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[1];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[1];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[1];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[1];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[1];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[1];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[1];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[1];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[1];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[1];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[1];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[1];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[1];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[1];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[1];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[1];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[1];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[1];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[1];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[1];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[1];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[1];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[1];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[1];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[1];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[1];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[1];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[1];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[1];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[1];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[1];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[1];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[1];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[1];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[1];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[1];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[1];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[1];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[1];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[1];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[1];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[1];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[1];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[1];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[1];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[1];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[1];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[1];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[1];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[1];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[1];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[1];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[1];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[1];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[1];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[1];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[1];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[1];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[1];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[1];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[1];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[1];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[1];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[1];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[1];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[1];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[1];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[1];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[1];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[1];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[1];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[1];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[1];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[1];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[1];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[1];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[1];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[1];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[1];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[1];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[1];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[1];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[1];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[1];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[1];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[1];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[1];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[1];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[1];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[2];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[2];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[2];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[2];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[2];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[2];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[2];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[2];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[2];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[2];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[2];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[2];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[2];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[2];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[2];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[2];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[2];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[2];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[2];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[2];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[2];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[2];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[2];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[2];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[2];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[2];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[2];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[2];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[2];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[2];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[2];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[2];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[2];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[2];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[2];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[2];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[2];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[2];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[2];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[2];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[2];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[2];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[2];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[2];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[2];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[2];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[2];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[2];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[2];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[2];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[2];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[2];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[2];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[2];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[2];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[2];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[2];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[2];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[2];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[2];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[2];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[2];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[2];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[2];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[2];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[2];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[2];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[2];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[2];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[2];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[2];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[2];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[2];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[2];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[2];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[2];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[2];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[2];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[2];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[2];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[2];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[2];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[2];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[2];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[2];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[2];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[2];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[2];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[2];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[2];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[2];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[2];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[2];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[2];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[2];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[2];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[2];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[2];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[2];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[2];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[2];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[2];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[2];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[2];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[2];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[2];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[2];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[2];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[2];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[2];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[2];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[2];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[2];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[2];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[2];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[2];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[2];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[2];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[2];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[2];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[2];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[2];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[2];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[2];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[2];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[2];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[2];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[2];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[2];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[2];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[2];
  assign data_masked[523] = data_i[523] & sel_one_hot_i[3];
  assign data_masked[522] = data_i[522] & sel_one_hot_i[3];
  assign data_masked[521] = data_i[521] & sel_one_hot_i[3];
  assign data_masked[520] = data_i[520] & sel_one_hot_i[3];
  assign data_masked[519] = data_i[519] & sel_one_hot_i[3];
  assign data_masked[518] = data_i[518] & sel_one_hot_i[3];
  assign data_masked[517] = data_i[517] & sel_one_hot_i[3];
  assign data_masked[516] = data_i[516] & sel_one_hot_i[3];
  assign data_masked[515] = data_i[515] & sel_one_hot_i[3];
  assign data_masked[514] = data_i[514] & sel_one_hot_i[3];
  assign data_masked[513] = data_i[513] & sel_one_hot_i[3];
  assign data_masked[512] = data_i[512] & sel_one_hot_i[3];
  assign data_masked[511] = data_i[511] & sel_one_hot_i[3];
  assign data_masked[510] = data_i[510] & sel_one_hot_i[3];
  assign data_masked[509] = data_i[509] & sel_one_hot_i[3];
  assign data_masked[508] = data_i[508] & sel_one_hot_i[3];
  assign data_masked[507] = data_i[507] & sel_one_hot_i[3];
  assign data_masked[506] = data_i[506] & sel_one_hot_i[3];
  assign data_masked[505] = data_i[505] & sel_one_hot_i[3];
  assign data_masked[504] = data_i[504] & sel_one_hot_i[3];
  assign data_masked[503] = data_i[503] & sel_one_hot_i[3];
  assign data_masked[502] = data_i[502] & sel_one_hot_i[3];
  assign data_masked[501] = data_i[501] & sel_one_hot_i[3];
  assign data_masked[500] = data_i[500] & sel_one_hot_i[3];
  assign data_masked[499] = data_i[499] & sel_one_hot_i[3];
  assign data_masked[498] = data_i[498] & sel_one_hot_i[3];
  assign data_masked[497] = data_i[497] & sel_one_hot_i[3];
  assign data_masked[496] = data_i[496] & sel_one_hot_i[3];
  assign data_masked[495] = data_i[495] & sel_one_hot_i[3];
  assign data_masked[494] = data_i[494] & sel_one_hot_i[3];
  assign data_masked[493] = data_i[493] & sel_one_hot_i[3];
  assign data_masked[492] = data_i[492] & sel_one_hot_i[3];
  assign data_masked[491] = data_i[491] & sel_one_hot_i[3];
  assign data_masked[490] = data_i[490] & sel_one_hot_i[3];
  assign data_masked[489] = data_i[489] & sel_one_hot_i[3];
  assign data_masked[488] = data_i[488] & sel_one_hot_i[3];
  assign data_masked[487] = data_i[487] & sel_one_hot_i[3];
  assign data_masked[486] = data_i[486] & sel_one_hot_i[3];
  assign data_masked[485] = data_i[485] & sel_one_hot_i[3];
  assign data_masked[484] = data_i[484] & sel_one_hot_i[3];
  assign data_masked[483] = data_i[483] & sel_one_hot_i[3];
  assign data_masked[482] = data_i[482] & sel_one_hot_i[3];
  assign data_masked[481] = data_i[481] & sel_one_hot_i[3];
  assign data_masked[480] = data_i[480] & sel_one_hot_i[3];
  assign data_masked[479] = data_i[479] & sel_one_hot_i[3];
  assign data_masked[478] = data_i[478] & sel_one_hot_i[3];
  assign data_masked[477] = data_i[477] & sel_one_hot_i[3];
  assign data_masked[476] = data_i[476] & sel_one_hot_i[3];
  assign data_masked[475] = data_i[475] & sel_one_hot_i[3];
  assign data_masked[474] = data_i[474] & sel_one_hot_i[3];
  assign data_masked[473] = data_i[473] & sel_one_hot_i[3];
  assign data_masked[472] = data_i[472] & sel_one_hot_i[3];
  assign data_masked[471] = data_i[471] & sel_one_hot_i[3];
  assign data_masked[470] = data_i[470] & sel_one_hot_i[3];
  assign data_masked[469] = data_i[469] & sel_one_hot_i[3];
  assign data_masked[468] = data_i[468] & sel_one_hot_i[3];
  assign data_masked[467] = data_i[467] & sel_one_hot_i[3];
  assign data_masked[466] = data_i[466] & sel_one_hot_i[3];
  assign data_masked[465] = data_i[465] & sel_one_hot_i[3];
  assign data_masked[464] = data_i[464] & sel_one_hot_i[3];
  assign data_masked[463] = data_i[463] & sel_one_hot_i[3];
  assign data_masked[462] = data_i[462] & sel_one_hot_i[3];
  assign data_masked[461] = data_i[461] & sel_one_hot_i[3];
  assign data_masked[460] = data_i[460] & sel_one_hot_i[3];
  assign data_masked[459] = data_i[459] & sel_one_hot_i[3];
  assign data_masked[458] = data_i[458] & sel_one_hot_i[3];
  assign data_masked[457] = data_i[457] & sel_one_hot_i[3];
  assign data_masked[456] = data_i[456] & sel_one_hot_i[3];
  assign data_masked[455] = data_i[455] & sel_one_hot_i[3];
  assign data_masked[454] = data_i[454] & sel_one_hot_i[3];
  assign data_masked[453] = data_i[453] & sel_one_hot_i[3];
  assign data_masked[452] = data_i[452] & sel_one_hot_i[3];
  assign data_masked[451] = data_i[451] & sel_one_hot_i[3];
  assign data_masked[450] = data_i[450] & sel_one_hot_i[3];
  assign data_masked[449] = data_i[449] & sel_one_hot_i[3];
  assign data_masked[448] = data_i[448] & sel_one_hot_i[3];
  assign data_masked[447] = data_i[447] & sel_one_hot_i[3];
  assign data_masked[446] = data_i[446] & sel_one_hot_i[3];
  assign data_masked[445] = data_i[445] & sel_one_hot_i[3];
  assign data_masked[444] = data_i[444] & sel_one_hot_i[3];
  assign data_masked[443] = data_i[443] & sel_one_hot_i[3];
  assign data_masked[442] = data_i[442] & sel_one_hot_i[3];
  assign data_masked[441] = data_i[441] & sel_one_hot_i[3];
  assign data_masked[440] = data_i[440] & sel_one_hot_i[3];
  assign data_masked[439] = data_i[439] & sel_one_hot_i[3];
  assign data_masked[438] = data_i[438] & sel_one_hot_i[3];
  assign data_masked[437] = data_i[437] & sel_one_hot_i[3];
  assign data_masked[436] = data_i[436] & sel_one_hot_i[3];
  assign data_masked[435] = data_i[435] & sel_one_hot_i[3];
  assign data_masked[434] = data_i[434] & sel_one_hot_i[3];
  assign data_masked[433] = data_i[433] & sel_one_hot_i[3];
  assign data_masked[432] = data_i[432] & sel_one_hot_i[3];
  assign data_masked[431] = data_i[431] & sel_one_hot_i[3];
  assign data_masked[430] = data_i[430] & sel_one_hot_i[3];
  assign data_masked[429] = data_i[429] & sel_one_hot_i[3];
  assign data_masked[428] = data_i[428] & sel_one_hot_i[3];
  assign data_masked[427] = data_i[427] & sel_one_hot_i[3];
  assign data_masked[426] = data_i[426] & sel_one_hot_i[3];
  assign data_masked[425] = data_i[425] & sel_one_hot_i[3];
  assign data_masked[424] = data_i[424] & sel_one_hot_i[3];
  assign data_masked[423] = data_i[423] & sel_one_hot_i[3];
  assign data_masked[422] = data_i[422] & sel_one_hot_i[3];
  assign data_masked[421] = data_i[421] & sel_one_hot_i[3];
  assign data_masked[420] = data_i[420] & sel_one_hot_i[3];
  assign data_masked[419] = data_i[419] & sel_one_hot_i[3];
  assign data_masked[418] = data_i[418] & sel_one_hot_i[3];
  assign data_masked[417] = data_i[417] & sel_one_hot_i[3];
  assign data_masked[416] = data_i[416] & sel_one_hot_i[3];
  assign data_masked[415] = data_i[415] & sel_one_hot_i[3];
  assign data_masked[414] = data_i[414] & sel_one_hot_i[3];
  assign data_masked[413] = data_i[413] & sel_one_hot_i[3];
  assign data_masked[412] = data_i[412] & sel_one_hot_i[3];
  assign data_masked[411] = data_i[411] & sel_one_hot_i[3];
  assign data_masked[410] = data_i[410] & sel_one_hot_i[3];
  assign data_masked[409] = data_i[409] & sel_one_hot_i[3];
  assign data_masked[408] = data_i[408] & sel_one_hot_i[3];
  assign data_masked[407] = data_i[407] & sel_one_hot_i[3];
  assign data_masked[406] = data_i[406] & sel_one_hot_i[3];
  assign data_masked[405] = data_i[405] & sel_one_hot_i[3];
  assign data_masked[404] = data_i[404] & sel_one_hot_i[3];
  assign data_masked[403] = data_i[403] & sel_one_hot_i[3];
  assign data_masked[402] = data_i[402] & sel_one_hot_i[3];
  assign data_masked[401] = data_i[401] & sel_one_hot_i[3];
  assign data_masked[400] = data_i[400] & sel_one_hot_i[3];
  assign data_masked[399] = data_i[399] & sel_one_hot_i[3];
  assign data_masked[398] = data_i[398] & sel_one_hot_i[3];
  assign data_masked[397] = data_i[397] & sel_one_hot_i[3];
  assign data_masked[396] = data_i[396] & sel_one_hot_i[3];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[3];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[3];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[3];
  assign data_masked[654] = data_i[654] & sel_one_hot_i[4];
  assign data_masked[653] = data_i[653] & sel_one_hot_i[4];
  assign data_masked[652] = data_i[652] & sel_one_hot_i[4];
  assign data_masked[651] = data_i[651] & sel_one_hot_i[4];
  assign data_masked[650] = data_i[650] & sel_one_hot_i[4];
  assign data_masked[649] = data_i[649] & sel_one_hot_i[4];
  assign data_masked[648] = data_i[648] & sel_one_hot_i[4];
  assign data_masked[647] = data_i[647] & sel_one_hot_i[4];
  assign data_masked[646] = data_i[646] & sel_one_hot_i[4];
  assign data_masked[645] = data_i[645] & sel_one_hot_i[4];
  assign data_masked[644] = data_i[644] & sel_one_hot_i[4];
  assign data_masked[643] = data_i[643] & sel_one_hot_i[4];
  assign data_masked[642] = data_i[642] & sel_one_hot_i[4];
  assign data_masked[641] = data_i[641] & sel_one_hot_i[4];
  assign data_masked[640] = data_i[640] & sel_one_hot_i[4];
  assign data_masked[639] = data_i[639] & sel_one_hot_i[4];
  assign data_masked[638] = data_i[638] & sel_one_hot_i[4];
  assign data_masked[637] = data_i[637] & sel_one_hot_i[4];
  assign data_masked[636] = data_i[636] & sel_one_hot_i[4];
  assign data_masked[635] = data_i[635] & sel_one_hot_i[4];
  assign data_masked[634] = data_i[634] & sel_one_hot_i[4];
  assign data_masked[633] = data_i[633] & sel_one_hot_i[4];
  assign data_masked[632] = data_i[632] & sel_one_hot_i[4];
  assign data_masked[631] = data_i[631] & sel_one_hot_i[4];
  assign data_masked[630] = data_i[630] & sel_one_hot_i[4];
  assign data_masked[629] = data_i[629] & sel_one_hot_i[4];
  assign data_masked[628] = data_i[628] & sel_one_hot_i[4];
  assign data_masked[627] = data_i[627] & sel_one_hot_i[4];
  assign data_masked[626] = data_i[626] & sel_one_hot_i[4];
  assign data_masked[625] = data_i[625] & sel_one_hot_i[4];
  assign data_masked[624] = data_i[624] & sel_one_hot_i[4];
  assign data_masked[623] = data_i[623] & sel_one_hot_i[4];
  assign data_masked[622] = data_i[622] & sel_one_hot_i[4];
  assign data_masked[621] = data_i[621] & sel_one_hot_i[4];
  assign data_masked[620] = data_i[620] & sel_one_hot_i[4];
  assign data_masked[619] = data_i[619] & sel_one_hot_i[4];
  assign data_masked[618] = data_i[618] & sel_one_hot_i[4];
  assign data_masked[617] = data_i[617] & sel_one_hot_i[4];
  assign data_masked[616] = data_i[616] & sel_one_hot_i[4];
  assign data_masked[615] = data_i[615] & sel_one_hot_i[4];
  assign data_masked[614] = data_i[614] & sel_one_hot_i[4];
  assign data_masked[613] = data_i[613] & sel_one_hot_i[4];
  assign data_masked[612] = data_i[612] & sel_one_hot_i[4];
  assign data_masked[611] = data_i[611] & sel_one_hot_i[4];
  assign data_masked[610] = data_i[610] & sel_one_hot_i[4];
  assign data_masked[609] = data_i[609] & sel_one_hot_i[4];
  assign data_masked[608] = data_i[608] & sel_one_hot_i[4];
  assign data_masked[607] = data_i[607] & sel_one_hot_i[4];
  assign data_masked[606] = data_i[606] & sel_one_hot_i[4];
  assign data_masked[605] = data_i[605] & sel_one_hot_i[4];
  assign data_masked[604] = data_i[604] & sel_one_hot_i[4];
  assign data_masked[603] = data_i[603] & sel_one_hot_i[4];
  assign data_masked[602] = data_i[602] & sel_one_hot_i[4];
  assign data_masked[601] = data_i[601] & sel_one_hot_i[4];
  assign data_masked[600] = data_i[600] & sel_one_hot_i[4];
  assign data_masked[599] = data_i[599] & sel_one_hot_i[4];
  assign data_masked[598] = data_i[598] & sel_one_hot_i[4];
  assign data_masked[597] = data_i[597] & sel_one_hot_i[4];
  assign data_masked[596] = data_i[596] & sel_one_hot_i[4];
  assign data_masked[595] = data_i[595] & sel_one_hot_i[4];
  assign data_masked[594] = data_i[594] & sel_one_hot_i[4];
  assign data_masked[593] = data_i[593] & sel_one_hot_i[4];
  assign data_masked[592] = data_i[592] & sel_one_hot_i[4];
  assign data_masked[591] = data_i[591] & sel_one_hot_i[4];
  assign data_masked[590] = data_i[590] & sel_one_hot_i[4];
  assign data_masked[589] = data_i[589] & sel_one_hot_i[4];
  assign data_masked[588] = data_i[588] & sel_one_hot_i[4];
  assign data_masked[587] = data_i[587] & sel_one_hot_i[4];
  assign data_masked[586] = data_i[586] & sel_one_hot_i[4];
  assign data_masked[585] = data_i[585] & sel_one_hot_i[4];
  assign data_masked[584] = data_i[584] & sel_one_hot_i[4];
  assign data_masked[583] = data_i[583] & sel_one_hot_i[4];
  assign data_masked[582] = data_i[582] & sel_one_hot_i[4];
  assign data_masked[581] = data_i[581] & sel_one_hot_i[4];
  assign data_masked[580] = data_i[580] & sel_one_hot_i[4];
  assign data_masked[579] = data_i[579] & sel_one_hot_i[4];
  assign data_masked[578] = data_i[578] & sel_one_hot_i[4];
  assign data_masked[577] = data_i[577] & sel_one_hot_i[4];
  assign data_masked[576] = data_i[576] & sel_one_hot_i[4];
  assign data_masked[575] = data_i[575] & sel_one_hot_i[4];
  assign data_masked[574] = data_i[574] & sel_one_hot_i[4];
  assign data_masked[573] = data_i[573] & sel_one_hot_i[4];
  assign data_masked[572] = data_i[572] & sel_one_hot_i[4];
  assign data_masked[571] = data_i[571] & sel_one_hot_i[4];
  assign data_masked[570] = data_i[570] & sel_one_hot_i[4];
  assign data_masked[569] = data_i[569] & sel_one_hot_i[4];
  assign data_masked[568] = data_i[568] & sel_one_hot_i[4];
  assign data_masked[567] = data_i[567] & sel_one_hot_i[4];
  assign data_masked[566] = data_i[566] & sel_one_hot_i[4];
  assign data_masked[565] = data_i[565] & sel_one_hot_i[4];
  assign data_masked[564] = data_i[564] & sel_one_hot_i[4];
  assign data_masked[563] = data_i[563] & sel_one_hot_i[4];
  assign data_masked[562] = data_i[562] & sel_one_hot_i[4];
  assign data_masked[561] = data_i[561] & sel_one_hot_i[4];
  assign data_masked[560] = data_i[560] & sel_one_hot_i[4];
  assign data_masked[559] = data_i[559] & sel_one_hot_i[4];
  assign data_masked[558] = data_i[558] & sel_one_hot_i[4];
  assign data_masked[557] = data_i[557] & sel_one_hot_i[4];
  assign data_masked[556] = data_i[556] & sel_one_hot_i[4];
  assign data_masked[555] = data_i[555] & sel_one_hot_i[4];
  assign data_masked[554] = data_i[554] & sel_one_hot_i[4];
  assign data_masked[553] = data_i[553] & sel_one_hot_i[4];
  assign data_masked[552] = data_i[552] & sel_one_hot_i[4];
  assign data_masked[551] = data_i[551] & sel_one_hot_i[4];
  assign data_masked[550] = data_i[550] & sel_one_hot_i[4];
  assign data_masked[549] = data_i[549] & sel_one_hot_i[4];
  assign data_masked[548] = data_i[548] & sel_one_hot_i[4];
  assign data_masked[547] = data_i[547] & sel_one_hot_i[4];
  assign data_masked[546] = data_i[546] & sel_one_hot_i[4];
  assign data_masked[545] = data_i[545] & sel_one_hot_i[4];
  assign data_masked[544] = data_i[544] & sel_one_hot_i[4];
  assign data_masked[543] = data_i[543] & sel_one_hot_i[4];
  assign data_masked[542] = data_i[542] & sel_one_hot_i[4];
  assign data_masked[541] = data_i[541] & sel_one_hot_i[4];
  assign data_masked[540] = data_i[540] & sel_one_hot_i[4];
  assign data_masked[539] = data_i[539] & sel_one_hot_i[4];
  assign data_masked[538] = data_i[538] & sel_one_hot_i[4];
  assign data_masked[537] = data_i[537] & sel_one_hot_i[4];
  assign data_masked[536] = data_i[536] & sel_one_hot_i[4];
  assign data_masked[535] = data_i[535] & sel_one_hot_i[4];
  assign data_masked[534] = data_i[534] & sel_one_hot_i[4];
  assign data_masked[533] = data_i[533] & sel_one_hot_i[4];
  assign data_masked[532] = data_i[532] & sel_one_hot_i[4];
  assign data_masked[531] = data_i[531] & sel_one_hot_i[4];
  assign data_masked[530] = data_i[530] & sel_one_hot_i[4];
  assign data_masked[529] = data_i[529] & sel_one_hot_i[4];
  assign data_masked[528] = data_i[528] & sel_one_hot_i[4];
  assign data_masked[527] = data_i[527] & sel_one_hot_i[4];
  assign data_masked[526] = data_i[526] & sel_one_hot_i[4];
  assign data_masked[525] = data_i[525] & sel_one_hot_i[4];
  assign data_masked[524] = data_i[524] & sel_one_hot_i[4];
  assign data_o[0] = N2 | data_masked[0];
  assign N2 = N1 | data_masked[131];
  assign N1 = N0 | data_masked[262];
  assign N0 = data_masked[524] | data_masked[393];
  assign data_o[1] = N5 | data_masked[1];
  assign N5 = N4 | data_masked[132];
  assign N4 = N3 | data_masked[263];
  assign N3 = data_masked[525] | data_masked[394];
  assign data_o[2] = N8 | data_masked[2];
  assign N8 = N7 | data_masked[133];
  assign N7 = N6 | data_masked[264];
  assign N6 = data_masked[526] | data_masked[395];
  assign data_o[3] = N11 | data_masked[3];
  assign N11 = N10 | data_masked[134];
  assign N10 = N9 | data_masked[265];
  assign N9 = data_masked[527] | data_masked[396];
  assign data_o[4] = N14 | data_masked[4];
  assign N14 = N13 | data_masked[135];
  assign N13 = N12 | data_masked[266];
  assign N12 = data_masked[528] | data_masked[397];
  assign data_o[5] = N17 | data_masked[5];
  assign N17 = N16 | data_masked[136];
  assign N16 = N15 | data_masked[267];
  assign N15 = data_masked[529] | data_masked[398];
  assign data_o[6] = N20 | data_masked[6];
  assign N20 = N19 | data_masked[137];
  assign N19 = N18 | data_masked[268];
  assign N18 = data_masked[530] | data_masked[399];
  assign data_o[7] = N23 | data_masked[7];
  assign N23 = N22 | data_masked[138];
  assign N22 = N21 | data_masked[269];
  assign N21 = data_masked[531] | data_masked[400];
  assign data_o[8] = N26 | data_masked[8];
  assign N26 = N25 | data_masked[139];
  assign N25 = N24 | data_masked[270];
  assign N24 = data_masked[532] | data_masked[401];
  assign data_o[9] = N29 | data_masked[9];
  assign N29 = N28 | data_masked[140];
  assign N28 = N27 | data_masked[271];
  assign N27 = data_masked[533] | data_masked[402];
  assign data_o[10] = N32 | data_masked[10];
  assign N32 = N31 | data_masked[141];
  assign N31 = N30 | data_masked[272];
  assign N30 = data_masked[534] | data_masked[403];
  assign data_o[11] = N35 | data_masked[11];
  assign N35 = N34 | data_masked[142];
  assign N34 = N33 | data_masked[273];
  assign N33 = data_masked[535] | data_masked[404];
  assign data_o[12] = N38 | data_masked[12];
  assign N38 = N37 | data_masked[143];
  assign N37 = N36 | data_masked[274];
  assign N36 = data_masked[536] | data_masked[405];
  assign data_o[13] = N41 | data_masked[13];
  assign N41 = N40 | data_masked[144];
  assign N40 = N39 | data_masked[275];
  assign N39 = data_masked[537] | data_masked[406];
  assign data_o[14] = N44 | data_masked[14];
  assign N44 = N43 | data_masked[145];
  assign N43 = N42 | data_masked[276];
  assign N42 = data_masked[538] | data_masked[407];
  assign data_o[15] = N47 | data_masked[15];
  assign N47 = N46 | data_masked[146];
  assign N46 = N45 | data_masked[277];
  assign N45 = data_masked[539] | data_masked[408];
  assign data_o[16] = N50 | data_masked[16];
  assign N50 = N49 | data_masked[147];
  assign N49 = N48 | data_masked[278];
  assign N48 = data_masked[540] | data_masked[409];
  assign data_o[17] = N53 | data_masked[17];
  assign N53 = N52 | data_masked[148];
  assign N52 = N51 | data_masked[279];
  assign N51 = data_masked[541] | data_masked[410];
  assign data_o[18] = N56 | data_masked[18];
  assign N56 = N55 | data_masked[149];
  assign N55 = N54 | data_masked[280];
  assign N54 = data_masked[542] | data_masked[411];
  assign data_o[19] = N59 | data_masked[19];
  assign N59 = N58 | data_masked[150];
  assign N58 = N57 | data_masked[281];
  assign N57 = data_masked[543] | data_masked[412];
  assign data_o[20] = N62 | data_masked[20];
  assign N62 = N61 | data_masked[151];
  assign N61 = N60 | data_masked[282];
  assign N60 = data_masked[544] | data_masked[413];
  assign data_o[21] = N65 | data_masked[21];
  assign N65 = N64 | data_masked[152];
  assign N64 = N63 | data_masked[283];
  assign N63 = data_masked[545] | data_masked[414];
  assign data_o[22] = N68 | data_masked[22];
  assign N68 = N67 | data_masked[153];
  assign N67 = N66 | data_masked[284];
  assign N66 = data_masked[546] | data_masked[415];
  assign data_o[23] = N71 | data_masked[23];
  assign N71 = N70 | data_masked[154];
  assign N70 = N69 | data_masked[285];
  assign N69 = data_masked[547] | data_masked[416];
  assign data_o[24] = N74 | data_masked[24];
  assign N74 = N73 | data_masked[155];
  assign N73 = N72 | data_masked[286];
  assign N72 = data_masked[548] | data_masked[417];
  assign data_o[25] = N77 | data_masked[25];
  assign N77 = N76 | data_masked[156];
  assign N76 = N75 | data_masked[287];
  assign N75 = data_masked[549] | data_masked[418];
  assign data_o[26] = N80 | data_masked[26];
  assign N80 = N79 | data_masked[157];
  assign N79 = N78 | data_masked[288];
  assign N78 = data_masked[550] | data_masked[419];
  assign data_o[27] = N83 | data_masked[27];
  assign N83 = N82 | data_masked[158];
  assign N82 = N81 | data_masked[289];
  assign N81 = data_masked[551] | data_masked[420];
  assign data_o[28] = N86 | data_masked[28];
  assign N86 = N85 | data_masked[159];
  assign N85 = N84 | data_masked[290];
  assign N84 = data_masked[552] | data_masked[421];
  assign data_o[29] = N89 | data_masked[29];
  assign N89 = N88 | data_masked[160];
  assign N88 = N87 | data_masked[291];
  assign N87 = data_masked[553] | data_masked[422];
  assign data_o[30] = N92 | data_masked[30];
  assign N92 = N91 | data_masked[161];
  assign N91 = N90 | data_masked[292];
  assign N90 = data_masked[554] | data_masked[423];
  assign data_o[31] = N95 | data_masked[31];
  assign N95 = N94 | data_masked[162];
  assign N94 = N93 | data_masked[293];
  assign N93 = data_masked[555] | data_masked[424];
  assign data_o[32] = N98 | data_masked[32];
  assign N98 = N97 | data_masked[163];
  assign N97 = N96 | data_masked[294];
  assign N96 = data_masked[556] | data_masked[425];
  assign data_o[33] = N101 | data_masked[33];
  assign N101 = N100 | data_masked[164];
  assign N100 = N99 | data_masked[295];
  assign N99 = data_masked[557] | data_masked[426];
  assign data_o[34] = N104 | data_masked[34];
  assign N104 = N103 | data_masked[165];
  assign N103 = N102 | data_masked[296];
  assign N102 = data_masked[558] | data_masked[427];
  assign data_o[35] = N107 | data_masked[35];
  assign N107 = N106 | data_masked[166];
  assign N106 = N105 | data_masked[297];
  assign N105 = data_masked[559] | data_masked[428];
  assign data_o[36] = N110 | data_masked[36];
  assign N110 = N109 | data_masked[167];
  assign N109 = N108 | data_masked[298];
  assign N108 = data_masked[560] | data_masked[429];
  assign data_o[37] = N113 | data_masked[37];
  assign N113 = N112 | data_masked[168];
  assign N112 = N111 | data_masked[299];
  assign N111 = data_masked[561] | data_masked[430];
  assign data_o[38] = N116 | data_masked[38];
  assign N116 = N115 | data_masked[169];
  assign N115 = N114 | data_masked[300];
  assign N114 = data_masked[562] | data_masked[431];
  assign data_o[39] = N119 | data_masked[39];
  assign N119 = N118 | data_masked[170];
  assign N118 = N117 | data_masked[301];
  assign N117 = data_masked[563] | data_masked[432];
  assign data_o[40] = N122 | data_masked[40];
  assign N122 = N121 | data_masked[171];
  assign N121 = N120 | data_masked[302];
  assign N120 = data_masked[564] | data_masked[433];
  assign data_o[41] = N125 | data_masked[41];
  assign N125 = N124 | data_masked[172];
  assign N124 = N123 | data_masked[303];
  assign N123 = data_masked[565] | data_masked[434];
  assign data_o[42] = N128 | data_masked[42];
  assign N128 = N127 | data_masked[173];
  assign N127 = N126 | data_masked[304];
  assign N126 = data_masked[566] | data_masked[435];
  assign data_o[43] = N131 | data_masked[43];
  assign N131 = N130 | data_masked[174];
  assign N130 = N129 | data_masked[305];
  assign N129 = data_masked[567] | data_masked[436];
  assign data_o[44] = N134 | data_masked[44];
  assign N134 = N133 | data_masked[175];
  assign N133 = N132 | data_masked[306];
  assign N132 = data_masked[568] | data_masked[437];
  assign data_o[45] = N137 | data_masked[45];
  assign N137 = N136 | data_masked[176];
  assign N136 = N135 | data_masked[307];
  assign N135 = data_masked[569] | data_masked[438];
  assign data_o[46] = N140 | data_masked[46];
  assign N140 = N139 | data_masked[177];
  assign N139 = N138 | data_masked[308];
  assign N138 = data_masked[570] | data_masked[439];
  assign data_o[47] = N143 | data_masked[47];
  assign N143 = N142 | data_masked[178];
  assign N142 = N141 | data_masked[309];
  assign N141 = data_masked[571] | data_masked[440];
  assign data_o[48] = N146 | data_masked[48];
  assign N146 = N145 | data_masked[179];
  assign N145 = N144 | data_masked[310];
  assign N144 = data_masked[572] | data_masked[441];
  assign data_o[49] = N149 | data_masked[49];
  assign N149 = N148 | data_masked[180];
  assign N148 = N147 | data_masked[311];
  assign N147 = data_masked[573] | data_masked[442];
  assign data_o[50] = N152 | data_masked[50];
  assign N152 = N151 | data_masked[181];
  assign N151 = N150 | data_masked[312];
  assign N150 = data_masked[574] | data_masked[443];
  assign data_o[51] = N155 | data_masked[51];
  assign N155 = N154 | data_masked[182];
  assign N154 = N153 | data_masked[313];
  assign N153 = data_masked[575] | data_masked[444];
  assign data_o[52] = N158 | data_masked[52];
  assign N158 = N157 | data_masked[183];
  assign N157 = N156 | data_masked[314];
  assign N156 = data_masked[576] | data_masked[445];
  assign data_o[53] = N161 | data_masked[53];
  assign N161 = N160 | data_masked[184];
  assign N160 = N159 | data_masked[315];
  assign N159 = data_masked[577] | data_masked[446];
  assign data_o[54] = N164 | data_masked[54];
  assign N164 = N163 | data_masked[185];
  assign N163 = N162 | data_masked[316];
  assign N162 = data_masked[578] | data_masked[447];
  assign data_o[55] = N167 | data_masked[55];
  assign N167 = N166 | data_masked[186];
  assign N166 = N165 | data_masked[317];
  assign N165 = data_masked[579] | data_masked[448];
  assign data_o[56] = N170 | data_masked[56];
  assign N170 = N169 | data_masked[187];
  assign N169 = N168 | data_masked[318];
  assign N168 = data_masked[580] | data_masked[449];
  assign data_o[57] = N173 | data_masked[57];
  assign N173 = N172 | data_masked[188];
  assign N172 = N171 | data_masked[319];
  assign N171 = data_masked[581] | data_masked[450];
  assign data_o[58] = N176 | data_masked[58];
  assign N176 = N175 | data_masked[189];
  assign N175 = N174 | data_masked[320];
  assign N174 = data_masked[582] | data_masked[451];
  assign data_o[59] = N179 | data_masked[59];
  assign N179 = N178 | data_masked[190];
  assign N178 = N177 | data_masked[321];
  assign N177 = data_masked[583] | data_masked[452];
  assign data_o[60] = N182 | data_masked[60];
  assign N182 = N181 | data_masked[191];
  assign N181 = N180 | data_masked[322];
  assign N180 = data_masked[584] | data_masked[453];
  assign data_o[61] = N185 | data_masked[61];
  assign N185 = N184 | data_masked[192];
  assign N184 = N183 | data_masked[323];
  assign N183 = data_masked[585] | data_masked[454];
  assign data_o[62] = N188 | data_masked[62];
  assign N188 = N187 | data_masked[193];
  assign N187 = N186 | data_masked[324];
  assign N186 = data_masked[586] | data_masked[455];
  assign data_o[63] = N191 | data_masked[63];
  assign N191 = N190 | data_masked[194];
  assign N190 = N189 | data_masked[325];
  assign N189 = data_masked[587] | data_masked[456];
  assign data_o[64] = N194 | data_masked[64];
  assign N194 = N193 | data_masked[195];
  assign N193 = N192 | data_masked[326];
  assign N192 = data_masked[588] | data_masked[457];
  assign data_o[65] = N197 | data_masked[65];
  assign N197 = N196 | data_masked[196];
  assign N196 = N195 | data_masked[327];
  assign N195 = data_masked[589] | data_masked[458];
  assign data_o[66] = N200 | data_masked[66];
  assign N200 = N199 | data_masked[197];
  assign N199 = N198 | data_masked[328];
  assign N198 = data_masked[590] | data_masked[459];
  assign data_o[67] = N203 | data_masked[67];
  assign N203 = N202 | data_masked[198];
  assign N202 = N201 | data_masked[329];
  assign N201 = data_masked[591] | data_masked[460];
  assign data_o[68] = N206 | data_masked[68];
  assign N206 = N205 | data_masked[199];
  assign N205 = N204 | data_masked[330];
  assign N204 = data_masked[592] | data_masked[461];
  assign data_o[69] = N209 | data_masked[69];
  assign N209 = N208 | data_masked[200];
  assign N208 = N207 | data_masked[331];
  assign N207 = data_masked[593] | data_masked[462];
  assign data_o[70] = N212 | data_masked[70];
  assign N212 = N211 | data_masked[201];
  assign N211 = N210 | data_masked[332];
  assign N210 = data_masked[594] | data_masked[463];
  assign data_o[71] = N215 | data_masked[71];
  assign N215 = N214 | data_masked[202];
  assign N214 = N213 | data_masked[333];
  assign N213 = data_masked[595] | data_masked[464];
  assign data_o[72] = N218 | data_masked[72];
  assign N218 = N217 | data_masked[203];
  assign N217 = N216 | data_masked[334];
  assign N216 = data_masked[596] | data_masked[465];
  assign data_o[73] = N221 | data_masked[73];
  assign N221 = N220 | data_masked[204];
  assign N220 = N219 | data_masked[335];
  assign N219 = data_masked[597] | data_masked[466];
  assign data_o[74] = N224 | data_masked[74];
  assign N224 = N223 | data_masked[205];
  assign N223 = N222 | data_masked[336];
  assign N222 = data_masked[598] | data_masked[467];
  assign data_o[75] = N227 | data_masked[75];
  assign N227 = N226 | data_masked[206];
  assign N226 = N225 | data_masked[337];
  assign N225 = data_masked[599] | data_masked[468];
  assign data_o[76] = N230 | data_masked[76];
  assign N230 = N229 | data_masked[207];
  assign N229 = N228 | data_masked[338];
  assign N228 = data_masked[600] | data_masked[469];
  assign data_o[77] = N233 | data_masked[77];
  assign N233 = N232 | data_masked[208];
  assign N232 = N231 | data_masked[339];
  assign N231 = data_masked[601] | data_masked[470];
  assign data_o[78] = N236 | data_masked[78];
  assign N236 = N235 | data_masked[209];
  assign N235 = N234 | data_masked[340];
  assign N234 = data_masked[602] | data_masked[471];
  assign data_o[79] = N239 | data_masked[79];
  assign N239 = N238 | data_masked[210];
  assign N238 = N237 | data_masked[341];
  assign N237 = data_masked[603] | data_masked[472];
  assign data_o[80] = N242 | data_masked[80];
  assign N242 = N241 | data_masked[211];
  assign N241 = N240 | data_masked[342];
  assign N240 = data_masked[604] | data_masked[473];
  assign data_o[81] = N245 | data_masked[81];
  assign N245 = N244 | data_masked[212];
  assign N244 = N243 | data_masked[343];
  assign N243 = data_masked[605] | data_masked[474];
  assign data_o[82] = N248 | data_masked[82];
  assign N248 = N247 | data_masked[213];
  assign N247 = N246 | data_masked[344];
  assign N246 = data_masked[606] | data_masked[475];
  assign data_o[83] = N251 | data_masked[83];
  assign N251 = N250 | data_masked[214];
  assign N250 = N249 | data_masked[345];
  assign N249 = data_masked[607] | data_masked[476];
  assign data_o[84] = N254 | data_masked[84];
  assign N254 = N253 | data_masked[215];
  assign N253 = N252 | data_masked[346];
  assign N252 = data_masked[608] | data_masked[477];
  assign data_o[85] = N257 | data_masked[85];
  assign N257 = N256 | data_masked[216];
  assign N256 = N255 | data_masked[347];
  assign N255 = data_masked[609] | data_masked[478];
  assign data_o[86] = N260 | data_masked[86];
  assign N260 = N259 | data_masked[217];
  assign N259 = N258 | data_masked[348];
  assign N258 = data_masked[610] | data_masked[479];
  assign data_o[87] = N263 | data_masked[87];
  assign N263 = N262 | data_masked[218];
  assign N262 = N261 | data_masked[349];
  assign N261 = data_masked[611] | data_masked[480];
  assign data_o[88] = N266 | data_masked[88];
  assign N266 = N265 | data_masked[219];
  assign N265 = N264 | data_masked[350];
  assign N264 = data_masked[612] | data_masked[481];
  assign data_o[89] = N269 | data_masked[89];
  assign N269 = N268 | data_masked[220];
  assign N268 = N267 | data_masked[351];
  assign N267 = data_masked[613] | data_masked[482];
  assign data_o[90] = N272 | data_masked[90];
  assign N272 = N271 | data_masked[221];
  assign N271 = N270 | data_masked[352];
  assign N270 = data_masked[614] | data_masked[483];
  assign data_o[91] = N275 | data_masked[91];
  assign N275 = N274 | data_masked[222];
  assign N274 = N273 | data_masked[353];
  assign N273 = data_masked[615] | data_masked[484];
  assign data_o[92] = N278 | data_masked[92];
  assign N278 = N277 | data_masked[223];
  assign N277 = N276 | data_masked[354];
  assign N276 = data_masked[616] | data_masked[485];
  assign data_o[93] = N281 | data_masked[93];
  assign N281 = N280 | data_masked[224];
  assign N280 = N279 | data_masked[355];
  assign N279 = data_masked[617] | data_masked[486];
  assign data_o[94] = N284 | data_masked[94];
  assign N284 = N283 | data_masked[225];
  assign N283 = N282 | data_masked[356];
  assign N282 = data_masked[618] | data_masked[487];
  assign data_o[95] = N287 | data_masked[95];
  assign N287 = N286 | data_masked[226];
  assign N286 = N285 | data_masked[357];
  assign N285 = data_masked[619] | data_masked[488];
  assign data_o[96] = N290 | data_masked[96];
  assign N290 = N289 | data_masked[227];
  assign N289 = N288 | data_masked[358];
  assign N288 = data_masked[620] | data_masked[489];
  assign data_o[97] = N293 | data_masked[97];
  assign N293 = N292 | data_masked[228];
  assign N292 = N291 | data_masked[359];
  assign N291 = data_masked[621] | data_masked[490];
  assign data_o[98] = N296 | data_masked[98];
  assign N296 = N295 | data_masked[229];
  assign N295 = N294 | data_masked[360];
  assign N294 = data_masked[622] | data_masked[491];
  assign data_o[99] = N299 | data_masked[99];
  assign N299 = N298 | data_masked[230];
  assign N298 = N297 | data_masked[361];
  assign N297 = data_masked[623] | data_masked[492];
  assign data_o[100] = N302 | data_masked[100];
  assign N302 = N301 | data_masked[231];
  assign N301 = N300 | data_masked[362];
  assign N300 = data_masked[624] | data_masked[493];
  assign data_o[101] = N305 | data_masked[101];
  assign N305 = N304 | data_masked[232];
  assign N304 = N303 | data_masked[363];
  assign N303 = data_masked[625] | data_masked[494];
  assign data_o[102] = N308 | data_masked[102];
  assign N308 = N307 | data_masked[233];
  assign N307 = N306 | data_masked[364];
  assign N306 = data_masked[626] | data_masked[495];
  assign data_o[103] = N311 | data_masked[103];
  assign N311 = N310 | data_masked[234];
  assign N310 = N309 | data_masked[365];
  assign N309 = data_masked[627] | data_masked[496];
  assign data_o[104] = N314 | data_masked[104];
  assign N314 = N313 | data_masked[235];
  assign N313 = N312 | data_masked[366];
  assign N312 = data_masked[628] | data_masked[497];
  assign data_o[105] = N317 | data_masked[105];
  assign N317 = N316 | data_masked[236];
  assign N316 = N315 | data_masked[367];
  assign N315 = data_masked[629] | data_masked[498];
  assign data_o[106] = N320 | data_masked[106];
  assign N320 = N319 | data_masked[237];
  assign N319 = N318 | data_masked[368];
  assign N318 = data_masked[630] | data_masked[499];
  assign data_o[107] = N323 | data_masked[107];
  assign N323 = N322 | data_masked[238];
  assign N322 = N321 | data_masked[369];
  assign N321 = data_masked[631] | data_masked[500];
  assign data_o[108] = N326 | data_masked[108];
  assign N326 = N325 | data_masked[239];
  assign N325 = N324 | data_masked[370];
  assign N324 = data_masked[632] | data_masked[501];
  assign data_o[109] = N329 | data_masked[109];
  assign N329 = N328 | data_masked[240];
  assign N328 = N327 | data_masked[371];
  assign N327 = data_masked[633] | data_masked[502];
  assign data_o[110] = N332 | data_masked[110];
  assign N332 = N331 | data_masked[241];
  assign N331 = N330 | data_masked[372];
  assign N330 = data_masked[634] | data_masked[503];
  assign data_o[111] = N335 | data_masked[111];
  assign N335 = N334 | data_masked[242];
  assign N334 = N333 | data_masked[373];
  assign N333 = data_masked[635] | data_masked[504];
  assign data_o[112] = N338 | data_masked[112];
  assign N338 = N337 | data_masked[243];
  assign N337 = N336 | data_masked[374];
  assign N336 = data_masked[636] | data_masked[505];
  assign data_o[113] = N341 | data_masked[113];
  assign N341 = N340 | data_masked[244];
  assign N340 = N339 | data_masked[375];
  assign N339 = data_masked[637] | data_masked[506];
  assign data_o[114] = N344 | data_masked[114];
  assign N344 = N343 | data_masked[245];
  assign N343 = N342 | data_masked[376];
  assign N342 = data_masked[638] | data_masked[507];
  assign data_o[115] = N347 | data_masked[115];
  assign N347 = N346 | data_masked[246];
  assign N346 = N345 | data_masked[377];
  assign N345 = data_masked[639] | data_masked[508];
  assign data_o[116] = N350 | data_masked[116];
  assign N350 = N349 | data_masked[247];
  assign N349 = N348 | data_masked[378];
  assign N348 = data_masked[640] | data_masked[509];
  assign data_o[117] = N353 | data_masked[117];
  assign N353 = N352 | data_masked[248];
  assign N352 = N351 | data_masked[379];
  assign N351 = data_masked[641] | data_masked[510];
  assign data_o[118] = N356 | data_masked[118];
  assign N356 = N355 | data_masked[249];
  assign N355 = N354 | data_masked[380];
  assign N354 = data_masked[642] | data_masked[511];
  assign data_o[119] = N359 | data_masked[119];
  assign N359 = N358 | data_masked[250];
  assign N358 = N357 | data_masked[381];
  assign N357 = data_masked[643] | data_masked[512];
  assign data_o[120] = N362 | data_masked[120];
  assign N362 = N361 | data_masked[251];
  assign N361 = N360 | data_masked[382];
  assign N360 = data_masked[644] | data_masked[513];
  assign data_o[121] = N365 | data_masked[121];
  assign N365 = N364 | data_masked[252];
  assign N364 = N363 | data_masked[383];
  assign N363 = data_masked[645] | data_masked[514];
  assign data_o[122] = N368 | data_masked[122];
  assign N368 = N367 | data_masked[253];
  assign N367 = N366 | data_masked[384];
  assign N366 = data_masked[646] | data_masked[515];
  assign data_o[123] = N371 | data_masked[123];
  assign N371 = N370 | data_masked[254];
  assign N370 = N369 | data_masked[385];
  assign N369 = data_masked[647] | data_masked[516];
  assign data_o[124] = N374 | data_masked[124];
  assign N374 = N373 | data_masked[255];
  assign N373 = N372 | data_masked[386];
  assign N372 = data_masked[648] | data_masked[517];
  assign data_o[125] = N377 | data_masked[125];
  assign N377 = N376 | data_masked[256];
  assign N376 = N375 | data_masked[387];
  assign N375 = data_masked[649] | data_masked[518];
  assign data_o[126] = N380 | data_masked[126];
  assign N380 = N379 | data_masked[257];
  assign N379 = N378 | data_masked[388];
  assign N378 = data_masked[650] | data_masked[519];
  assign data_o[127] = N383 | data_masked[127];
  assign N383 = N382 | data_masked[258];
  assign N382 = N381 | data_masked[389];
  assign N381 = data_masked[651] | data_masked[520];
  assign data_o[128] = N386 | data_masked[128];
  assign N386 = N385 | data_masked[259];
  assign N385 = N384 | data_masked[390];
  assign N384 = data_masked[652] | data_masked[521];
  assign data_o[129] = N389 | data_masked[129];
  assign N389 = N388 | data_masked[260];
  assign N388 = N387 | data_masked[391];
  assign N387 = data_masked[653] | data_masked[522];
  assign data_o[130] = N392 | data_masked[130];
  assign N392 = N391 | data_masked[261];
  assign N391 = N390 | data_masked[392];
  assign N390 = data_masked[654] | data_masked[523];

endmodule



module bsg_wormhole_router_131_1_1_2_1_1_1_00000003_0000001a
(
  clk_i,
  reset_i,
  local_x_cord_i,
  local_y_cord_i,
  valid_i,
  data_i,
  ready_o,
  valid_o,
  data_o,
  ready_i
);

  input [0:0] local_x_cord_i;
  input [0:0] local_y_cord_i;
  input [4:0] valid_i;
  input [654:0] data_i;
  output [4:0] ready_o;
  output [4:0] valid_o;
  output [654:0] data_o;
  input [4:0] ready_i;
  input clk_i;
  input reset_i;
  wire [4:0] ready_o,valid_o,fifo_yumi_i;
  wire [654:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,fifo_data_o_4__130_,fifo_data_o_4__129_,
  fifo_data_o_4__128_,fifo_data_o_4__127_,fifo_data_o_4__126_,fifo_data_o_4__125_,
  fifo_data_o_4__124_,fifo_data_o_4__123_,fifo_data_o_4__122_,fifo_data_o_4__121_,
  fifo_data_o_4__120_,fifo_data_o_4__119_,fifo_data_o_4__118_,fifo_data_o_4__117_,
  fifo_data_o_4__116_,fifo_data_o_4__115_,fifo_data_o_4__114_,fifo_data_o_4__113_,
  fifo_data_o_4__112_,fifo_data_o_4__111_,fifo_data_o_4__110_,fifo_data_o_4__109_,
  fifo_data_o_4__108_,fifo_data_o_4__107_,fifo_data_o_4__106_,fifo_data_o_4__105_,
  fifo_data_o_4__104_,fifo_data_o_4__103_,fifo_data_o_4__102_,fifo_data_o_4__101_,
  fifo_data_o_4__100_,fifo_data_o_4__99_,fifo_data_o_4__98_,fifo_data_o_4__97_,
  fifo_data_o_4__96_,fifo_data_o_4__95_,fifo_data_o_4__94_,fifo_data_o_4__93_,
  fifo_data_o_4__92_,fifo_data_o_4__91_,fifo_data_o_4__90_,fifo_data_o_4__89_,
  fifo_data_o_4__88_,fifo_data_o_4__87_,fifo_data_o_4__86_,fifo_data_o_4__85_,
  fifo_data_o_4__84_,fifo_data_o_4__83_,fifo_data_o_4__82_,fifo_data_o_4__81_,fifo_data_o_4__80_,
  fifo_data_o_4__79_,fifo_data_o_4__78_,fifo_data_o_4__77_,fifo_data_o_4__76_,
  fifo_data_o_4__75_,fifo_data_o_4__74_,fifo_data_o_4__73_,fifo_data_o_4__72_,
  fifo_data_o_4__71_,fifo_data_o_4__70_,fifo_data_o_4__69_,fifo_data_o_4__68_,
  fifo_data_o_4__67_,fifo_data_o_4__66_,fifo_data_o_4__65_,fifo_data_o_4__64_,
  fifo_data_o_4__63_,fifo_data_o_4__62_,fifo_data_o_4__61_,fifo_data_o_4__60_,fifo_data_o_4__59_,
  fifo_data_o_4__58_,fifo_data_o_4__57_,fifo_data_o_4__56_,fifo_data_o_4__55_,
  fifo_data_o_4__54_,fifo_data_o_4__53_,fifo_data_o_4__52_,fifo_data_o_4__51_,
  fifo_data_o_4__50_,fifo_data_o_4__49_,fifo_data_o_4__48_,fifo_data_o_4__47_,
  fifo_data_o_4__46_,fifo_data_o_4__45_,fifo_data_o_4__44_,fifo_data_o_4__43_,
  fifo_data_o_4__42_,fifo_data_o_4__41_,fifo_data_o_4__40_,fifo_data_o_4__39_,fifo_data_o_4__38_,
  fifo_data_o_4__37_,fifo_data_o_4__36_,fifo_data_o_4__35_,fifo_data_o_4__34_,
  fifo_data_o_4__33_,fifo_data_o_4__32_,fifo_data_o_4__31_,fifo_data_o_4__30_,
  fifo_data_o_4__29_,fifo_data_o_4__28_,fifo_data_o_4__27_,fifo_data_o_4__26_,
  fifo_data_o_4__25_,fifo_data_o_4__24_,fifo_data_o_4__23_,fifo_data_o_4__22_,
  fifo_data_o_4__21_,fifo_data_o_4__20_,fifo_data_o_4__19_,fifo_data_o_4__18_,fifo_data_o_4__17_,
  fifo_data_o_4__16_,fifo_data_o_4__15_,fifo_data_o_4__14_,fifo_data_o_4__13_,
  fifo_data_o_4__12_,fifo_data_o_4__11_,fifo_data_o_4__10_,fifo_data_o_4__9_,
  fifo_data_o_4__8_,fifo_data_o_4__7_,fifo_data_o_4__6_,fifo_data_o_4__5_,fifo_data_o_4__4_,
  fifo_data_o_4__3_,fifo_data_o_4__2_,fifo_data_o_4__1_,fifo_data_o_4__0_,
  fifo_data_o_3__130_,fifo_data_o_3__129_,fifo_data_o_3__128_,fifo_data_o_3__127_,
  fifo_data_o_3__126_,fifo_data_o_3__125_,fifo_data_o_3__124_,fifo_data_o_3__123_,
  fifo_data_o_3__122_,fifo_data_o_3__121_,fifo_data_o_3__120_,fifo_data_o_3__119_,
  fifo_data_o_3__118_,fifo_data_o_3__117_,fifo_data_o_3__116_,fifo_data_o_3__115_,
  fifo_data_o_3__114_,fifo_data_o_3__113_,fifo_data_o_3__112_,fifo_data_o_3__111_,
  fifo_data_o_3__110_,fifo_data_o_3__109_,fifo_data_o_3__108_,fifo_data_o_3__107_,
  fifo_data_o_3__106_,fifo_data_o_3__105_,fifo_data_o_3__104_,fifo_data_o_3__103_,
  fifo_data_o_3__102_,fifo_data_o_3__101_,fifo_data_o_3__100_,fifo_data_o_3__99_,
  fifo_data_o_3__98_,fifo_data_o_3__97_,fifo_data_o_3__96_,fifo_data_o_3__95_,
  fifo_data_o_3__94_,fifo_data_o_3__93_,fifo_data_o_3__92_,fifo_data_o_3__91_,fifo_data_o_3__90_,
  fifo_data_o_3__89_,fifo_data_o_3__88_,fifo_data_o_3__87_,fifo_data_o_3__86_,
  fifo_data_o_3__85_,fifo_data_o_3__84_,fifo_data_o_3__83_,fifo_data_o_3__82_,
  fifo_data_o_3__81_,fifo_data_o_3__80_,fifo_data_o_3__79_,fifo_data_o_3__78_,
  fifo_data_o_3__77_,fifo_data_o_3__76_,fifo_data_o_3__75_,fifo_data_o_3__74_,
  fifo_data_o_3__73_,fifo_data_o_3__72_,fifo_data_o_3__71_,fifo_data_o_3__70_,fifo_data_o_3__69_,
  fifo_data_o_3__68_,fifo_data_o_3__67_,fifo_data_o_3__66_,fifo_data_o_3__65_,
  fifo_data_o_3__64_,fifo_data_o_3__63_,fifo_data_o_3__62_,fifo_data_o_3__61_,
  fifo_data_o_3__60_,fifo_data_o_3__59_,fifo_data_o_3__58_,fifo_data_o_3__57_,
  fifo_data_o_3__56_,fifo_data_o_3__55_,fifo_data_o_3__54_,fifo_data_o_3__53_,
  fifo_data_o_3__52_,fifo_data_o_3__51_,fifo_data_o_3__50_,fifo_data_o_3__49_,fifo_data_o_3__48_,
  fifo_data_o_3__47_,fifo_data_o_3__46_,fifo_data_o_3__45_,fifo_data_o_3__44_,
  fifo_data_o_3__43_,fifo_data_o_3__42_,fifo_data_o_3__41_,fifo_data_o_3__40_,
  fifo_data_o_3__39_,fifo_data_o_3__38_,fifo_data_o_3__37_,fifo_data_o_3__36_,
  fifo_data_o_3__35_,fifo_data_o_3__34_,fifo_data_o_3__33_,fifo_data_o_3__32_,
  fifo_data_o_3__31_,fifo_data_o_3__30_,fifo_data_o_3__29_,fifo_data_o_3__28_,fifo_data_o_3__27_,
  fifo_data_o_3__26_,fifo_data_o_3__25_,fifo_data_o_3__24_,fifo_data_o_3__23_,
  fifo_data_o_3__22_,fifo_data_o_3__21_,fifo_data_o_3__20_,fifo_data_o_3__19_,
  fifo_data_o_3__18_,fifo_data_o_3__17_,fifo_data_o_3__16_,fifo_data_o_3__15_,
  fifo_data_o_3__14_,fifo_data_o_3__13_,fifo_data_o_3__12_,fifo_data_o_3__11_,fifo_data_o_3__10_,
  fifo_data_o_3__9_,fifo_data_o_3__8_,fifo_data_o_3__7_,fifo_data_o_3__6_,
  fifo_data_o_3__5_,fifo_data_o_3__4_,fifo_data_o_3__3_,fifo_data_o_3__2_,
  fifo_data_o_3__1_,fifo_data_o_3__0_,fifo_data_o_2__130_,fifo_data_o_2__129_,fifo_data_o_2__128_,
  fifo_data_o_2__127_,fifo_data_o_2__126_,fifo_data_o_2__125_,fifo_data_o_2__124_,
  fifo_data_o_2__123_,fifo_data_o_2__122_,fifo_data_o_2__121_,fifo_data_o_2__120_,
  fifo_data_o_2__119_,fifo_data_o_2__118_,fifo_data_o_2__117_,fifo_data_o_2__116_,
  fifo_data_o_2__115_,fifo_data_o_2__114_,fifo_data_o_2__113_,fifo_data_o_2__112_,
  fifo_data_o_2__111_,fifo_data_o_2__110_,fifo_data_o_2__109_,fifo_data_o_2__108_,
  fifo_data_o_2__107_,fifo_data_o_2__106_,fifo_data_o_2__105_,fifo_data_o_2__104_,
  fifo_data_o_2__103_,fifo_data_o_2__102_,fifo_data_o_2__101_,fifo_data_o_2__100_,
  fifo_data_o_2__99_,fifo_data_o_2__98_,fifo_data_o_2__97_,fifo_data_o_2__96_,
  fifo_data_o_2__95_,fifo_data_o_2__94_,fifo_data_o_2__93_,fifo_data_o_2__92_,
  fifo_data_o_2__91_,fifo_data_o_2__90_,fifo_data_o_2__89_,fifo_data_o_2__88_,
  fifo_data_o_2__87_,fifo_data_o_2__86_,fifo_data_o_2__85_,fifo_data_o_2__84_,
  fifo_data_o_2__83_,fifo_data_o_2__82_,fifo_data_o_2__81_,fifo_data_o_2__80_,fifo_data_o_2__79_,
  fifo_data_o_2__78_,fifo_data_o_2__77_,fifo_data_o_2__76_,fifo_data_o_2__75_,
  fifo_data_o_2__74_,fifo_data_o_2__73_,fifo_data_o_2__72_,fifo_data_o_2__71_,
  fifo_data_o_2__70_,fifo_data_o_2__69_,fifo_data_o_2__68_,fifo_data_o_2__67_,
  fifo_data_o_2__66_,fifo_data_o_2__65_,fifo_data_o_2__64_,fifo_data_o_2__63_,
  fifo_data_o_2__62_,fifo_data_o_2__61_,fifo_data_o_2__60_,fifo_data_o_2__59_,fifo_data_o_2__58_,
  fifo_data_o_2__57_,fifo_data_o_2__56_,fifo_data_o_2__55_,fifo_data_o_2__54_,
  fifo_data_o_2__53_,fifo_data_o_2__52_,fifo_data_o_2__51_,fifo_data_o_2__50_,
  fifo_data_o_2__49_,fifo_data_o_2__48_,fifo_data_o_2__47_,fifo_data_o_2__46_,
  fifo_data_o_2__45_,fifo_data_o_2__44_,fifo_data_o_2__43_,fifo_data_o_2__42_,
  fifo_data_o_2__41_,fifo_data_o_2__40_,fifo_data_o_2__39_,fifo_data_o_2__38_,fifo_data_o_2__37_,
  fifo_data_o_2__36_,fifo_data_o_2__35_,fifo_data_o_2__34_,fifo_data_o_2__33_,
  fifo_data_o_2__32_,fifo_data_o_2__31_,fifo_data_o_2__30_,fifo_data_o_2__29_,
  fifo_data_o_2__28_,fifo_data_o_2__27_,fifo_data_o_2__26_,fifo_data_o_2__25_,
  fifo_data_o_2__24_,fifo_data_o_2__23_,fifo_data_o_2__22_,fifo_data_o_2__21_,fifo_data_o_2__20_,
  fifo_data_o_2__19_,fifo_data_o_2__18_,fifo_data_o_2__17_,fifo_data_o_2__16_,
  fifo_data_o_2__15_,fifo_data_o_2__14_,fifo_data_o_2__13_,fifo_data_o_2__12_,
  fifo_data_o_2__11_,fifo_data_o_2__10_,fifo_data_o_2__9_,fifo_data_o_2__8_,
  fifo_data_o_2__7_,fifo_data_o_2__6_,fifo_data_o_2__5_,fifo_data_o_2__4_,fifo_data_o_2__3_,
  fifo_data_o_2__2_,fifo_data_o_2__1_,fifo_data_o_2__0_,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
  dest_n_4__3_,dest_n_4__2_,dest_n_4__1_,dest_n_4__0_,dest_n_3__4_,dest_n_3__2_,
  dest_n_3__1_,dest_n_3__0_,dest_n_2__4_,dest_n_2__3_,dest_n_2__1_,dest_n_2__0_,dest_n_1__4_,
  dest_n_1__3_,dest_n_1__2_,dest_n_1__0_,dest_n_0__4_,dest_n_0__3_,dest_n_0__2_,
  dest_n_0__1_,dest_n_0__0_,new_valid_4__3_,new_valid_4__2_,new_valid_4__1_,
  new_valid_4__0_,new_valid_3__4_,new_valid_3__2_,new_valid_3__1_,new_valid_3__0_,
  new_valid_2__4_,new_valid_2__3_,new_valid_2__1_,new_valid_2__0_,new_valid_1__4_,
  new_valid_1__3_,new_valid_1__2_,new_valid_1__0_,new_valid_0__4_,new_valid_0__3_,
  new_valid_0__2_,new_valid_0__1_,new_valid_0__0_,arb_grants_o_4__3_,arb_grants_o_4__2_,
  arb_grants_o_4__1_,arb_grants_o_4__0_,arb_grants_o_3__4_,arb_grants_o_3__2_,
  arb_grants_o_3__1_,arb_grants_o_3__0_,arb_grants_o_2__4_,arb_grants_o_2__3_,
  arb_grants_o_2__1_,arb_grants_o_2__0_,arb_grants_o_1__4_,arb_grants_o_1__3_,
  arb_grants_o_1__2_,arb_grants_o_1__0_,arb_grants_o_0__4_,arb_grants_o_0__3_,arb_grants_o_0__2_,
  arb_grants_o_0__1_,arb_grants_o_0__0_,N194,N195,N196,N197,N198,N199,N200,N201,
  N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,
  N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,
  N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,
  N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,
  arb_valid_4__3_,arb_valid_4__2_,arb_valid_4__1_,arb_valid_4__0_,arb_valid_3__4_,
  arb_valid_3__2_,arb_valid_3__1_,arb_valid_3__0_,arb_valid_2__4_,arb_valid_2__3_,
  arb_valid_2__1_,arb_valid_2__0_,arb_valid_1__4_,arb_valid_1__3_,arb_valid_1__2_,
  arb_valid_1__0_,arb_valid_0__4_,arb_valid_0__3_,arb_valid_0__2_,arb_valid_0__1_,
  arb_valid_0__0_,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,
  N279,N280,N281,N282,N283,N284,n_3_net_,arb_sel_o_4__3_,arb_sel_o_4__2_,
  arb_sel_o_4__1_,arb_sel_o_4__0_,arb_sel_o_3__3_,arb_sel_o_3__2_,arb_sel_o_3__1_,
  arb_sel_o_3__0_,arb_sel_o_2__3_,arb_sel_o_2__2_,arb_sel_o_2__1_,arb_sel_o_2__0_,
  arb_sel_o_1__3_,arb_sel_o_1__2_,arb_sel_o_1__1_,arb_sel_o_1__0_,arb_sel_o_0__4_,
  arb_sel_o_0__3_,arb_sel_o_0__2_,arb_sel_o_0__1_,arb_sel_o_0__0_,n_9_net_,n_15_net_,
  n_21_net_,n_27_net_,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,
  N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,
  N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,
  N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,
  N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,
  N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,
  N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,
  N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,
  N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,
  N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,
  N442,N443,N444,N445,N446,N447,N448,SV2V_UNCONNECTED_1,SV2V_UNCONNECTED_2,
  SV2V_UNCONNECTED_3,SV2V_UNCONNECTED_4,SV2V_UNCONNECTED_5,
  SV2V_UNCONNECTED_6,SV2V_UNCONNECTED_7,SV2V_UNCONNECTED_8,SV2V_UNCONNECTED_9,
  SV2V_UNCONNECTED_10,SV2V_UNCONNECTED_11;
  wire [4:2] fifo_valid_o;
  reg [9:0] count_r,out_count_r;
  reg dest_r_0__4_,dest_r_0__3_,dest_r_0__2_,dest_r_0__1_,dest_r_0__0_,dest_r_1__4_,
  dest_r_1__3_,dest_r_1__2_,dest_r_1__0_,dest_r_2__4_,dest_r_2__3_,dest_r_2__1_,
  dest_r_2__0_,dest_r_3__4_,dest_r_3__2_,dest_r_3__1_,dest_r_3__0_,dest_r_4__3_,
  dest_r_4__2_,dest_r_4__1_,dest_r_4__0_,arb_grants_r_0__0_,arb_grants_r_0__1_,
  arb_grants_r_0__2_,arb_grants_r_0__3_,arb_grants_r_0__4_,arb_grants_r_1__0_,
  arb_grants_r_1__2_,arb_grants_r_1__3_,arb_grants_r_1__4_,arb_grants_r_2__0_,
  arb_grants_r_2__1_,arb_grants_r_2__3_,arb_grants_r_2__4_,arb_grants_r_3__0_,arb_grants_r_3__1_,
  arb_grants_r_3__2_,arb_grants_r_3__4_,arb_grants_r_4__0_,arb_grants_r_4__1_,
  arb_grants_r_4__2_,arb_grants_r_4__3_;
  assign ready_o[1] = 1'b1;
  assign ready_o[0] = 1'b1;

  bsg_two_fifo_width_p131
  in_ff_2__no_stub_two_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(ready_o[2]),
    .data_i(data_i[392:262]),
    .v_i(valid_i[2]),
    .v_o(fifo_valid_o[2]),
    .data_o({ fifo_data_o_2__130_, fifo_data_o_2__129_, fifo_data_o_2__128_, fifo_data_o_2__127_, fifo_data_o_2__126_, fifo_data_o_2__125_, fifo_data_o_2__124_, fifo_data_o_2__123_, fifo_data_o_2__122_, fifo_data_o_2__121_, fifo_data_o_2__120_, fifo_data_o_2__119_, fifo_data_o_2__118_, fifo_data_o_2__117_, fifo_data_o_2__116_, fifo_data_o_2__115_, fifo_data_o_2__114_, fifo_data_o_2__113_, fifo_data_o_2__112_, fifo_data_o_2__111_, fifo_data_o_2__110_, fifo_data_o_2__109_, fifo_data_o_2__108_, fifo_data_o_2__107_, fifo_data_o_2__106_, fifo_data_o_2__105_, fifo_data_o_2__104_, fifo_data_o_2__103_, fifo_data_o_2__102_, fifo_data_o_2__101_, fifo_data_o_2__100_, fifo_data_o_2__99_, fifo_data_o_2__98_, fifo_data_o_2__97_, fifo_data_o_2__96_, fifo_data_o_2__95_, fifo_data_o_2__94_, fifo_data_o_2__93_, fifo_data_o_2__92_, fifo_data_o_2__91_, fifo_data_o_2__90_, fifo_data_o_2__89_, fifo_data_o_2__88_, fifo_data_o_2__87_, fifo_data_o_2__86_, fifo_data_o_2__85_, fifo_data_o_2__84_, fifo_data_o_2__83_, fifo_data_o_2__82_, fifo_data_o_2__81_, fifo_data_o_2__80_, fifo_data_o_2__79_, fifo_data_o_2__78_, fifo_data_o_2__77_, fifo_data_o_2__76_, fifo_data_o_2__75_, fifo_data_o_2__74_, fifo_data_o_2__73_, fifo_data_o_2__72_, fifo_data_o_2__71_, fifo_data_o_2__70_, fifo_data_o_2__69_, fifo_data_o_2__68_, fifo_data_o_2__67_, fifo_data_o_2__66_, fifo_data_o_2__65_, fifo_data_o_2__64_, fifo_data_o_2__63_, fifo_data_o_2__62_, fifo_data_o_2__61_, fifo_data_o_2__60_, fifo_data_o_2__59_, fifo_data_o_2__58_, fifo_data_o_2__57_, fifo_data_o_2__56_, fifo_data_o_2__55_, fifo_data_o_2__54_, fifo_data_o_2__53_, fifo_data_o_2__52_, fifo_data_o_2__51_, fifo_data_o_2__50_, fifo_data_o_2__49_, fifo_data_o_2__48_, fifo_data_o_2__47_, fifo_data_o_2__46_, fifo_data_o_2__45_, fifo_data_o_2__44_, fifo_data_o_2__43_, fifo_data_o_2__42_, fifo_data_o_2__41_, fifo_data_o_2__40_, fifo_data_o_2__39_, fifo_data_o_2__38_, fifo_data_o_2__37_, fifo_data_o_2__36_, fifo_data_o_2__35_, fifo_data_o_2__34_, fifo_data_o_2__33_, fifo_data_o_2__32_, fifo_data_o_2__31_, fifo_data_o_2__30_, fifo_data_o_2__29_, fifo_data_o_2__28_, fifo_data_o_2__27_, fifo_data_o_2__26_, fifo_data_o_2__25_, fifo_data_o_2__24_, fifo_data_o_2__23_, fifo_data_o_2__22_, fifo_data_o_2__21_, fifo_data_o_2__20_, fifo_data_o_2__19_, fifo_data_o_2__18_, fifo_data_o_2__17_, fifo_data_o_2__16_, fifo_data_o_2__15_, fifo_data_o_2__14_, fifo_data_o_2__13_, fifo_data_o_2__12_, fifo_data_o_2__11_, fifo_data_o_2__10_, fifo_data_o_2__9_, fifo_data_o_2__8_, fifo_data_o_2__7_, fifo_data_o_2__6_, fifo_data_o_2__5_, fifo_data_o_2__4_, fifo_data_o_2__3_, fifo_data_o_2__2_, fifo_data_o_2__1_, fifo_data_o_2__0_ }),
    .yumi_i(fifo_yumi_i[2])
  );


  bsg_two_fifo_width_p131
  in_ff_3__no_stub_two_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(ready_o[3]),
    .data_i(data_i[523:393]),
    .v_i(valid_i[3]),
    .v_o(fifo_valid_o[3]),
    .data_o({ fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_ }),
    .yumi_i(fifo_yumi_i[3])
  );


  bsg_two_fifo_width_p131
  in_ff_4__no_stub_two_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(ready_o[4]),
    .data_i(data_i[654:524]),
    .v_i(valid_i[4]),
    .v_o(fifo_valid_o[4]),
    .data_o({ fifo_data_o_4__130_, fifo_data_o_4__129_, fifo_data_o_4__128_, fifo_data_o_4__127_, fifo_data_o_4__126_, fifo_data_o_4__125_, fifo_data_o_4__124_, fifo_data_o_4__123_, fifo_data_o_4__122_, fifo_data_o_4__121_, fifo_data_o_4__120_, fifo_data_o_4__119_, fifo_data_o_4__118_, fifo_data_o_4__117_, fifo_data_o_4__116_, fifo_data_o_4__115_, fifo_data_o_4__114_, fifo_data_o_4__113_, fifo_data_o_4__112_, fifo_data_o_4__111_, fifo_data_o_4__110_, fifo_data_o_4__109_, fifo_data_o_4__108_, fifo_data_o_4__107_, fifo_data_o_4__106_, fifo_data_o_4__105_, fifo_data_o_4__104_, fifo_data_o_4__103_, fifo_data_o_4__102_, fifo_data_o_4__101_, fifo_data_o_4__100_, fifo_data_o_4__99_, fifo_data_o_4__98_, fifo_data_o_4__97_, fifo_data_o_4__96_, fifo_data_o_4__95_, fifo_data_o_4__94_, fifo_data_o_4__93_, fifo_data_o_4__92_, fifo_data_o_4__91_, fifo_data_o_4__90_, fifo_data_o_4__89_, fifo_data_o_4__88_, fifo_data_o_4__87_, fifo_data_o_4__86_, fifo_data_o_4__85_, fifo_data_o_4__84_, fifo_data_o_4__83_, fifo_data_o_4__82_, fifo_data_o_4__81_, fifo_data_o_4__80_, fifo_data_o_4__79_, fifo_data_o_4__78_, fifo_data_o_4__77_, fifo_data_o_4__76_, fifo_data_o_4__75_, fifo_data_o_4__74_, fifo_data_o_4__73_, fifo_data_o_4__72_, fifo_data_o_4__71_, fifo_data_o_4__70_, fifo_data_o_4__69_, fifo_data_o_4__68_, fifo_data_o_4__67_, fifo_data_o_4__66_, fifo_data_o_4__65_, fifo_data_o_4__64_, fifo_data_o_4__63_, fifo_data_o_4__62_, fifo_data_o_4__61_, fifo_data_o_4__60_, fifo_data_o_4__59_, fifo_data_o_4__58_, fifo_data_o_4__57_, fifo_data_o_4__56_, fifo_data_o_4__55_, fifo_data_o_4__54_, fifo_data_o_4__53_, fifo_data_o_4__52_, fifo_data_o_4__51_, fifo_data_o_4__50_, fifo_data_o_4__49_, fifo_data_o_4__48_, fifo_data_o_4__47_, fifo_data_o_4__46_, fifo_data_o_4__45_, fifo_data_o_4__44_, fifo_data_o_4__43_, fifo_data_o_4__42_, fifo_data_o_4__41_, fifo_data_o_4__40_, fifo_data_o_4__39_, fifo_data_o_4__38_, fifo_data_o_4__37_, fifo_data_o_4__36_, fifo_data_o_4__35_, fifo_data_o_4__34_, fifo_data_o_4__33_, fifo_data_o_4__32_, fifo_data_o_4__31_, fifo_data_o_4__30_, fifo_data_o_4__29_, fifo_data_o_4__28_, fifo_data_o_4__27_, fifo_data_o_4__26_, fifo_data_o_4__25_, fifo_data_o_4__24_, fifo_data_o_4__23_, fifo_data_o_4__22_, fifo_data_o_4__21_, fifo_data_o_4__20_, fifo_data_o_4__19_, fifo_data_o_4__18_, fifo_data_o_4__17_, fifo_data_o_4__16_, fifo_data_o_4__15_, fifo_data_o_4__14_, fifo_data_o_4__13_, fifo_data_o_4__12_, fifo_data_o_4__11_, fifo_data_o_4__10_, fifo_data_o_4__9_, fifo_data_o_4__8_, fifo_data_o_4__7_, fifo_data_o_4__6_, fifo_data_o_4__5_, fifo_data_o_4__4_, fifo_data_o_4__3_, fifo_data_o_4__2_, fifo_data_o_4__1_, fifo_data_o_4__0_ }),
    .yumi_i(fifo_yumi_i[4])
  );


  bsg_round_robin_arb_inputs_p4
  out_side_1__rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ arb_valid_4__1_, arb_valid_3__1_, arb_valid_2__1_, arb_valid_0__1_ }),
    .grants_o({ arb_grants_o_4__1_, arb_grants_o_3__1_, arb_grants_o_2__1_, arb_grants_o_0__1_ }),
    .sel_one_hot_o({ arb_sel_o_1__3_, arb_sel_o_1__2_, arb_sel_o_1__1_, arb_sel_o_1__0_ }),
    .v_o(valid_o[1]),
    .tag_o({ SV2V_UNCONNECTED_1, SV2V_UNCONNECTED_2 }),
    .yumi_i(n_3_net_)
  );


  bsg_mux_one_hot_width_p131_els_p4
  out_side_1__mux
  (
    .data_i({ fifo_data_o_4__130_, fifo_data_o_4__129_, fifo_data_o_4__128_, fifo_data_o_4__127_, fifo_data_o_4__126_, fifo_data_o_4__125_, fifo_data_o_4__124_, fifo_data_o_4__123_, fifo_data_o_4__122_, fifo_data_o_4__121_, fifo_data_o_4__120_, fifo_data_o_4__119_, fifo_data_o_4__118_, fifo_data_o_4__117_, fifo_data_o_4__116_, fifo_data_o_4__115_, fifo_data_o_4__114_, fifo_data_o_4__113_, fifo_data_o_4__112_, fifo_data_o_4__111_, fifo_data_o_4__110_, fifo_data_o_4__109_, fifo_data_o_4__108_, fifo_data_o_4__107_, fifo_data_o_4__106_, fifo_data_o_4__105_, fifo_data_o_4__104_, fifo_data_o_4__103_, fifo_data_o_4__102_, fifo_data_o_4__101_, fifo_data_o_4__100_, fifo_data_o_4__99_, fifo_data_o_4__98_, fifo_data_o_4__97_, fifo_data_o_4__96_, fifo_data_o_4__95_, fifo_data_o_4__94_, fifo_data_o_4__93_, fifo_data_o_4__92_, fifo_data_o_4__91_, fifo_data_o_4__90_, fifo_data_o_4__89_, fifo_data_o_4__88_, fifo_data_o_4__87_, fifo_data_o_4__86_, fifo_data_o_4__85_, fifo_data_o_4__84_, fifo_data_o_4__83_, fifo_data_o_4__82_, fifo_data_o_4__81_, fifo_data_o_4__80_, fifo_data_o_4__79_, fifo_data_o_4__78_, fifo_data_o_4__77_, fifo_data_o_4__76_, fifo_data_o_4__75_, fifo_data_o_4__74_, fifo_data_o_4__73_, fifo_data_o_4__72_, fifo_data_o_4__71_, fifo_data_o_4__70_, fifo_data_o_4__69_, fifo_data_o_4__68_, fifo_data_o_4__67_, fifo_data_o_4__66_, fifo_data_o_4__65_, fifo_data_o_4__64_, fifo_data_o_4__63_, fifo_data_o_4__62_, fifo_data_o_4__61_, fifo_data_o_4__60_, fifo_data_o_4__59_, fifo_data_o_4__58_, fifo_data_o_4__57_, fifo_data_o_4__56_, fifo_data_o_4__55_, fifo_data_o_4__54_, fifo_data_o_4__53_, fifo_data_o_4__52_, fifo_data_o_4__51_, fifo_data_o_4__50_, fifo_data_o_4__49_, fifo_data_o_4__48_, fifo_data_o_4__47_, fifo_data_o_4__46_, fifo_data_o_4__45_, fifo_data_o_4__44_, fifo_data_o_4__43_, fifo_data_o_4__42_, fifo_data_o_4__41_, fifo_data_o_4__40_, fifo_data_o_4__39_, fifo_data_o_4__38_, fifo_data_o_4__37_, fifo_data_o_4__36_, fifo_data_o_4__35_, fifo_data_o_4__34_, fifo_data_o_4__33_, fifo_data_o_4__32_, fifo_data_o_4__31_, fifo_data_o_4__30_, fifo_data_o_4__29_, fifo_data_o_4__28_, fifo_data_o_4__27_, fifo_data_o_4__26_, fifo_data_o_4__25_, fifo_data_o_4__24_, fifo_data_o_4__23_, fifo_data_o_4__22_, fifo_data_o_4__21_, fifo_data_o_4__20_, fifo_data_o_4__19_, fifo_data_o_4__18_, fifo_data_o_4__17_, fifo_data_o_4__16_, fifo_data_o_4__15_, fifo_data_o_4__14_, fifo_data_o_4__13_, fifo_data_o_4__12_, fifo_data_o_4__11_, fifo_data_o_4__10_, fifo_data_o_4__9_, fifo_data_o_4__8_, fifo_data_o_4__7_, fifo_data_o_4__6_, fifo_data_o_4__5_, fifo_data_o_4__4_, fifo_data_o_4__3_, fifo_data_o_4__2_, fifo_data_o_4__1_, fifo_data_o_4__0_, fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_, fifo_data_o_2__130_, fifo_data_o_2__129_, fifo_data_o_2__128_, fifo_data_o_2__127_, fifo_data_o_2__126_, fifo_data_o_2__125_, fifo_data_o_2__124_, fifo_data_o_2__123_, fifo_data_o_2__122_, fifo_data_o_2__121_, fifo_data_o_2__120_, fifo_data_o_2__119_, fifo_data_o_2__118_, fifo_data_o_2__117_, fifo_data_o_2__116_, fifo_data_o_2__115_, fifo_data_o_2__114_, fifo_data_o_2__113_, fifo_data_o_2__112_, fifo_data_o_2__111_, fifo_data_o_2__110_, fifo_data_o_2__109_, fifo_data_o_2__108_, fifo_data_o_2__107_, fifo_data_o_2__106_, fifo_data_o_2__105_, fifo_data_o_2__104_, fifo_data_o_2__103_, fifo_data_o_2__102_, fifo_data_o_2__101_, fifo_data_o_2__100_, fifo_data_o_2__99_, fifo_data_o_2__98_, fifo_data_o_2__97_, fifo_data_o_2__96_, fifo_data_o_2__95_, fifo_data_o_2__94_, fifo_data_o_2__93_, fifo_data_o_2__92_, fifo_data_o_2__91_, fifo_data_o_2__90_, fifo_data_o_2__89_, fifo_data_o_2__88_, fifo_data_o_2__87_, fifo_data_o_2__86_, fifo_data_o_2__85_, fifo_data_o_2__84_, fifo_data_o_2__83_, fifo_data_o_2__82_, fifo_data_o_2__81_, fifo_data_o_2__80_, fifo_data_o_2__79_, fifo_data_o_2__78_, fifo_data_o_2__77_, fifo_data_o_2__76_, fifo_data_o_2__75_, fifo_data_o_2__74_, fifo_data_o_2__73_, fifo_data_o_2__72_, fifo_data_o_2__71_, fifo_data_o_2__70_, fifo_data_o_2__69_, fifo_data_o_2__68_, fifo_data_o_2__67_, fifo_data_o_2__66_, fifo_data_o_2__65_, fifo_data_o_2__64_, fifo_data_o_2__63_, fifo_data_o_2__62_, fifo_data_o_2__61_, fifo_data_o_2__60_, fifo_data_o_2__59_, fifo_data_o_2__58_, fifo_data_o_2__57_, fifo_data_o_2__56_, fifo_data_o_2__55_, fifo_data_o_2__54_, fifo_data_o_2__53_, fifo_data_o_2__52_, fifo_data_o_2__51_, fifo_data_o_2__50_, fifo_data_o_2__49_, fifo_data_o_2__48_, fifo_data_o_2__47_, fifo_data_o_2__46_, fifo_data_o_2__45_, fifo_data_o_2__44_, fifo_data_o_2__43_, fifo_data_o_2__42_, fifo_data_o_2__41_, fifo_data_o_2__40_, fifo_data_o_2__39_, fifo_data_o_2__38_, fifo_data_o_2__37_, fifo_data_o_2__36_, fifo_data_o_2__35_, fifo_data_o_2__34_, fifo_data_o_2__33_, fifo_data_o_2__32_, fifo_data_o_2__31_, fifo_data_o_2__30_, fifo_data_o_2__29_, fifo_data_o_2__28_, fifo_data_o_2__27_, fifo_data_o_2__26_, fifo_data_o_2__25_, fifo_data_o_2__24_, fifo_data_o_2__23_, fifo_data_o_2__22_, fifo_data_o_2__21_, fifo_data_o_2__20_, fifo_data_o_2__19_, fifo_data_o_2__18_, fifo_data_o_2__17_, fifo_data_o_2__16_, fifo_data_o_2__15_, fifo_data_o_2__14_, fifo_data_o_2__13_, fifo_data_o_2__12_, fifo_data_o_2__11_, fifo_data_o_2__10_, fifo_data_o_2__9_, fifo_data_o_2__8_, fifo_data_o_2__7_, fifo_data_o_2__6_, fifo_data_o_2__5_, fifo_data_o_2__4_, fifo_data_o_2__3_, fifo_data_o_2__2_, fifo_data_o_2__1_, fifo_data_o_2__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_1__3_, arb_sel_o_1__2_, arb_sel_o_1__1_, arb_sel_o_1__0_ }),
    .data_o(data_o[261:131])
  );


  bsg_round_robin_arb_inputs_p4
  out_side_2__rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[2]),
    .reqs_i({ arb_valid_4__2_, arb_valid_3__2_, arb_valid_1__2_, arb_valid_0__2_ }),
    .grants_o({ arb_grants_o_4__2_, arb_grants_o_3__2_, arb_grants_o_1__2_, arb_grants_o_0__2_ }),
    .sel_one_hot_o({ arb_sel_o_2__3_, arb_sel_o_2__2_, arb_sel_o_2__1_, arb_sel_o_2__0_ }),
    .v_o(valid_o[2]),
    .tag_o({ SV2V_UNCONNECTED_3, SV2V_UNCONNECTED_4 }),
    .yumi_i(n_9_net_)
  );


  bsg_mux_one_hot_width_p131_els_p4
  out_side_2__mux
  (
    .data_i({ fifo_data_o_4__130_, fifo_data_o_4__129_, fifo_data_o_4__128_, fifo_data_o_4__127_, fifo_data_o_4__126_, fifo_data_o_4__125_, fifo_data_o_4__124_, fifo_data_o_4__123_, fifo_data_o_4__122_, fifo_data_o_4__121_, fifo_data_o_4__120_, fifo_data_o_4__119_, fifo_data_o_4__118_, fifo_data_o_4__117_, fifo_data_o_4__116_, fifo_data_o_4__115_, fifo_data_o_4__114_, fifo_data_o_4__113_, fifo_data_o_4__112_, fifo_data_o_4__111_, fifo_data_o_4__110_, fifo_data_o_4__109_, fifo_data_o_4__108_, fifo_data_o_4__107_, fifo_data_o_4__106_, fifo_data_o_4__105_, fifo_data_o_4__104_, fifo_data_o_4__103_, fifo_data_o_4__102_, fifo_data_o_4__101_, fifo_data_o_4__100_, fifo_data_o_4__99_, fifo_data_o_4__98_, fifo_data_o_4__97_, fifo_data_o_4__96_, fifo_data_o_4__95_, fifo_data_o_4__94_, fifo_data_o_4__93_, fifo_data_o_4__92_, fifo_data_o_4__91_, fifo_data_o_4__90_, fifo_data_o_4__89_, fifo_data_o_4__88_, fifo_data_o_4__87_, fifo_data_o_4__86_, fifo_data_o_4__85_, fifo_data_o_4__84_, fifo_data_o_4__83_, fifo_data_o_4__82_, fifo_data_o_4__81_, fifo_data_o_4__80_, fifo_data_o_4__79_, fifo_data_o_4__78_, fifo_data_o_4__77_, fifo_data_o_4__76_, fifo_data_o_4__75_, fifo_data_o_4__74_, fifo_data_o_4__73_, fifo_data_o_4__72_, fifo_data_o_4__71_, fifo_data_o_4__70_, fifo_data_o_4__69_, fifo_data_o_4__68_, fifo_data_o_4__67_, fifo_data_o_4__66_, fifo_data_o_4__65_, fifo_data_o_4__64_, fifo_data_o_4__63_, fifo_data_o_4__62_, fifo_data_o_4__61_, fifo_data_o_4__60_, fifo_data_o_4__59_, fifo_data_o_4__58_, fifo_data_o_4__57_, fifo_data_o_4__56_, fifo_data_o_4__55_, fifo_data_o_4__54_, fifo_data_o_4__53_, fifo_data_o_4__52_, fifo_data_o_4__51_, fifo_data_o_4__50_, fifo_data_o_4__49_, fifo_data_o_4__48_, fifo_data_o_4__47_, fifo_data_o_4__46_, fifo_data_o_4__45_, fifo_data_o_4__44_, fifo_data_o_4__43_, fifo_data_o_4__42_, fifo_data_o_4__41_, fifo_data_o_4__40_, fifo_data_o_4__39_, fifo_data_o_4__38_, fifo_data_o_4__37_, fifo_data_o_4__36_, fifo_data_o_4__35_, fifo_data_o_4__34_, fifo_data_o_4__33_, fifo_data_o_4__32_, fifo_data_o_4__31_, fifo_data_o_4__30_, fifo_data_o_4__29_, fifo_data_o_4__28_, fifo_data_o_4__27_, fifo_data_o_4__26_, fifo_data_o_4__25_, fifo_data_o_4__24_, fifo_data_o_4__23_, fifo_data_o_4__22_, fifo_data_o_4__21_, fifo_data_o_4__20_, fifo_data_o_4__19_, fifo_data_o_4__18_, fifo_data_o_4__17_, fifo_data_o_4__16_, fifo_data_o_4__15_, fifo_data_o_4__14_, fifo_data_o_4__13_, fifo_data_o_4__12_, fifo_data_o_4__11_, fifo_data_o_4__10_, fifo_data_o_4__9_, fifo_data_o_4__8_, fifo_data_o_4__7_, fifo_data_o_4__6_, fifo_data_o_4__5_, fifo_data_o_4__4_, fifo_data_o_4__3_, fifo_data_o_4__2_, fifo_data_o_4__1_, fifo_data_o_4__0_, fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_2__3_, arb_sel_o_2__2_, arb_sel_o_2__1_, arb_sel_o_2__0_ }),
    .data_o(data_o[392:262])
  );


  bsg_round_robin_arb_inputs_p4
  out_side_3__rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ arb_valid_4__3_, arb_valid_2__3_, arb_valid_1__3_, arb_valid_0__3_ }),
    .grants_o({ arb_grants_o_4__3_, arb_grants_o_2__3_, arb_grants_o_1__3_, arb_grants_o_0__3_ }),
    .sel_one_hot_o({ arb_sel_o_3__3_, arb_sel_o_3__2_, arb_sel_o_3__1_, arb_sel_o_3__0_ }),
    .v_o(valid_o[3]),
    .tag_o({ SV2V_UNCONNECTED_5, SV2V_UNCONNECTED_6 }),
    .yumi_i(n_15_net_)
  );


  bsg_mux_one_hot_width_p131_els_p4
  out_side_3__mux
  (
    .data_i({ fifo_data_o_4__130_, fifo_data_o_4__129_, fifo_data_o_4__128_, fifo_data_o_4__127_, fifo_data_o_4__126_, fifo_data_o_4__125_, fifo_data_o_4__124_, fifo_data_o_4__123_, fifo_data_o_4__122_, fifo_data_o_4__121_, fifo_data_o_4__120_, fifo_data_o_4__119_, fifo_data_o_4__118_, fifo_data_o_4__117_, fifo_data_o_4__116_, fifo_data_o_4__115_, fifo_data_o_4__114_, fifo_data_o_4__113_, fifo_data_o_4__112_, fifo_data_o_4__111_, fifo_data_o_4__110_, fifo_data_o_4__109_, fifo_data_o_4__108_, fifo_data_o_4__107_, fifo_data_o_4__106_, fifo_data_o_4__105_, fifo_data_o_4__104_, fifo_data_o_4__103_, fifo_data_o_4__102_, fifo_data_o_4__101_, fifo_data_o_4__100_, fifo_data_o_4__99_, fifo_data_o_4__98_, fifo_data_o_4__97_, fifo_data_o_4__96_, fifo_data_o_4__95_, fifo_data_o_4__94_, fifo_data_o_4__93_, fifo_data_o_4__92_, fifo_data_o_4__91_, fifo_data_o_4__90_, fifo_data_o_4__89_, fifo_data_o_4__88_, fifo_data_o_4__87_, fifo_data_o_4__86_, fifo_data_o_4__85_, fifo_data_o_4__84_, fifo_data_o_4__83_, fifo_data_o_4__82_, fifo_data_o_4__81_, fifo_data_o_4__80_, fifo_data_o_4__79_, fifo_data_o_4__78_, fifo_data_o_4__77_, fifo_data_o_4__76_, fifo_data_o_4__75_, fifo_data_o_4__74_, fifo_data_o_4__73_, fifo_data_o_4__72_, fifo_data_o_4__71_, fifo_data_o_4__70_, fifo_data_o_4__69_, fifo_data_o_4__68_, fifo_data_o_4__67_, fifo_data_o_4__66_, fifo_data_o_4__65_, fifo_data_o_4__64_, fifo_data_o_4__63_, fifo_data_o_4__62_, fifo_data_o_4__61_, fifo_data_o_4__60_, fifo_data_o_4__59_, fifo_data_o_4__58_, fifo_data_o_4__57_, fifo_data_o_4__56_, fifo_data_o_4__55_, fifo_data_o_4__54_, fifo_data_o_4__53_, fifo_data_o_4__52_, fifo_data_o_4__51_, fifo_data_o_4__50_, fifo_data_o_4__49_, fifo_data_o_4__48_, fifo_data_o_4__47_, fifo_data_o_4__46_, fifo_data_o_4__45_, fifo_data_o_4__44_, fifo_data_o_4__43_, fifo_data_o_4__42_, fifo_data_o_4__41_, fifo_data_o_4__40_, fifo_data_o_4__39_, fifo_data_o_4__38_, fifo_data_o_4__37_, fifo_data_o_4__36_, fifo_data_o_4__35_, fifo_data_o_4__34_, fifo_data_o_4__33_, fifo_data_o_4__32_, fifo_data_o_4__31_, fifo_data_o_4__30_, fifo_data_o_4__29_, fifo_data_o_4__28_, fifo_data_o_4__27_, fifo_data_o_4__26_, fifo_data_o_4__25_, fifo_data_o_4__24_, fifo_data_o_4__23_, fifo_data_o_4__22_, fifo_data_o_4__21_, fifo_data_o_4__20_, fifo_data_o_4__19_, fifo_data_o_4__18_, fifo_data_o_4__17_, fifo_data_o_4__16_, fifo_data_o_4__15_, fifo_data_o_4__14_, fifo_data_o_4__13_, fifo_data_o_4__12_, fifo_data_o_4__11_, fifo_data_o_4__10_, fifo_data_o_4__9_, fifo_data_o_4__8_, fifo_data_o_4__7_, fifo_data_o_4__6_, fifo_data_o_4__5_, fifo_data_o_4__4_, fifo_data_o_4__3_, fifo_data_o_4__2_, fifo_data_o_4__1_, fifo_data_o_4__0_, fifo_data_o_2__130_, fifo_data_o_2__129_, fifo_data_o_2__128_, fifo_data_o_2__127_, fifo_data_o_2__126_, fifo_data_o_2__125_, fifo_data_o_2__124_, fifo_data_o_2__123_, fifo_data_o_2__122_, fifo_data_o_2__121_, fifo_data_o_2__120_, fifo_data_o_2__119_, fifo_data_o_2__118_, fifo_data_o_2__117_, fifo_data_o_2__116_, fifo_data_o_2__115_, fifo_data_o_2__114_, fifo_data_o_2__113_, fifo_data_o_2__112_, fifo_data_o_2__111_, fifo_data_o_2__110_, fifo_data_o_2__109_, fifo_data_o_2__108_, fifo_data_o_2__107_, fifo_data_o_2__106_, fifo_data_o_2__105_, fifo_data_o_2__104_, fifo_data_o_2__103_, fifo_data_o_2__102_, fifo_data_o_2__101_, fifo_data_o_2__100_, fifo_data_o_2__99_, fifo_data_o_2__98_, fifo_data_o_2__97_, fifo_data_o_2__96_, fifo_data_o_2__95_, fifo_data_o_2__94_, fifo_data_o_2__93_, fifo_data_o_2__92_, fifo_data_o_2__91_, fifo_data_o_2__90_, fifo_data_o_2__89_, fifo_data_o_2__88_, fifo_data_o_2__87_, fifo_data_o_2__86_, fifo_data_o_2__85_, fifo_data_o_2__84_, fifo_data_o_2__83_, fifo_data_o_2__82_, fifo_data_o_2__81_, fifo_data_o_2__80_, fifo_data_o_2__79_, fifo_data_o_2__78_, fifo_data_o_2__77_, fifo_data_o_2__76_, fifo_data_o_2__75_, fifo_data_o_2__74_, fifo_data_o_2__73_, fifo_data_o_2__72_, fifo_data_o_2__71_, fifo_data_o_2__70_, fifo_data_o_2__69_, fifo_data_o_2__68_, fifo_data_o_2__67_, fifo_data_o_2__66_, fifo_data_o_2__65_, fifo_data_o_2__64_, fifo_data_o_2__63_, fifo_data_o_2__62_, fifo_data_o_2__61_, fifo_data_o_2__60_, fifo_data_o_2__59_, fifo_data_o_2__58_, fifo_data_o_2__57_, fifo_data_o_2__56_, fifo_data_o_2__55_, fifo_data_o_2__54_, fifo_data_o_2__53_, fifo_data_o_2__52_, fifo_data_o_2__51_, fifo_data_o_2__50_, fifo_data_o_2__49_, fifo_data_o_2__48_, fifo_data_o_2__47_, fifo_data_o_2__46_, fifo_data_o_2__45_, fifo_data_o_2__44_, fifo_data_o_2__43_, fifo_data_o_2__42_, fifo_data_o_2__41_, fifo_data_o_2__40_, fifo_data_o_2__39_, fifo_data_o_2__38_, fifo_data_o_2__37_, fifo_data_o_2__36_, fifo_data_o_2__35_, fifo_data_o_2__34_, fifo_data_o_2__33_, fifo_data_o_2__32_, fifo_data_o_2__31_, fifo_data_o_2__30_, fifo_data_o_2__29_, fifo_data_o_2__28_, fifo_data_o_2__27_, fifo_data_o_2__26_, fifo_data_o_2__25_, fifo_data_o_2__24_, fifo_data_o_2__23_, fifo_data_o_2__22_, fifo_data_o_2__21_, fifo_data_o_2__20_, fifo_data_o_2__19_, fifo_data_o_2__18_, fifo_data_o_2__17_, fifo_data_o_2__16_, fifo_data_o_2__15_, fifo_data_o_2__14_, fifo_data_o_2__13_, fifo_data_o_2__12_, fifo_data_o_2__11_, fifo_data_o_2__10_, fifo_data_o_2__9_, fifo_data_o_2__8_, fifo_data_o_2__7_, fifo_data_o_2__6_, fifo_data_o_2__5_, fifo_data_o_2__4_, fifo_data_o_2__3_, fifo_data_o_2__2_, fifo_data_o_2__1_, fifo_data_o_2__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_3__3_, arb_sel_o_3__2_, arb_sel_o_3__1_, arb_sel_o_3__0_ }),
    .data_o(data_o[523:393])
  );


  bsg_round_robin_arb_inputs_p4
  out_side_4__rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ arb_valid_3__4_, arb_valid_2__4_, arb_valid_1__4_, arb_valid_0__4_ }),
    .grants_o({ arb_grants_o_3__4_, arb_grants_o_2__4_, arb_grants_o_1__4_, arb_grants_o_0__4_ }),
    .sel_one_hot_o({ arb_sel_o_4__3_, arb_sel_o_4__2_, arb_sel_o_4__1_, arb_sel_o_4__0_ }),
    .v_o(valid_o[4]),
    .tag_o({ SV2V_UNCONNECTED_7, SV2V_UNCONNECTED_8 }),
    .yumi_i(n_21_net_)
  );


  bsg_mux_one_hot_width_p131_els_p4
  out_side_4__mux
  (
    .data_i({ fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_, fifo_data_o_2__130_, fifo_data_o_2__129_, fifo_data_o_2__128_, fifo_data_o_2__127_, fifo_data_o_2__126_, fifo_data_o_2__125_, fifo_data_o_2__124_, fifo_data_o_2__123_, fifo_data_o_2__122_, fifo_data_o_2__121_, fifo_data_o_2__120_, fifo_data_o_2__119_, fifo_data_o_2__118_, fifo_data_o_2__117_, fifo_data_o_2__116_, fifo_data_o_2__115_, fifo_data_o_2__114_, fifo_data_o_2__113_, fifo_data_o_2__112_, fifo_data_o_2__111_, fifo_data_o_2__110_, fifo_data_o_2__109_, fifo_data_o_2__108_, fifo_data_o_2__107_, fifo_data_o_2__106_, fifo_data_o_2__105_, fifo_data_o_2__104_, fifo_data_o_2__103_, fifo_data_o_2__102_, fifo_data_o_2__101_, fifo_data_o_2__100_, fifo_data_o_2__99_, fifo_data_o_2__98_, fifo_data_o_2__97_, fifo_data_o_2__96_, fifo_data_o_2__95_, fifo_data_o_2__94_, fifo_data_o_2__93_, fifo_data_o_2__92_, fifo_data_o_2__91_, fifo_data_o_2__90_, fifo_data_o_2__89_, fifo_data_o_2__88_, fifo_data_o_2__87_, fifo_data_o_2__86_, fifo_data_o_2__85_, fifo_data_o_2__84_, fifo_data_o_2__83_, fifo_data_o_2__82_, fifo_data_o_2__81_, fifo_data_o_2__80_, fifo_data_o_2__79_, fifo_data_o_2__78_, fifo_data_o_2__77_, fifo_data_o_2__76_, fifo_data_o_2__75_, fifo_data_o_2__74_, fifo_data_o_2__73_, fifo_data_o_2__72_, fifo_data_o_2__71_, fifo_data_o_2__70_, fifo_data_o_2__69_, fifo_data_o_2__68_, fifo_data_o_2__67_, fifo_data_o_2__66_, fifo_data_o_2__65_, fifo_data_o_2__64_, fifo_data_o_2__63_, fifo_data_o_2__62_, fifo_data_o_2__61_, fifo_data_o_2__60_, fifo_data_o_2__59_, fifo_data_o_2__58_, fifo_data_o_2__57_, fifo_data_o_2__56_, fifo_data_o_2__55_, fifo_data_o_2__54_, fifo_data_o_2__53_, fifo_data_o_2__52_, fifo_data_o_2__51_, fifo_data_o_2__50_, fifo_data_o_2__49_, fifo_data_o_2__48_, fifo_data_o_2__47_, fifo_data_o_2__46_, fifo_data_o_2__45_, fifo_data_o_2__44_, fifo_data_o_2__43_, fifo_data_o_2__42_, fifo_data_o_2__41_, fifo_data_o_2__40_, fifo_data_o_2__39_, fifo_data_o_2__38_, fifo_data_o_2__37_, fifo_data_o_2__36_, fifo_data_o_2__35_, fifo_data_o_2__34_, fifo_data_o_2__33_, fifo_data_o_2__32_, fifo_data_o_2__31_, fifo_data_o_2__30_, fifo_data_o_2__29_, fifo_data_o_2__28_, fifo_data_o_2__27_, fifo_data_o_2__26_, fifo_data_o_2__25_, fifo_data_o_2__24_, fifo_data_o_2__23_, fifo_data_o_2__22_, fifo_data_o_2__21_, fifo_data_o_2__20_, fifo_data_o_2__19_, fifo_data_o_2__18_, fifo_data_o_2__17_, fifo_data_o_2__16_, fifo_data_o_2__15_, fifo_data_o_2__14_, fifo_data_o_2__13_, fifo_data_o_2__12_, fifo_data_o_2__11_, fifo_data_o_2__10_, fifo_data_o_2__9_, fifo_data_o_2__8_, fifo_data_o_2__7_, fifo_data_o_2__6_, fifo_data_o_2__5_, fifo_data_o_2__4_, fifo_data_o_2__3_, fifo_data_o_2__2_, fifo_data_o_2__1_, fifo_data_o_2__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_4__3_, arb_sel_o_4__2_, arb_sel_o_4__1_, arb_sel_o_4__0_ }),
    .data_o(data_o[654:524])
  );


  bsg_round_robin_arb_inputs_p5
  rr_arb_proc
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[0]),
    .reqs_i({ arb_valid_4__0_, arb_valid_3__0_, arb_valid_2__0_, arb_valid_1__0_, arb_valid_0__0_ }),
    .grants_o({ arb_grants_o_4__0_, arb_grants_o_3__0_, arb_grants_o_2__0_, arb_grants_o_1__0_, arb_grants_o_0__0_ }),
    .sel_one_hot_o({ arb_sel_o_0__4_, arb_sel_o_0__3_, arb_sel_o_0__2_, arb_sel_o_0__1_, arb_sel_o_0__0_ }),
    .v_o(valid_o[0]),
    .tag_o({ SV2V_UNCONNECTED_9, SV2V_UNCONNECTED_10, SV2V_UNCONNECTED_11 }),
    .yumi_i(n_27_net_)
  );


  bsg_mux_one_hot_width_p131_els_p5
  mux_proc
  (
    .data_i({ fifo_data_o_4__130_, fifo_data_o_4__129_, fifo_data_o_4__128_, fifo_data_o_4__127_, fifo_data_o_4__126_, fifo_data_o_4__125_, fifo_data_o_4__124_, fifo_data_o_4__123_, fifo_data_o_4__122_, fifo_data_o_4__121_, fifo_data_o_4__120_, fifo_data_o_4__119_, fifo_data_o_4__118_, fifo_data_o_4__117_, fifo_data_o_4__116_, fifo_data_o_4__115_, fifo_data_o_4__114_, fifo_data_o_4__113_, fifo_data_o_4__112_, fifo_data_o_4__111_, fifo_data_o_4__110_, fifo_data_o_4__109_, fifo_data_o_4__108_, fifo_data_o_4__107_, fifo_data_o_4__106_, fifo_data_o_4__105_, fifo_data_o_4__104_, fifo_data_o_4__103_, fifo_data_o_4__102_, fifo_data_o_4__101_, fifo_data_o_4__100_, fifo_data_o_4__99_, fifo_data_o_4__98_, fifo_data_o_4__97_, fifo_data_o_4__96_, fifo_data_o_4__95_, fifo_data_o_4__94_, fifo_data_o_4__93_, fifo_data_o_4__92_, fifo_data_o_4__91_, fifo_data_o_4__90_, fifo_data_o_4__89_, fifo_data_o_4__88_, fifo_data_o_4__87_, fifo_data_o_4__86_, fifo_data_o_4__85_, fifo_data_o_4__84_, fifo_data_o_4__83_, fifo_data_o_4__82_, fifo_data_o_4__81_, fifo_data_o_4__80_, fifo_data_o_4__79_, fifo_data_o_4__78_, fifo_data_o_4__77_, fifo_data_o_4__76_, fifo_data_o_4__75_, fifo_data_o_4__74_, fifo_data_o_4__73_, fifo_data_o_4__72_, fifo_data_o_4__71_, fifo_data_o_4__70_, fifo_data_o_4__69_, fifo_data_o_4__68_, fifo_data_o_4__67_, fifo_data_o_4__66_, fifo_data_o_4__65_, fifo_data_o_4__64_, fifo_data_o_4__63_, fifo_data_o_4__62_, fifo_data_o_4__61_, fifo_data_o_4__60_, fifo_data_o_4__59_, fifo_data_o_4__58_, fifo_data_o_4__57_, fifo_data_o_4__56_, fifo_data_o_4__55_, fifo_data_o_4__54_, fifo_data_o_4__53_, fifo_data_o_4__52_, fifo_data_o_4__51_, fifo_data_o_4__50_, fifo_data_o_4__49_, fifo_data_o_4__48_, fifo_data_o_4__47_, fifo_data_o_4__46_, fifo_data_o_4__45_, fifo_data_o_4__44_, fifo_data_o_4__43_, fifo_data_o_4__42_, fifo_data_o_4__41_, fifo_data_o_4__40_, fifo_data_o_4__39_, fifo_data_o_4__38_, fifo_data_o_4__37_, fifo_data_o_4__36_, fifo_data_o_4__35_, fifo_data_o_4__34_, fifo_data_o_4__33_, fifo_data_o_4__32_, fifo_data_o_4__31_, fifo_data_o_4__30_, fifo_data_o_4__29_, fifo_data_o_4__28_, fifo_data_o_4__27_, fifo_data_o_4__26_, fifo_data_o_4__25_, fifo_data_o_4__24_, fifo_data_o_4__23_, fifo_data_o_4__22_, fifo_data_o_4__21_, fifo_data_o_4__20_, fifo_data_o_4__19_, fifo_data_o_4__18_, fifo_data_o_4__17_, fifo_data_o_4__16_, fifo_data_o_4__15_, fifo_data_o_4__14_, fifo_data_o_4__13_, fifo_data_o_4__12_, fifo_data_o_4__11_, fifo_data_o_4__10_, fifo_data_o_4__9_, fifo_data_o_4__8_, fifo_data_o_4__7_, fifo_data_o_4__6_, fifo_data_o_4__5_, fifo_data_o_4__4_, fifo_data_o_4__3_, fifo_data_o_4__2_, fifo_data_o_4__1_, fifo_data_o_4__0_, fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_, fifo_data_o_2__130_, fifo_data_o_2__129_, fifo_data_o_2__128_, fifo_data_o_2__127_, fifo_data_o_2__126_, fifo_data_o_2__125_, fifo_data_o_2__124_, fifo_data_o_2__123_, fifo_data_o_2__122_, fifo_data_o_2__121_, fifo_data_o_2__120_, fifo_data_o_2__119_, fifo_data_o_2__118_, fifo_data_o_2__117_, fifo_data_o_2__116_, fifo_data_o_2__115_, fifo_data_o_2__114_, fifo_data_o_2__113_, fifo_data_o_2__112_, fifo_data_o_2__111_, fifo_data_o_2__110_, fifo_data_o_2__109_, fifo_data_o_2__108_, fifo_data_o_2__107_, fifo_data_o_2__106_, fifo_data_o_2__105_, fifo_data_o_2__104_, fifo_data_o_2__103_, fifo_data_o_2__102_, fifo_data_o_2__101_, fifo_data_o_2__100_, fifo_data_o_2__99_, fifo_data_o_2__98_, fifo_data_o_2__97_, fifo_data_o_2__96_, fifo_data_o_2__95_, fifo_data_o_2__94_, fifo_data_o_2__93_, fifo_data_o_2__92_, fifo_data_o_2__91_, fifo_data_o_2__90_, fifo_data_o_2__89_, fifo_data_o_2__88_, fifo_data_o_2__87_, fifo_data_o_2__86_, fifo_data_o_2__85_, fifo_data_o_2__84_, fifo_data_o_2__83_, fifo_data_o_2__82_, fifo_data_o_2__81_, fifo_data_o_2__80_, fifo_data_o_2__79_, fifo_data_o_2__78_, fifo_data_o_2__77_, fifo_data_o_2__76_, fifo_data_o_2__75_, fifo_data_o_2__74_, fifo_data_o_2__73_, fifo_data_o_2__72_, fifo_data_o_2__71_, fifo_data_o_2__70_, fifo_data_o_2__69_, fifo_data_o_2__68_, fifo_data_o_2__67_, fifo_data_o_2__66_, fifo_data_o_2__65_, fifo_data_o_2__64_, fifo_data_o_2__63_, fifo_data_o_2__62_, fifo_data_o_2__61_, fifo_data_o_2__60_, fifo_data_o_2__59_, fifo_data_o_2__58_, fifo_data_o_2__57_, fifo_data_o_2__56_, fifo_data_o_2__55_, fifo_data_o_2__54_, fifo_data_o_2__53_, fifo_data_o_2__52_, fifo_data_o_2__51_, fifo_data_o_2__50_, fifo_data_o_2__49_, fifo_data_o_2__48_, fifo_data_o_2__47_, fifo_data_o_2__46_, fifo_data_o_2__45_, fifo_data_o_2__44_, fifo_data_o_2__43_, fifo_data_o_2__42_, fifo_data_o_2__41_, fifo_data_o_2__40_, fifo_data_o_2__39_, fifo_data_o_2__38_, fifo_data_o_2__37_, fifo_data_o_2__36_, fifo_data_o_2__35_, fifo_data_o_2__34_, fifo_data_o_2__33_, fifo_data_o_2__32_, fifo_data_o_2__31_, fifo_data_o_2__30_, fifo_data_o_2__29_, fifo_data_o_2__28_, fifo_data_o_2__27_, fifo_data_o_2__26_, fifo_data_o_2__25_, fifo_data_o_2__24_, fifo_data_o_2__23_, fifo_data_o_2__22_, fifo_data_o_2__21_, fifo_data_o_2__20_, fifo_data_o_2__19_, fifo_data_o_2__18_, fifo_data_o_2__17_, fifo_data_o_2__16_, fifo_data_o_2__15_, fifo_data_o_2__14_, fifo_data_o_2__13_, fifo_data_o_2__12_, fifo_data_o_2__11_, fifo_data_o_2__10_, fifo_data_o_2__9_, fifo_data_o_2__8_, fifo_data_o_2__7_, fifo_data_o_2__6_, fifo_data_o_2__5_, fifo_data_o_2__4_, fifo_data_o_2__3_, fifo_data_o_2__2_, fifo_data_o_2__1_, fifo_data_o_2__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_0__4_, arb_sel_o_0__3_, arb_sel_o_0__2_, arb_sel_o_0__1_, arb_sel_o_0__0_ }),
    .data_o(data_o[130:0])
  );

  assign N285 = N0 & local_x_cord_i[0];
  assign N0 = ~1'b0;
  assign N286 = 1'b0 & N1;
  assign N1 = ~local_x_cord_i[0];
  assign N290 = N2 & local_y_cord_i[0];
  assign N2 = ~1'b0;
  assign N291 = 1'b0 & N3;
  assign N3 = ~local_y_cord_i[0];
  assign N4 = fifo_data_o_2__1_ ^ local_y_cord_i[0];
  assign N292 = ~N4;
  assign N5 = fifo_data_o_2__0_ ^ local_x_cord_i[0];
  assign N294 = ~N5;
  assign N295 = N6 & local_x_cord_i[0];
  assign N6 = ~fifo_data_o_2__0_;
  assign N298 = N7 & local_y_cord_i[0];
  assign N7 = ~fifo_data_o_2__1_;
  assign N299 = fifo_data_o_2__1_ & N8;
  assign N8 = ~local_y_cord_i[0];
  assign N9 = fifo_data_o_3__1_ ^ local_y_cord_i[0];
  assign N300 = ~N9;
  assign N10 = fifo_data_o_3__0_ ^ local_x_cord_i[0];
  assign N302 = ~N10;
  assign N303 = N11 & local_x_cord_i[0];
  assign N11 = ~fifo_data_o_3__0_;
  assign N304 = fifo_data_o_3__0_ & N12;
  assign N12 = ~local_x_cord_i[0];
  assign N308 = fifo_data_o_3__1_ & N13;
  assign N13 = ~local_y_cord_i[0];
  assign N14 = fifo_data_o_4__1_ ^ local_y_cord_i[0];
  assign N309 = ~N14;
  assign N15 = fifo_data_o_4__0_ ^ local_x_cord_i[0];
  assign N311 = ~N15;
  assign N312 = N16 & local_x_cord_i[0];
  assign N16 = ~fifo_data_o_4__0_;
  assign N313 = fifo_data_o_4__0_ & N17;
  assign N17 = ~local_x_cord_i[0];
  assign N317 = N18 & local_y_cord_i[0];
  assign N18 = ~fifo_data_o_4__1_;
  assign N339 = out_count_r[2] | out_count_r[3];
  assign N340 = ~N339;
  assign N341 = out_count_r[2] | out_count_r[3];
  assign N342 = ~N341;
  assign N343 = out_count_r[2] | out_count_r[3];
  assign N344 = ~N343;
  assign N345 = out_count_r[2] | out_count_r[3];
  assign N346 = ~N345;
  assign N347 = out_count_r[4] | out_count_r[5];
  assign N348 = ~N347;
  assign N349 = out_count_r[4] | out_count_r[5];
  assign N350 = ~N349;
  assign N351 = out_count_r[4] | out_count_r[5];
  assign N352 = ~N351;
  assign N353 = out_count_r[4] | out_count_r[5];
  assign N354 = ~N353;
  assign N355 = out_count_r[6] | out_count_r[7];
  assign N356 = ~N355;
  assign N357 = out_count_r[6] | out_count_r[7];
  assign N358 = ~N357;
  assign N359 = out_count_r[6] | out_count_r[7];
  assign N360 = ~N359;
  assign N361 = out_count_r[6] | out_count_r[7];
  assign N362 = ~N361;
  assign N363 = out_count_r[8] | out_count_r[9];
  assign N364 = ~N363;
  assign N365 = out_count_r[8] | out_count_r[9];
  assign N366 = ~N365;
  assign N367 = out_count_r[8] | out_count_r[9];
  assign N368 = ~N367;
  assign N369 = out_count_r[8] | out_count_r[9];
  assign N370 = ~N369;
  assign N371 = out_count_r[0] | out_count_r[1];
  assign N372 = ~N371;
  assign N373 = out_count_r[0] | out_count_r[1];
  assign N374 = ~N373;
  assign N375 = out_count_r[0] | out_count_r[1];
  assign N376 = ~N375;
  assign N377 = out_count_r[0] | out_count_r[1];
  assign N378 = ~N377;
  assign N379 = out_count_r[0] | out_count_r[1];
  assign N380 = ~N379;
  assign N381 = out_count_r[0] | out_count_r[1];
  assign N382 = out_count_r[2] | out_count_r[3];
  assign N383 = out_count_r[4] | out_count_r[5];
  assign N384 = out_count_r[6] | out_count_r[7];
  assign N385 = out_count_r[8] | out_count_r[9];
  assign N386 = out_count_r[0] | out_count_r[1];
  assign N387 = out_count_r[4] | out_count_r[5];
  assign N388 = out_count_r[6] | out_count_r[7];
  assign N389 = out_count_r[8] | out_count_r[9];
  assign N390 = out_count_r[0] | out_count_r[1];
  assign N391 = out_count_r[2] | out_count_r[3];
  assign N392 = out_count_r[6] | out_count_r[7];
  assign N393 = out_count_r[8] | out_count_r[9];
  assign N394 = out_count_r[0] | out_count_r[1];
  assign N395 = out_count_r[2] | out_count_r[3];
  assign N396 = out_count_r[4] | out_count_r[5];
  assign N397 = out_count_r[8] | out_count_r[9];
  assign N398 = out_count_r[0] | out_count_r[1];
  assign N399 = out_count_r[2] | out_count_r[3];
  assign N400 = out_count_r[4] | out_count_r[5];
  assign N401 = out_count_r[6] | out_count_r[7];
  assign N402 = count_r[8] | count_r[9];
  assign N403 = ~N402;
  assign N404 = count_r[6] | count_r[7];
  assign N405 = ~N404;
  assign N406 = count_r[4] | count_r[5];
  assign N407 = ~N406;
  assign N408 = count_r[2] | count_r[3];
  assign N409 = ~N408;
  assign N410 = count_r[0] | count_r[1];
  assign N411 = ~N410;
  assign N412 = ~local_y_cord_i[0];
  assign N413 = ~local_x_cord_i[0];
  assign N414 = count_r[0] | count_r[1];
  assign N415 = ~N414;
  assign N416 = count_r[2] | count_r[3];
  assign N417 = ~N416;
  assign N418 = count_r[4] | count_r[5];
  assign N419 = ~N418;
  assign N420 = count_r[6] | count_r[7];
  assign N421 = ~N420;
  assign N422 = count_r[8] | count_r[9];
  assign N423 = ~N422;
  assign N424 = out_count_r[0] | out_count_r[1];
  assign N425 = ~N424;
  assign N426 = out_count_r[2] | out_count_r[3];
  assign N427 = ~N426;
  assign N428 = out_count_r[4] | out_count_r[5];
  assign N429 = ~N428;
  assign N430 = out_count_r[6] | out_count_r[7];
  assign N431 = ~N430;
  assign N432 = out_count_r[8] | out_count_r[9];
  assign N433 = ~N432;
  assign { N132, N131 } = count_r[1:0] - 1'b1;
  assign { N145, N144 } = count_r[3:2] - 1'b1;
  assign { N159, N158 } = count_r[5:4] - 1'b1;
  assign { N173, N172 } = count_r[7:6] - 1'b1;
  assign { N187, N186 } = count_r[9:8] - 1'b1;
  assign { N201, N200 } = out_count_r[1:0] - 1'b1;
  assign { N215, N214 } = out_count_r[3:2] - 1'b1;
  assign { N229, N228 } = out_count_r[5:4] - 1'b1;
  assign { N243, N242 } = out_count_r[7:6] - 1'b1;
  assign { N257, N256 } = out_count_r[9:8] - 1'b1;
  assign { N134, N133 } = (N19)? { 1'b0, 1'b0 } :
                          (N20)? { N132, N131 } : 1'b0;
  assign N19 = N415;
  assign N20 = N414;
  assign { N136, N135 } = (N21)? { N134, N133 } :
                          (N129)? count_r[1:0] : 1'b0;
  assign N21 = fifo_yumi_i[0];
  assign { N138, N137 } = (N22)? { 1'b0, 1'b0 } :
                          (N23)? { N136, N135 } : 1'b0;
  assign N22 = N127;
  assign N23 = N126;
  assign { N147, N146 } = (N24)? { 1'b0, 1'b0 } :
                          (N25)? { N145, N144 } : 1'b0;
  assign N24 = N417;
  assign N25 = N416;
  assign { N149, N148 } = (N26)? { N147, N146 } :
                          (N142)? count_r[3:2] : 1'b0;
  assign N26 = fifo_yumi_i[1];
  assign { N151, N150 } = (N27)? { 1'b0, 1'b0 } :
                          (N28)? { N149, N148 } : 1'b0;
  assign N27 = N140;
  assign N28 = N139;
  assign { N161, N160 } = (N29)? { fifo_data_o_2__3_, fifo_data_o_2__2_ } :
                          (N30)? { N159, N158 } : 1'b0;
  assign N29 = N419;
  assign N30 = N418;
  assign { N163, N162 } = (N31)? { N161, N160 } :
                          (N156)? count_r[5:4] : 1'b0;
  assign N31 = N155;
  assign { N165, N164 } = (N32)? { 1'b0, 1'b0 } :
                          (N33)? { N163, N162 } : 1'b0;
  assign N32 = N153;
  assign N33 = N152;
  assign { N175, N174 } = (N34)? { fifo_data_o_3__3_, fifo_data_o_3__2_ } :
                          (N35)? { N173, N172 } : 1'b0;
  assign N34 = N421;
  assign N35 = N420;
  assign { N177, N176 } = (N36)? { N175, N174 } :
                          (N170)? count_r[7:6] : 1'b0;
  assign N36 = N169;
  assign { N179, N178 } = (N37)? { 1'b0, 1'b0 } :
                          (N38)? { N177, N176 } : 1'b0;
  assign N37 = N167;
  assign N38 = N166;
  assign { N189, N188 } = (N39)? { fifo_data_o_4__3_, fifo_data_o_4__2_ } :
                          (N40)? { N187, N186 } : 1'b0;
  assign N39 = N423;
  assign N40 = N422;
  assign { N191, N190 } = (N41)? { N189, N188 } :
                          (N184)? count_r[9:8] : 1'b0;
  assign N41 = N183;
  assign { N193, N192 } = (N42)? { 1'b0, 1'b0 } :
                          (N43)? { N191, N190 } : 1'b0;
  assign N42 = N181;
  assign N43 = N180;
  assign { N203, N202 } = (N44)? data_o[3:2] :
                          (N45)? { N201, N200 } : 1'b0;
  assign N44 = N425;
  assign N45 = N424;
  assign { N205, N204 } = (N46)? { N203, N202 } :
                          (N198)? out_count_r[1:0] : 1'b0;
  assign N46 = N197;
  assign { N207, N206 } = (N47)? { 1'b0, 1'b0 } :
                          (N48)? { N205, N204 } : 1'b0;
  assign N47 = N195;
  assign N48 = N194;
  assign { N217, N216 } = (N49)? data_o[134:133] :
                          (N50)? { N215, N214 } : 1'b0;
  assign N49 = N427;
  assign N50 = N426;
  assign { N219, N218 } = (N51)? { N217, N216 } :
                          (N212)? out_count_r[3:2] : 1'b0;
  assign N51 = N211;
  assign { N221, N220 } = (N52)? { 1'b0, 1'b0 } :
                          (N53)? { N219, N218 } : 1'b0;
  assign N52 = N209;
  assign N53 = N208;
  assign { N231, N230 } = (N54)? data_o[265:264] :
                          (N55)? { N229, N228 } : 1'b0;
  assign N54 = N429;
  assign N55 = N428;
  assign { N233, N232 } = (N56)? { N231, N230 } :
                          (N226)? out_count_r[5:4] : 1'b0;
  assign N56 = N225;
  assign { N235, N234 } = (N57)? { 1'b0, 1'b0 } :
                          (N58)? { N233, N232 } : 1'b0;
  assign N57 = N223;
  assign N58 = N222;
  assign { N245, N244 } = (N59)? data_o[396:395] :
                          (N60)? { N243, N242 } : 1'b0;
  assign N59 = N431;
  assign N60 = N430;
  assign { N247, N246 } = (N61)? { N245, N244 } :
                          (N240)? out_count_r[7:6] : 1'b0;
  assign N61 = N239;
  assign { N249, N248 } = (N62)? { 1'b0, 1'b0 } :
                          (N63)? { N247, N246 } : 1'b0;
  assign N62 = N237;
  assign N63 = N236;
  assign { N259, N258 } = (N64)? data_o[527:526] :
                          (N65)? { N257, N256 } : 1'b0;
  assign N64 = N433;
  assign N65 = N432;
  assign { N261, N260 } = (N66)? { N259, N258 } :
                          (N254)? out_count_r[9:8] : 1'b0;
  assign N66 = N253;
  assign { N263, N262 } = (N67)? { 1'b0, 1'b0 } :
                          (N68)? { N261, N260 } : 1'b0;
  assign N67 = N251;
  assign N68 = N250;
  assign arb_valid_0__0_ = (N69)? new_valid_0__0_ :
                           (N70)? N264 : 1'b0;
  assign N69 = N380;
  assign N70 = N379;
  assign arb_valid_0__1_ = (N71)? new_valid_0__1_ :
                           (N72)? N265 : 1'b0;
  assign N71 = N346;
  assign N72 = N345;
  assign arb_valid_0__2_ = (N73)? new_valid_0__2_ :
                           (N74)? N266 : 1'b0;
  assign N73 = N354;
  assign N74 = N353;
  assign arb_valid_0__3_ = (N75)? new_valid_0__3_ :
                           (N76)? N267 : 1'b0;
  assign N75 = N362;
  assign N76 = N361;
  assign arb_valid_0__4_ = (N77)? new_valid_0__4_ :
                           (N78)? N268 : 1'b0;
  assign N77 = N370;
  assign N78 = N369;
  assign arb_valid_1__0_ = (N79)? new_valid_1__0_ :
                           (N80)? N269 : 1'b0;
  assign N79 = N378;
  assign N80 = N377;
  assign arb_valid_1__2_ = (N81)? new_valid_1__2_ :
                           (N82)? N270 : 1'b0;
  assign N81 = N352;
  assign N82 = N351;
  assign arb_valid_1__3_ = (N83)? new_valid_1__3_ :
                           (N84)? N271 : 1'b0;
  assign N83 = N360;
  assign N84 = N359;
  assign arb_valid_1__4_ = (N85)? new_valid_1__4_ :
                           (N86)? N272 : 1'b0;
  assign N85 = N368;
  assign N86 = N367;
  assign arb_valid_2__0_ = (N87)? new_valid_2__0_ :
                           (N88)? N273 : 1'b0;
  assign N87 = N376;
  assign N88 = N375;
  assign arb_valid_2__1_ = (N89)? new_valid_2__1_ :
                           (N90)? N274 : 1'b0;
  assign N89 = N344;
  assign N90 = N343;
  assign arb_valid_2__3_ = (N91)? new_valid_2__3_ :
                           (N92)? N275 : 1'b0;
  assign N91 = N358;
  assign N92 = N357;
  assign arb_valid_2__4_ = (N93)? new_valid_2__4_ :
                           (N94)? N276 : 1'b0;
  assign N93 = N366;
  assign N94 = N365;
  assign arb_valid_3__0_ = (N95)? new_valid_3__0_ :
                           (N96)? N277 : 1'b0;
  assign N95 = N374;
  assign N96 = N373;
  assign arb_valid_3__1_ = (N97)? new_valid_3__1_ :
                           (N98)? N278 : 1'b0;
  assign N97 = N342;
  assign N98 = N341;
  assign arb_valid_3__2_ = (N99)? new_valid_3__2_ :
                           (N100)? N279 : 1'b0;
  assign N99 = N350;
  assign N100 = N349;
  assign arb_valid_3__4_ = (N101)? new_valid_3__4_ :
                           (N102)? N280 : 1'b0;
  assign N101 = N364;
  assign N102 = N363;
  assign arb_valid_4__0_ = (N103)? new_valid_4__0_ :
                           (N104)? N281 : 1'b0;
  assign N103 = N372;
  assign N104 = N371;
  assign arb_valid_4__1_ = (N105)? new_valid_4__1_ :
                           (N106)? N282 : 1'b0;
  assign N105 = N340;
  assign N106 = N339;
  assign arb_valid_4__2_ = (N107)? new_valid_4__2_ :
                           (N108)? N283 : 1'b0;
  assign N107 = N348;
  assign N108 = N347;
  assign arb_valid_4__3_ = (N109)? new_valid_4__3_ :
                           (N110)? N284 : 1'b0;
  assign N109 = N356;
  assign N110 = N355;
  assign { N289, N288, N287 } = (N111)? { N286, N285, N413 } :
                                (N112)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N111 = N412;
  assign N112 = local_y_cord_i[0];
  assign { dest_n_0__4_, dest_n_0__3_, dest_n_0__2_, dest_n_0__1_, dest_n_0__0_ } = (N113)? { N291, N290, N289, N288, N287 } :
                                                                                    (N114)? { dest_r_0__4_, dest_r_0__3_, dest_r_0__2_, dest_r_0__1_, dest_r_0__0_ } : 1'b0;
  assign N113 = N411;
  assign N114 = N410;
  assign { dest_n_1__4_, dest_n_1__3_, dest_n_1__2_, dest_n_1__0_ } = (N115)? { N291, N290, N289, N287 } :
                                                                      (N116)? { dest_r_1__4_, dest_r_1__3_, dest_r_1__2_, dest_r_1__0_ } : 1'b0;
  assign N115 = N409;
  assign N116 = N408;
  assign { N297, N296 } = (N117)? { N295, N294 } :
                          (N293)? { 1'b0, 1'b0 } : 1'b0;
  assign N117 = N292;
  assign { dest_n_2__4_, dest_n_2__3_, dest_n_2__1_, dest_n_2__0_ } = (N118)? { N299, N298, N297, N296 } :
                                                                      (N119)? { dest_r_2__4_, dest_r_2__3_, dest_r_2__1_, dest_r_2__0_ } : 1'b0;
  assign N118 = N407;
  assign N119 = N406;
  assign { N307, N306, N305 } = (N120)? { N304, N303, N302 } :
                                (N301)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N120 = N300;
  assign { dest_n_3__4_, dest_n_3__2_, dest_n_3__1_, dest_n_3__0_ } = (N121)? { N308, N307, N306, N305 } :
                                                                      (N122)? { dest_r_3__4_, dest_r_3__2_, dest_r_3__1_, dest_r_3__0_ } : 1'b0;
  assign N121 = N405;
  assign N122 = N404;
  assign { N316, N315, N314 } = (N123)? { N313, N312, N311 } :
                                (N310)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N123 = N309;
  assign { dest_n_4__3_, dest_n_4__2_, dest_n_4__1_, dest_n_4__0_ } = (N124)? { N317, N316, N315, N314 } :
                                                                      (N125)? { dest_r_4__3_, dest_r_4__2_, dest_r_4__1_, dest_r_4__0_ } : 1'b0;
  assign N124 = N403;
  assign N125 = N402;
  assign N126 = ~reset_i;
  assign N127 = reset_i;
  assign N128 = N126;
  assign N129 = ~fifo_yumi_i[0];
  assign N130 = N128 & fifo_yumi_i[0];
  assign N139 = ~reset_i;
  assign N140 = reset_i;
  assign N141 = N139;
  assign N142 = ~fifo_yumi_i[1];
  assign N143 = N141 & fifo_yumi_i[1];
  assign N152 = ~reset_i;
  assign N153 = reset_i;
  assign N154 = N152;
  assign N155 = fifo_yumi_i[2];
  assign N156 = ~N155;
  assign N157 = N154 & N155;
  assign N166 = ~reset_i;
  assign N167 = reset_i;
  assign N168 = N166;
  assign N169 = fifo_yumi_i[3];
  assign N170 = ~N169;
  assign N171 = N168 & N169;
  assign N180 = ~reset_i;
  assign N181 = reset_i;
  assign N182 = N180;
  assign N183 = fifo_yumi_i[4];
  assign N184 = ~N183;
  assign N185 = N182 & N183;
  assign new_valid_0__0_ = 1'b0 & dest_n_0__0_;
  assign new_valid_0__1_ = 1'b0 & dest_n_0__1_;
  assign new_valid_0__2_ = 1'b0 & dest_n_0__2_;
  assign new_valid_0__3_ = 1'b0 & dest_n_0__3_;
  assign new_valid_0__4_ = 1'b0 & dest_n_0__4_;
  assign new_valid_1__0_ = 1'b0 & dest_n_1__0_;
  assign new_valid_1__2_ = 1'b0 & dest_n_1__2_;
  assign new_valid_1__3_ = 1'b0 & dest_n_1__3_;
  assign new_valid_1__4_ = 1'b0 & dest_n_1__4_;
  assign new_valid_2__0_ = fifo_valid_o[2] & dest_n_2__0_;
  assign new_valid_2__1_ = fifo_valid_o[2] & dest_n_2__1_;
  assign new_valid_2__3_ = fifo_valid_o[2] & dest_n_2__3_;
  assign new_valid_2__4_ = fifo_valid_o[2] & dest_n_2__4_;
  assign new_valid_3__0_ = fifo_valid_o[3] & dest_n_3__0_;
  assign new_valid_3__1_ = fifo_valid_o[3] & dest_n_3__1_;
  assign new_valid_3__2_ = fifo_valid_o[3] & dest_n_3__2_;
  assign new_valid_3__4_ = fifo_valid_o[3] & dest_n_3__4_;
  assign new_valid_4__0_ = fifo_valid_o[4] & dest_n_4__0_;
  assign new_valid_4__1_ = fifo_valid_o[4] & dest_n_4__1_;
  assign new_valid_4__2_ = fifo_valid_o[4] & dest_n_4__2_;
  assign new_valid_4__3_ = fifo_valid_o[4] & dest_n_4__3_;
  assign fifo_yumi_i[0] = N436 | arb_grants_o_0__0_;
  assign N436 = N435 | arb_grants_o_0__1_;
  assign N435 = N434 | arb_grants_o_0__2_;
  assign N434 = arb_grants_o_0__4_ | arb_grants_o_0__3_;
  assign fifo_yumi_i[1] = N439 | arb_grants_o_1__0_;
  assign N439 = N438 | 1'b0;
  assign N438 = N437 | arb_grants_o_1__2_;
  assign N437 = arb_grants_o_1__4_ | arb_grants_o_1__3_;
  assign fifo_yumi_i[2] = N442 | arb_grants_o_2__0_;
  assign N442 = N441 | arb_grants_o_2__1_;
  assign N441 = N440 | 1'b0;
  assign N440 = arb_grants_o_2__4_ | arb_grants_o_2__3_;
  assign fifo_yumi_i[3] = N445 | arb_grants_o_3__0_;
  assign N445 = N444 | arb_grants_o_3__1_;
  assign N444 = N443 | arb_grants_o_3__2_;
  assign N443 = arb_grants_o_3__4_ | 1'b0;
  assign fifo_yumi_i[4] = N448 | arb_grants_o_4__0_;
  assign N448 = N447 | arb_grants_o_4__1_;
  assign N447 = N446 | arb_grants_o_4__2_;
  assign N446 = 1'b0 | arb_grants_o_4__3_;
  assign N194 = ~reset_i;
  assign N195 = reset_i;
  assign N196 = N194;
  assign N197 = valid_o[0] & ready_i[0];
  assign N198 = ~N197;
  assign N199 = N196 & N197;
  assign N208 = ~reset_i;
  assign N209 = reset_i;
  assign N210 = N208;
  assign N211 = valid_o[1] & 1'b1;
  assign N212 = ~N211;
  assign N213 = N210 & N211;
  assign N222 = ~reset_i;
  assign N223 = reset_i;
  assign N224 = N222;
  assign N225 = valid_o[2] & ready_i[2];
  assign N226 = ~N225;
  assign N227 = N224 & N225;
  assign N236 = ~reset_i;
  assign N237 = reset_i;
  assign N238 = N236;
  assign N239 = valid_o[3] & 1'b1;
  assign N240 = ~N239;
  assign N241 = N238 & N239;
  assign N250 = ~reset_i;
  assign N251 = reset_i;
  assign N252 = N250;
  assign N253 = valid_o[4] & 1'b1;
  assign N254 = ~N253;
  assign N255 = N252 & N253;
  assign N264 = new_valid_0__0_ & arb_grants_r_0__0_;
  assign N265 = new_valid_0__1_ & arb_grants_r_0__1_;
  assign N266 = new_valid_0__2_ & arb_grants_r_0__2_;
  assign N267 = new_valid_0__3_ & arb_grants_r_0__3_;
  assign N268 = new_valid_0__4_ & arb_grants_r_0__4_;
  assign N269 = new_valid_1__0_ & arb_grants_r_1__0_;
  assign N270 = new_valid_1__2_ & arb_grants_r_1__2_;
  assign N271 = new_valid_1__3_ & arb_grants_r_1__3_;
  assign N272 = new_valid_1__4_ & arb_grants_r_1__4_;
  assign N273 = new_valid_2__0_ & arb_grants_r_2__0_;
  assign N274 = new_valid_2__1_ & arb_grants_r_2__1_;
  assign N275 = new_valid_2__3_ & arb_grants_r_2__3_;
  assign N276 = new_valid_2__4_ & arb_grants_r_2__4_;
  assign N277 = new_valid_3__0_ & arb_grants_r_3__0_;
  assign N278 = new_valid_3__1_ & arb_grants_r_3__1_;
  assign N279 = new_valid_3__2_ & arb_grants_r_3__2_;
  assign N280 = new_valid_3__4_ & arb_grants_r_3__4_;
  assign N281 = new_valid_4__0_ & arb_grants_r_4__0_;
  assign N282 = new_valid_4__1_ & arb_grants_r_4__1_;
  assign N283 = new_valid_4__2_ & arb_grants_r_4__2_;
  assign N284 = new_valid_4__3_ & arb_grants_r_4__3_;
  assign n_3_net_ = valid_o[1] & 1'b1;
  assign n_9_net_ = valid_o[2] & ready_i[2];
  assign n_15_net_ = valid_o[3] & 1'b1;
  assign n_21_net_ = valid_o[4] & 1'b1;
  assign n_27_net_ = valid_o[0] & ready_i[0];
  assign N293 = ~N292;
  assign N301 = ~N300;
  assign N310 = ~N309;
  assign N318 = ~N381;
  assign N319 = ~N382;
  assign N320 = ~N383;
  assign N321 = ~N384;
  assign N322 = ~N385;
  assign N323 = ~N386;
  assign N324 = ~N387;
  assign N325 = ~N388;
  assign N326 = ~N389;
  assign N327 = ~N390;
  assign N328 = ~N391;
  assign N329 = ~N392;
  assign N330 = ~N393;
  assign N331 = ~N394;
  assign N332 = ~N395;
  assign N333 = ~N396;
  assign N334 = ~N397;
  assign N335 = ~N398;
  assign N336 = ~N399;
  assign N337 = ~N400;
  assign N338 = ~N401;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { count_r[9:0] } <= { N193, N192, N179, N178, N165, N164, N151, N150, N138, N137 };
      dest_r_0__4_ <= dest_n_0__4_;
      dest_r_0__3_ <= dest_n_0__3_;
      dest_r_0__2_ <= dest_n_0__2_;
      dest_r_0__1_ <= dest_n_0__1_;
      dest_r_0__0_ <= dest_n_0__0_;
      dest_r_1__4_ <= dest_n_1__4_;
      dest_r_1__3_ <= dest_n_1__3_;
      dest_r_1__2_ <= dest_n_1__2_;
      dest_r_1__0_ <= dest_n_1__0_;
      dest_r_2__4_ <= dest_n_2__4_;
      dest_r_2__3_ <= dest_n_2__3_;
      dest_r_2__1_ <= dest_n_2__1_;
      dest_r_2__0_ <= dest_n_2__0_;
      dest_r_3__4_ <= dest_n_3__4_;
      dest_r_3__2_ <= dest_n_3__2_;
      dest_r_3__1_ <= dest_n_3__1_;
      dest_r_3__0_ <= dest_n_3__0_;
      dest_r_4__3_ <= dest_n_4__3_;
      dest_r_4__2_ <= dest_n_4__2_;
      dest_r_4__1_ <= dest_n_4__1_;
      dest_r_4__0_ <= dest_n_4__0_;
      { out_count_r[9:0] } <= { N263, N262, N249, N248, N235, N234, N221, N220, N207, N206 };
    end
    if(N318) begin
      arb_grants_r_0__0_ <= arb_grants_o_0__0_;
    end
    if(N319) begin
      arb_grants_r_0__1_ <= arb_grants_o_0__1_;
    end
    if(N320) begin
      arb_grants_r_0__2_ <= arb_grants_o_0__2_;
    end
    if(N321) begin
      arb_grants_r_0__3_ <= arb_grants_o_0__3_;
    end
    if(N322) begin
      arb_grants_r_0__4_ <= arb_grants_o_0__4_;
    end
    if(N323) begin
      arb_grants_r_1__0_ <= arb_grants_o_1__0_;
    end
    if(N324) begin
      arb_grants_r_1__2_ <= arb_grants_o_1__2_;
    end
    if(N325) begin
      arb_grants_r_1__3_ <= arb_grants_o_1__3_;
    end
    if(N326) begin
      arb_grants_r_1__4_ <= arb_grants_o_1__4_;
    end
    if(N327) begin
      arb_grants_r_2__0_ <= arb_grants_o_2__0_;
    end
    if(N328) begin
      arb_grants_r_2__1_ <= arb_grants_o_2__1_;
    end
    if(N329) begin
      arb_grants_r_2__3_ <= arb_grants_o_2__3_;
    end
    if(N330) begin
      arb_grants_r_2__4_ <= arb_grants_o_2__4_;
    end
    if(N331) begin
      arb_grants_r_3__0_ <= arb_grants_o_3__0_;
    end
    if(N332) begin
      arb_grants_r_3__1_ <= arb_grants_o_3__1_;
    end
    if(N333) begin
      arb_grants_r_3__2_ <= arb_grants_o_3__2_;
    end
    if(N334) begin
      arb_grants_r_3__4_ <= arb_grants_o_3__4_;
    end
    if(N335) begin
      arb_grants_r_4__0_ <= arb_grants_o_4__0_;
    end
    if(N336) begin
      arb_grants_r_4__1_ <= arb_grants_o_4__1_;
    end
    if(N337) begin
      arb_grants_r_4__2_ <= arb_grants_o_4__2_;
    end
    if(N338) begin
      arb_grants_r_4__3_ <= arb_grants_o_4__3_;
    end
  end


endmodule



module bsg_wormhole_router_131_1_1_2_1_1_1_00000015_0000001c
(
  clk_i,
  reset_i,
  local_x_cord_i,
  local_y_cord_i,
  valid_i,
  data_i,
  ready_o,
  valid_o,
  data_o,
  ready_i
);

  input [0:0] local_x_cord_i;
  input [0:0] local_y_cord_i;
  input [4:0] valid_i;
  input [654:0] data_i;
  output [4:0] ready_o;
  output [4:0] valid_o;
  output [654:0] data_o;
  input [4:0] ready_i;
  input clk_i;
  input reset_i;
  wire [4:0] ready_o,valid_o,fifo_yumi_i;
  wire [654:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,fifo_valid_o_1,fifo_data_o_3__130_,fifo_data_o_3__129_,
  fifo_data_o_3__128_,fifo_data_o_3__127_,fifo_data_o_3__126_,fifo_data_o_3__125_,
  fifo_data_o_3__124_,fifo_data_o_3__123_,fifo_data_o_3__122_,fifo_data_o_3__121_,
  fifo_data_o_3__120_,fifo_data_o_3__119_,fifo_data_o_3__118_,fifo_data_o_3__117_,
  fifo_data_o_3__116_,fifo_data_o_3__115_,fifo_data_o_3__114_,fifo_data_o_3__113_,
  fifo_data_o_3__112_,fifo_data_o_3__111_,fifo_data_o_3__110_,fifo_data_o_3__109_,
  fifo_data_o_3__108_,fifo_data_o_3__107_,fifo_data_o_3__106_,fifo_data_o_3__105_,
  fifo_data_o_3__104_,fifo_data_o_3__103_,fifo_data_o_3__102_,fifo_data_o_3__101_,
  fifo_data_o_3__100_,fifo_data_o_3__99_,fifo_data_o_3__98_,fifo_data_o_3__97_,
  fifo_data_o_3__96_,fifo_data_o_3__95_,fifo_data_o_3__94_,fifo_data_o_3__93_,fifo_data_o_3__92_,
  fifo_data_o_3__91_,fifo_data_o_3__90_,fifo_data_o_3__89_,fifo_data_o_3__88_,
  fifo_data_o_3__87_,fifo_data_o_3__86_,fifo_data_o_3__85_,fifo_data_o_3__84_,
  fifo_data_o_3__83_,fifo_data_o_3__82_,fifo_data_o_3__81_,fifo_data_o_3__80_,
  fifo_data_o_3__79_,fifo_data_o_3__78_,fifo_data_o_3__77_,fifo_data_o_3__76_,fifo_data_o_3__75_,
  fifo_data_o_3__74_,fifo_data_o_3__73_,fifo_data_o_3__72_,fifo_data_o_3__71_,
  fifo_data_o_3__70_,fifo_data_o_3__69_,fifo_data_o_3__68_,fifo_data_o_3__67_,
  fifo_data_o_3__66_,fifo_data_o_3__65_,fifo_data_o_3__64_,fifo_data_o_3__63_,
  fifo_data_o_3__62_,fifo_data_o_3__61_,fifo_data_o_3__60_,fifo_data_o_3__59_,
  fifo_data_o_3__58_,fifo_data_o_3__57_,fifo_data_o_3__56_,fifo_data_o_3__55_,fifo_data_o_3__54_,
  fifo_data_o_3__53_,fifo_data_o_3__52_,fifo_data_o_3__51_,fifo_data_o_3__50_,
  fifo_data_o_3__49_,fifo_data_o_3__48_,fifo_data_o_3__47_,fifo_data_o_3__46_,
  fifo_data_o_3__45_,fifo_data_o_3__44_,fifo_data_o_3__43_,fifo_data_o_3__42_,
  fifo_data_o_3__41_,fifo_data_o_3__40_,fifo_data_o_3__39_,fifo_data_o_3__38_,
  fifo_data_o_3__37_,fifo_data_o_3__36_,fifo_data_o_3__35_,fifo_data_o_3__34_,fifo_data_o_3__33_,
  fifo_data_o_3__32_,fifo_data_o_3__31_,fifo_data_o_3__30_,fifo_data_o_3__29_,
  fifo_data_o_3__28_,fifo_data_o_3__27_,fifo_data_o_3__26_,fifo_data_o_3__25_,
  fifo_data_o_3__24_,fifo_data_o_3__23_,fifo_data_o_3__22_,fifo_data_o_3__21_,
  fifo_data_o_3__20_,fifo_data_o_3__19_,fifo_data_o_3__18_,fifo_data_o_3__17_,
  fifo_data_o_3__16_,fifo_data_o_3__15_,fifo_data_o_3__14_,fifo_data_o_3__13_,fifo_data_o_3__12_,
  fifo_data_o_3__11_,fifo_data_o_3__10_,fifo_data_o_3__9_,fifo_data_o_3__8_,
  fifo_data_o_3__7_,fifo_data_o_3__6_,fifo_data_o_3__5_,fifo_data_o_3__4_,
  fifo_data_o_3__3_,fifo_data_o_3__2_,fifo_data_o_3__1_,fifo_data_o_3__0_,fifo_data_o_1__130_,
  fifo_data_o_1__129_,fifo_data_o_1__128_,fifo_data_o_1__127_,fifo_data_o_1__126_,
  fifo_data_o_1__125_,fifo_data_o_1__124_,fifo_data_o_1__123_,fifo_data_o_1__122_,
  fifo_data_o_1__121_,fifo_data_o_1__120_,fifo_data_o_1__119_,fifo_data_o_1__118_,
  fifo_data_o_1__117_,fifo_data_o_1__116_,fifo_data_o_1__115_,fifo_data_o_1__114_,
  fifo_data_o_1__113_,fifo_data_o_1__112_,fifo_data_o_1__111_,fifo_data_o_1__110_,
  fifo_data_o_1__109_,fifo_data_o_1__108_,fifo_data_o_1__107_,fifo_data_o_1__106_,
  fifo_data_o_1__105_,fifo_data_o_1__104_,fifo_data_o_1__103_,fifo_data_o_1__102_,
  fifo_data_o_1__101_,fifo_data_o_1__100_,fifo_data_o_1__99_,fifo_data_o_1__98_,
  fifo_data_o_1__97_,fifo_data_o_1__96_,fifo_data_o_1__95_,fifo_data_o_1__94_,
  fifo_data_o_1__93_,fifo_data_o_1__92_,fifo_data_o_1__91_,fifo_data_o_1__90_,
  fifo_data_o_1__89_,fifo_data_o_1__88_,fifo_data_o_1__87_,fifo_data_o_1__86_,fifo_data_o_1__85_,
  fifo_data_o_1__84_,fifo_data_o_1__83_,fifo_data_o_1__82_,fifo_data_o_1__81_,
  fifo_data_o_1__80_,fifo_data_o_1__79_,fifo_data_o_1__78_,fifo_data_o_1__77_,
  fifo_data_o_1__76_,fifo_data_o_1__75_,fifo_data_o_1__74_,fifo_data_o_1__73_,
  fifo_data_o_1__72_,fifo_data_o_1__71_,fifo_data_o_1__70_,fifo_data_o_1__69_,
  fifo_data_o_1__68_,fifo_data_o_1__67_,fifo_data_o_1__66_,fifo_data_o_1__65_,fifo_data_o_1__64_,
  fifo_data_o_1__63_,fifo_data_o_1__62_,fifo_data_o_1__61_,fifo_data_o_1__60_,
  fifo_data_o_1__59_,fifo_data_o_1__58_,fifo_data_o_1__57_,fifo_data_o_1__56_,
  fifo_data_o_1__55_,fifo_data_o_1__54_,fifo_data_o_1__53_,fifo_data_o_1__52_,
  fifo_data_o_1__51_,fifo_data_o_1__50_,fifo_data_o_1__49_,fifo_data_o_1__48_,
  fifo_data_o_1__47_,fifo_data_o_1__46_,fifo_data_o_1__45_,fifo_data_o_1__44_,fifo_data_o_1__43_,
  fifo_data_o_1__42_,fifo_data_o_1__41_,fifo_data_o_1__40_,fifo_data_o_1__39_,
  fifo_data_o_1__38_,fifo_data_o_1__37_,fifo_data_o_1__36_,fifo_data_o_1__35_,
  fifo_data_o_1__34_,fifo_data_o_1__33_,fifo_data_o_1__32_,fifo_data_o_1__31_,
  fifo_data_o_1__30_,fifo_data_o_1__29_,fifo_data_o_1__28_,fifo_data_o_1__27_,
  fifo_data_o_1__26_,fifo_data_o_1__25_,fifo_data_o_1__24_,fifo_data_o_1__23_,fifo_data_o_1__22_,
  fifo_data_o_1__21_,fifo_data_o_1__20_,fifo_data_o_1__19_,fifo_data_o_1__18_,
  fifo_data_o_1__17_,fifo_data_o_1__16_,fifo_data_o_1__15_,fifo_data_o_1__14_,
  fifo_data_o_1__13_,fifo_data_o_1__12_,fifo_data_o_1__11_,fifo_data_o_1__10_,
  fifo_data_o_1__9_,fifo_data_o_1__8_,fifo_data_o_1__7_,fifo_data_o_1__6_,fifo_data_o_1__5_,
  fifo_data_o_1__4_,fifo_data_o_1__3_,fifo_data_o_1__2_,fifo_data_o_1__1_,
  fifo_data_o_1__0_,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,
  N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,
  N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,
  N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,
  N183,N184,N185,N186,dest_n_4__3_,dest_n_4__2_,dest_n_4__1_,dest_n_4__0_,
  dest_n_3__4_,dest_n_3__2_,dest_n_3__1_,dest_n_3__0_,dest_n_2__4_,dest_n_2__3_,
  dest_n_2__1_,dest_n_2__0_,dest_n_1__4_,dest_n_1__3_,dest_n_1__2_,dest_n_1__0_,
  dest_n_0__4_,dest_n_0__3_,dest_n_0__2_,dest_n_0__1_,dest_n_0__0_,new_valid_4__3_,
  new_valid_4__2_,new_valid_4__1_,new_valid_4__0_,new_valid_3__4_,new_valid_3__2_,
  new_valid_3__1_,new_valid_3__0_,new_valid_2__4_,new_valid_2__3_,new_valid_2__1_,
  new_valid_2__0_,new_valid_1__4_,new_valid_1__3_,new_valid_1__2_,new_valid_1__0_,
  new_valid_0__4_,new_valid_0__3_,new_valid_0__2_,new_valid_0__1_,new_valid_0__0_,
  arb_grants_o_4__3_,arb_grants_o_4__2_,arb_grants_o_4__1_,arb_grants_o_4__0_,
  arb_grants_o_3__4_,arb_grants_o_3__2_,arb_grants_o_3__1_,arb_grants_o_3__0_,arb_grants_o_2__4_,
  arb_grants_o_2__3_,arb_grants_o_2__1_,arb_grants_o_2__0_,arb_grants_o_1__4_,
  arb_grants_o_1__3_,arb_grants_o_1__2_,arb_grants_o_1__0_,arb_grants_o_0__4_,
  arb_grants_o_0__3_,arb_grants_o_0__2_,arb_grants_o_0__1_,arb_grants_o_0__0_,N187,N188,
  N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,
  N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,
  N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,
  N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,
  N253,N254,N255,N256,N257,arb_valid_4__3_,arb_valid_4__2_,arb_valid_4__1_,
  arb_valid_4__0_,arb_valid_3__4_,arb_valid_3__2_,arb_valid_3__1_,arb_valid_3__0_,
  arb_valid_2__4_,arb_valid_2__3_,arb_valid_2__1_,arb_valid_2__0_,arb_valid_1__4_,
  arb_valid_1__3_,arb_valid_1__2_,arb_valid_1__0_,arb_valid_0__4_,arb_valid_0__3_,
  arb_valid_0__2_,arb_valid_0__1_,arb_valid_0__0_,N258,N259,N260,N261,N262,N263,N264,N265,
  N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,n_3_net_,
  arb_sel_o_4__3_,arb_sel_o_4__2_,arb_sel_o_4__1_,arb_sel_o_4__0_,arb_sel_o_3__3_,
  arb_sel_o_3__2_,arb_sel_o_3__1_,arb_sel_o_3__0_,arb_sel_o_2__3_,arb_sel_o_2__2_,
  arb_sel_o_2__1_,arb_sel_o_2__0_,arb_sel_o_1__3_,arb_sel_o_1__2_,arb_sel_o_1__1_,
  arb_sel_o_1__0_,arb_sel_o_0__4_,arb_sel_o_0__3_,arb_sel_o_0__2_,arb_sel_o_0__1_,
  arb_sel_o_0__0_,n_9_net_,n_15_net_,n_21_net_,n_27_net_,N278,N279,N280,N281,N282,N283,N284,
  N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,
  N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,
  N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,
  N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
  N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,
  N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,
  N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,
  N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,
  N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,
  N429,N430,N431,N432,SV2V_UNCONNECTED_1,SV2V_UNCONNECTED_2,
  SV2V_UNCONNECTED_3,SV2V_UNCONNECTED_4,SV2V_UNCONNECTED_5,SV2V_UNCONNECTED_6,
  SV2V_UNCONNECTED_7,SV2V_UNCONNECTED_8,SV2V_UNCONNECTED_9,
  SV2V_UNCONNECTED_10,SV2V_UNCONNECTED_11;
  wire [3:3] fifo_valid_o;
  reg [9:0] count_r,out_count_r;
  reg dest_r_0__4_,dest_r_0__3_,dest_r_0__2_,dest_r_0__1_,dest_r_0__0_,dest_r_1__4_,
  dest_r_1__3_,dest_r_1__2_,dest_r_1__0_,dest_r_2__4_,dest_r_2__3_,dest_r_2__1_,
  dest_r_2__0_,dest_r_3__4_,dest_r_3__2_,dest_r_3__1_,dest_r_3__0_,dest_r_4__3_,
  dest_r_4__2_,dest_r_4__1_,dest_r_4__0_,arb_grants_r_0__0_,arb_grants_r_0__1_,
  arb_grants_r_0__2_,arb_grants_r_0__3_,arb_grants_r_0__4_,arb_grants_r_1__0_,
  arb_grants_r_1__2_,arb_grants_r_1__3_,arb_grants_r_1__4_,arb_grants_r_2__0_,
  arb_grants_r_2__1_,arb_grants_r_2__3_,arb_grants_r_2__4_,arb_grants_r_3__0_,arb_grants_r_3__1_,
  arb_grants_r_3__2_,arb_grants_r_3__4_,arb_grants_r_4__0_,arb_grants_r_4__1_,
  arb_grants_r_4__2_,arb_grants_r_4__3_;
  assign ready_o[4] = 1'b1;
  assign ready_o[2] = 1'b1;
  assign ready_o[0] = 1'b1;

  bsg_two_fifo_width_p131
  in_ff_1__no_stub_two_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(ready_o[1]),
    .data_i(data_i[261:131]),
    .v_i(valid_i[1]),
    .v_o(fifo_valid_o_1),
    .data_o({ fifo_data_o_1__130_, fifo_data_o_1__129_, fifo_data_o_1__128_, fifo_data_o_1__127_, fifo_data_o_1__126_, fifo_data_o_1__125_, fifo_data_o_1__124_, fifo_data_o_1__123_, fifo_data_o_1__122_, fifo_data_o_1__121_, fifo_data_o_1__120_, fifo_data_o_1__119_, fifo_data_o_1__118_, fifo_data_o_1__117_, fifo_data_o_1__116_, fifo_data_o_1__115_, fifo_data_o_1__114_, fifo_data_o_1__113_, fifo_data_o_1__112_, fifo_data_o_1__111_, fifo_data_o_1__110_, fifo_data_o_1__109_, fifo_data_o_1__108_, fifo_data_o_1__107_, fifo_data_o_1__106_, fifo_data_o_1__105_, fifo_data_o_1__104_, fifo_data_o_1__103_, fifo_data_o_1__102_, fifo_data_o_1__101_, fifo_data_o_1__100_, fifo_data_o_1__99_, fifo_data_o_1__98_, fifo_data_o_1__97_, fifo_data_o_1__96_, fifo_data_o_1__95_, fifo_data_o_1__94_, fifo_data_o_1__93_, fifo_data_o_1__92_, fifo_data_o_1__91_, fifo_data_o_1__90_, fifo_data_o_1__89_, fifo_data_o_1__88_, fifo_data_o_1__87_, fifo_data_o_1__86_, fifo_data_o_1__85_, fifo_data_o_1__84_, fifo_data_o_1__83_, fifo_data_o_1__82_, fifo_data_o_1__81_, fifo_data_o_1__80_, fifo_data_o_1__79_, fifo_data_o_1__78_, fifo_data_o_1__77_, fifo_data_o_1__76_, fifo_data_o_1__75_, fifo_data_o_1__74_, fifo_data_o_1__73_, fifo_data_o_1__72_, fifo_data_o_1__71_, fifo_data_o_1__70_, fifo_data_o_1__69_, fifo_data_o_1__68_, fifo_data_o_1__67_, fifo_data_o_1__66_, fifo_data_o_1__65_, fifo_data_o_1__64_, fifo_data_o_1__63_, fifo_data_o_1__62_, fifo_data_o_1__61_, fifo_data_o_1__60_, fifo_data_o_1__59_, fifo_data_o_1__58_, fifo_data_o_1__57_, fifo_data_o_1__56_, fifo_data_o_1__55_, fifo_data_o_1__54_, fifo_data_o_1__53_, fifo_data_o_1__52_, fifo_data_o_1__51_, fifo_data_o_1__50_, fifo_data_o_1__49_, fifo_data_o_1__48_, fifo_data_o_1__47_, fifo_data_o_1__46_, fifo_data_o_1__45_, fifo_data_o_1__44_, fifo_data_o_1__43_, fifo_data_o_1__42_, fifo_data_o_1__41_, fifo_data_o_1__40_, fifo_data_o_1__39_, fifo_data_o_1__38_, fifo_data_o_1__37_, fifo_data_o_1__36_, fifo_data_o_1__35_, fifo_data_o_1__34_, fifo_data_o_1__33_, fifo_data_o_1__32_, fifo_data_o_1__31_, fifo_data_o_1__30_, fifo_data_o_1__29_, fifo_data_o_1__28_, fifo_data_o_1__27_, fifo_data_o_1__26_, fifo_data_o_1__25_, fifo_data_o_1__24_, fifo_data_o_1__23_, fifo_data_o_1__22_, fifo_data_o_1__21_, fifo_data_o_1__20_, fifo_data_o_1__19_, fifo_data_o_1__18_, fifo_data_o_1__17_, fifo_data_o_1__16_, fifo_data_o_1__15_, fifo_data_o_1__14_, fifo_data_o_1__13_, fifo_data_o_1__12_, fifo_data_o_1__11_, fifo_data_o_1__10_, fifo_data_o_1__9_, fifo_data_o_1__8_, fifo_data_o_1__7_, fifo_data_o_1__6_, fifo_data_o_1__5_, fifo_data_o_1__4_, fifo_data_o_1__3_, fifo_data_o_1__2_, fifo_data_o_1__1_, fifo_data_o_1__0_ }),
    .yumi_i(fifo_yumi_i[1])
  );


  bsg_two_fifo_width_p131
  in_ff_3__no_stub_two_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(ready_o[3]),
    .data_i(data_i[523:393]),
    .v_i(valid_i[3]),
    .v_o(fifo_valid_o[3]),
    .data_o({ fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_ }),
    .yumi_i(fifo_yumi_i[3])
  );


  bsg_round_robin_arb_inputs_p4
  out_side_1__rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[1]),
    .reqs_i({ arb_valid_4__1_, arb_valid_3__1_, arb_valid_2__1_, arb_valid_0__1_ }),
    .grants_o({ arb_grants_o_4__1_, arb_grants_o_3__1_, arb_grants_o_2__1_, arb_grants_o_0__1_ }),
    .sel_one_hot_o({ arb_sel_o_1__3_, arb_sel_o_1__2_, arb_sel_o_1__1_, arb_sel_o_1__0_ }),
    .v_o(valid_o[1]),
    .tag_o({ SV2V_UNCONNECTED_1, SV2V_UNCONNECTED_2 }),
    .yumi_i(n_3_net_)
  );


  bsg_mux_one_hot_width_p131_els_p4
  out_side_1__mux
  (
    .data_i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_1__3_, arb_sel_o_1__2_, arb_sel_o_1__1_, arb_sel_o_1__0_ }),
    .data_o(data_o[261:131])
  );


  bsg_round_robin_arb_inputs_p4
  out_side_2__rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ arb_valid_4__2_, arb_valid_3__2_, arb_valid_1__2_, arb_valid_0__2_ }),
    .grants_o({ arb_grants_o_4__2_, arb_grants_o_3__2_, arb_grants_o_1__2_, arb_grants_o_0__2_ }),
    .sel_one_hot_o({ arb_sel_o_2__3_, arb_sel_o_2__2_, arb_sel_o_2__1_, arb_sel_o_2__0_ }),
    .v_o(valid_o[2]),
    .tag_o({ SV2V_UNCONNECTED_3, SV2V_UNCONNECTED_4 }),
    .yumi_i(n_9_net_)
  );


  bsg_mux_one_hot_width_p131_els_p4
  out_side_2__mux
  (
    .data_i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_, fifo_data_o_1__130_, fifo_data_o_1__129_, fifo_data_o_1__128_, fifo_data_o_1__127_, fifo_data_o_1__126_, fifo_data_o_1__125_, fifo_data_o_1__124_, fifo_data_o_1__123_, fifo_data_o_1__122_, fifo_data_o_1__121_, fifo_data_o_1__120_, fifo_data_o_1__119_, fifo_data_o_1__118_, fifo_data_o_1__117_, fifo_data_o_1__116_, fifo_data_o_1__115_, fifo_data_o_1__114_, fifo_data_o_1__113_, fifo_data_o_1__112_, fifo_data_o_1__111_, fifo_data_o_1__110_, fifo_data_o_1__109_, fifo_data_o_1__108_, fifo_data_o_1__107_, fifo_data_o_1__106_, fifo_data_o_1__105_, fifo_data_o_1__104_, fifo_data_o_1__103_, fifo_data_o_1__102_, fifo_data_o_1__101_, fifo_data_o_1__100_, fifo_data_o_1__99_, fifo_data_o_1__98_, fifo_data_o_1__97_, fifo_data_o_1__96_, fifo_data_o_1__95_, fifo_data_o_1__94_, fifo_data_o_1__93_, fifo_data_o_1__92_, fifo_data_o_1__91_, fifo_data_o_1__90_, fifo_data_o_1__89_, fifo_data_o_1__88_, fifo_data_o_1__87_, fifo_data_o_1__86_, fifo_data_o_1__85_, fifo_data_o_1__84_, fifo_data_o_1__83_, fifo_data_o_1__82_, fifo_data_o_1__81_, fifo_data_o_1__80_, fifo_data_o_1__79_, fifo_data_o_1__78_, fifo_data_o_1__77_, fifo_data_o_1__76_, fifo_data_o_1__75_, fifo_data_o_1__74_, fifo_data_o_1__73_, fifo_data_o_1__72_, fifo_data_o_1__71_, fifo_data_o_1__70_, fifo_data_o_1__69_, fifo_data_o_1__68_, fifo_data_o_1__67_, fifo_data_o_1__66_, fifo_data_o_1__65_, fifo_data_o_1__64_, fifo_data_o_1__63_, fifo_data_o_1__62_, fifo_data_o_1__61_, fifo_data_o_1__60_, fifo_data_o_1__59_, fifo_data_o_1__58_, fifo_data_o_1__57_, fifo_data_o_1__56_, fifo_data_o_1__55_, fifo_data_o_1__54_, fifo_data_o_1__53_, fifo_data_o_1__52_, fifo_data_o_1__51_, fifo_data_o_1__50_, fifo_data_o_1__49_, fifo_data_o_1__48_, fifo_data_o_1__47_, fifo_data_o_1__46_, fifo_data_o_1__45_, fifo_data_o_1__44_, fifo_data_o_1__43_, fifo_data_o_1__42_, fifo_data_o_1__41_, fifo_data_o_1__40_, fifo_data_o_1__39_, fifo_data_o_1__38_, fifo_data_o_1__37_, fifo_data_o_1__36_, fifo_data_o_1__35_, fifo_data_o_1__34_, fifo_data_o_1__33_, fifo_data_o_1__32_, fifo_data_o_1__31_, fifo_data_o_1__30_, fifo_data_o_1__29_, fifo_data_o_1__28_, fifo_data_o_1__27_, fifo_data_o_1__26_, fifo_data_o_1__25_, fifo_data_o_1__24_, fifo_data_o_1__23_, fifo_data_o_1__22_, fifo_data_o_1__21_, fifo_data_o_1__20_, fifo_data_o_1__19_, fifo_data_o_1__18_, fifo_data_o_1__17_, fifo_data_o_1__16_, fifo_data_o_1__15_, fifo_data_o_1__14_, fifo_data_o_1__13_, fifo_data_o_1__12_, fifo_data_o_1__11_, fifo_data_o_1__10_, fifo_data_o_1__9_, fifo_data_o_1__8_, fifo_data_o_1__7_, fifo_data_o_1__6_, fifo_data_o_1__5_, fifo_data_o_1__4_, fifo_data_o_1__3_, fifo_data_o_1__2_, fifo_data_o_1__1_, fifo_data_o_1__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_2__3_, arb_sel_o_2__2_, arb_sel_o_2__1_, arb_sel_o_2__0_ }),
    .data_o(data_o[392:262])
  );


  bsg_round_robin_arb_inputs_p4
  out_side_3__rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ arb_valid_4__3_, arb_valid_2__3_, arb_valid_1__3_, arb_valid_0__3_ }),
    .grants_o({ arb_grants_o_4__3_, arb_grants_o_2__3_, arb_grants_o_1__3_, arb_grants_o_0__3_ }),
    .sel_one_hot_o({ arb_sel_o_3__3_, arb_sel_o_3__2_, arb_sel_o_3__1_, arb_sel_o_3__0_ }),
    .v_o(valid_o[3]),
    .tag_o({ SV2V_UNCONNECTED_5, SV2V_UNCONNECTED_6 }),
    .yumi_i(n_15_net_)
  );


  bsg_mux_one_hot_width_p131_els_p4
  out_side_3__mux
  (
    .data_i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_o_1__130_, fifo_data_o_1__129_, fifo_data_o_1__128_, fifo_data_o_1__127_, fifo_data_o_1__126_, fifo_data_o_1__125_, fifo_data_o_1__124_, fifo_data_o_1__123_, fifo_data_o_1__122_, fifo_data_o_1__121_, fifo_data_o_1__120_, fifo_data_o_1__119_, fifo_data_o_1__118_, fifo_data_o_1__117_, fifo_data_o_1__116_, fifo_data_o_1__115_, fifo_data_o_1__114_, fifo_data_o_1__113_, fifo_data_o_1__112_, fifo_data_o_1__111_, fifo_data_o_1__110_, fifo_data_o_1__109_, fifo_data_o_1__108_, fifo_data_o_1__107_, fifo_data_o_1__106_, fifo_data_o_1__105_, fifo_data_o_1__104_, fifo_data_o_1__103_, fifo_data_o_1__102_, fifo_data_o_1__101_, fifo_data_o_1__100_, fifo_data_o_1__99_, fifo_data_o_1__98_, fifo_data_o_1__97_, fifo_data_o_1__96_, fifo_data_o_1__95_, fifo_data_o_1__94_, fifo_data_o_1__93_, fifo_data_o_1__92_, fifo_data_o_1__91_, fifo_data_o_1__90_, fifo_data_o_1__89_, fifo_data_o_1__88_, fifo_data_o_1__87_, fifo_data_o_1__86_, fifo_data_o_1__85_, fifo_data_o_1__84_, fifo_data_o_1__83_, fifo_data_o_1__82_, fifo_data_o_1__81_, fifo_data_o_1__80_, fifo_data_o_1__79_, fifo_data_o_1__78_, fifo_data_o_1__77_, fifo_data_o_1__76_, fifo_data_o_1__75_, fifo_data_o_1__74_, fifo_data_o_1__73_, fifo_data_o_1__72_, fifo_data_o_1__71_, fifo_data_o_1__70_, fifo_data_o_1__69_, fifo_data_o_1__68_, fifo_data_o_1__67_, fifo_data_o_1__66_, fifo_data_o_1__65_, fifo_data_o_1__64_, fifo_data_o_1__63_, fifo_data_o_1__62_, fifo_data_o_1__61_, fifo_data_o_1__60_, fifo_data_o_1__59_, fifo_data_o_1__58_, fifo_data_o_1__57_, fifo_data_o_1__56_, fifo_data_o_1__55_, fifo_data_o_1__54_, fifo_data_o_1__53_, fifo_data_o_1__52_, fifo_data_o_1__51_, fifo_data_o_1__50_, fifo_data_o_1__49_, fifo_data_o_1__48_, fifo_data_o_1__47_, fifo_data_o_1__46_, fifo_data_o_1__45_, fifo_data_o_1__44_, fifo_data_o_1__43_, fifo_data_o_1__42_, fifo_data_o_1__41_, fifo_data_o_1__40_, fifo_data_o_1__39_, fifo_data_o_1__38_, fifo_data_o_1__37_, fifo_data_o_1__36_, fifo_data_o_1__35_, fifo_data_o_1__34_, fifo_data_o_1__33_, fifo_data_o_1__32_, fifo_data_o_1__31_, fifo_data_o_1__30_, fifo_data_o_1__29_, fifo_data_o_1__28_, fifo_data_o_1__27_, fifo_data_o_1__26_, fifo_data_o_1__25_, fifo_data_o_1__24_, fifo_data_o_1__23_, fifo_data_o_1__22_, fifo_data_o_1__21_, fifo_data_o_1__20_, fifo_data_o_1__19_, fifo_data_o_1__18_, fifo_data_o_1__17_, fifo_data_o_1__16_, fifo_data_o_1__15_, fifo_data_o_1__14_, fifo_data_o_1__13_, fifo_data_o_1__12_, fifo_data_o_1__11_, fifo_data_o_1__10_, fifo_data_o_1__9_, fifo_data_o_1__8_, fifo_data_o_1__7_, fifo_data_o_1__6_, fifo_data_o_1__5_, fifo_data_o_1__4_, fifo_data_o_1__3_, fifo_data_o_1__2_, fifo_data_o_1__1_, fifo_data_o_1__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_3__3_, arb_sel_o_3__2_, arb_sel_o_3__1_, arb_sel_o_3__0_ }),
    .data_o(data_o[523:393])
  );


  bsg_round_robin_arb_inputs_p4
  out_side_4__rr_arb
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(1'b1),
    .reqs_i({ arb_valid_3__4_, arb_valid_2__4_, arb_valid_1__4_, arb_valid_0__4_ }),
    .grants_o({ arb_grants_o_3__4_, arb_grants_o_2__4_, arb_grants_o_1__4_, arb_grants_o_0__4_ }),
    .sel_one_hot_o({ arb_sel_o_4__3_, arb_sel_o_4__2_, arb_sel_o_4__1_, arb_sel_o_4__0_ }),
    .v_o(valid_o[4]),
    .tag_o({ SV2V_UNCONNECTED_7, SV2V_UNCONNECTED_8 }),
    .yumi_i(n_21_net_)
  );


  bsg_mux_one_hot_width_p131_els_p4
  out_side_4__mux
  (
    .data_i({ fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_o_1__130_, fifo_data_o_1__129_, fifo_data_o_1__128_, fifo_data_o_1__127_, fifo_data_o_1__126_, fifo_data_o_1__125_, fifo_data_o_1__124_, fifo_data_o_1__123_, fifo_data_o_1__122_, fifo_data_o_1__121_, fifo_data_o_1__120_, fifo_data_o_1__119_, fifo_data_o_1__118_, fifo_data_o_1__117_, fifo_data_o_1__116_, fifo_data_o_1__115_, fifo_data_o_1__114_, fifo_data_o_1__113_, fifo_data_o_1__112_, fifo_data_o_1__111_, fifo_data_o_1__110_, fifo_data_o_1__109_, fifo_data_o_1__108_, fifo_data_o_1__107_, fifo_data_o_1__106_, fifo_data_o_1__105_, fifo_data_o_1__104_, fifo_data_o_1__103_, fifo_data_o_1__102_, fifo_data_o_1__101_, fifo_data_o_1__100_, fifo_data_o_1__99_, fifo_data_o_1__98_, fifo_data_o_1__97_, fifo_data_o_1__96_, fifo_data_o_1__95_, fifo_data_o_1__94_, fifo_data_o_1__93_, fifo_data_o_1__92_, fifo_data_o_1__91_, fifo_data_o_1__90_, fifo_data_o_1__89_, fifo_data_o_1__88_, fifo_data_o_1__87_, fifo_data_o_1__86_, fifo_data_o_1__85_, fifo_data_o_1__84_, fifo_data_o_1__83_, fifo_data_o_1__82_, fifo_data_o_1__81_, fifo_data_o_1__80_, fifo_data_o_1__79_, fifo_data_o_1__78_, fifo_data_o_1__77_, fifo_data_o_1__76_, fifo_data_o_1__75_, fifo_data_o_1__74_, fifo_data_o_1__73_, fifo_data_o_1__72_, fifo_data_o_1__71_, fifo_data_o_1__70_, fifo_data_o_1__69_, fifo_data_o_1__68_, fifo_data_o_1__67_, fifo_data_o_1__66_, fifo_data_o_1__65_, fifo_data_o_1__64_, fifo_data_o_1__63_, fifo_data_o_1__62_, fifo_data_o_1__61_, fifo_data_o_1__60_, fifo_data_o_1__59_, fifo_data_o_1__58_, fifo_data_o_1__57_, fifo_data_o_1__56_, fifo_data_o_1__55_, fifo_data_o_1__54_, fifo_data_o_1__53_, fifo_data_o_1__52_, fifo_data_o_1__51_, fifo_data_o_1__50_, fifo_data_o_1__49_, fifo_data_o_1__48_, fifo_data_o_1__47_, fifo_data_o_1__46_, fifo_data_o_1__45_, fifo_data_o_1__44_, fifo_data_o_1__43_, fifo_data_o_1__42_, fifo_data_o_1__41_, fifo_data_o_1__40_, fifo_data_o_1__39_, fifo_data_o_1__38_, fifo_data_o_1__37_, fifo_data_o_1__36_, fifo_data_o_1__35_, fifo_data_o_1__34_, fifo_data_o_1__33_, fifo_data_o_1__32_, fifo_data_o_1__31_, fifo_data_o_1__30_, fifo_data_o_1__29_, fifo_data_o_1__28_, fifo_data_o_1__27_, fifo_data_o_1__26_, fifo_data_o_1__25_, fifo_data_o_1__24_, fifo_data_o_1__23_, fifo_data_o_1__22_, fifo_data_o_1__21_, fifo_data_o_1__20_, fifo_data_o_1__19_, fifo_data_o_1__18_, fifo_data_o_1__17_, fifo_data_o_1__16_, fifo_data_o_1__15_, fifo_data_o_1__14_, fifo_data_o_1__13_, fifo_data_o_1__12_, fifo_data_o_1__11_, fifo_data_o_1__10_, fifo_data_o_1__9_, fifo_data_o_1__8_, fifo_data_o_1__7_, fifo_data_o_1__6_, fifo_data_o_1__5_, fifo_data_o_1__4_, fifo_data_o_1__3_, fifo_data_o_1__2_, fifo_data_o_1__1_, fifo_data_o_1__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_4__3_, arb_sel_o_4__2_, arb_sel_o_4__1_, arb_sel_o_4__0_ }),
    .data_o(data_o[654:524])
  );


  bsg_round_robin_arb_inputs_p5
  rr_arb_proc
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(ready_i[0]),
    .reqs_i({ arb_valid_4__0_, arb_valid_3__0_, arb_valid_2__0_, arb_valid_1__0_, arb_valid_0__0_ }),
    .grants_o({ arb_grants_o_4__0_, arb_grants_o_3__0_, arb_grants_o_2__0_, arb_grants_o_1__0_, arb_grants_o_0__0_ }),
    .sel_one_hot_o({ arb_sel_o_0__4_, arb_sel_o_0__3_, arb_sel_o_0__2_, arb_sel_o_0__1_, arb_sel_o_0__0_ }),
    .v_o(valid_o[0]),
    .tag_o({ SV2V_UNCONNECTED_9, SV2V_UNCONNECTED_10, SV2V_UNCONNECTED_11 }),
    .yumi_i(n_27_net_)
  );


  bsg_mux_one_hot_width_p131_els_p5
  mux_proc
  (
    .data_i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_o_3__130_, fifo_data_o_3__129_, fifo_data_o_3__128_, fifo_data_o_3__127_, fifo_data_o_3__126_, fifo_data_o_3__125_, fifo_data_o_3__124_, fifo_data_o_3__123_, fifo_data_o_3__122_, fifo_data_o_3__121_, fifo_data_o_3__120_, fifo_data_o_3__119_, fifo_data_o_3__118_, fifo_data_o_3__117_, fifo_data_o_3__116_, fifo_data_o_3__115_, fifo_data_o_3__114_, fifo_data_o_3__113_, fifo_data_o_3__112_, fifo_data_o_3__111_, fifo_data_o_3__110_, fifo_data_o_3__109_, fifo_data_o_3__108_, fifo_data_o_3__107_, fifo_data_o_3__106_, fifo_data_o_3__105_, fifo_data_o_3__104_, fifo_data_o_3__103_, fifo_data_o_3__102_, fifo_data_o_3__101_, fifo_data_o_3__100_, fifo_data_o_3__99_, fifo_data_o_3__98_, fifo_data_o_3__97_, fifo_data_o_3__96_, fifo_data_o_3__95_, fifo_data_o_3__94_, fifo_data_o_3__93_, fifo_data_o_3__92_, fifo_data_o_3__91_, fifo_data_o_3__90_, fifo_data_o_3__89_, fifo_data_o_3__88_, fifo_data_o_3__87_, fifo_data_o_3__86_, fifo_data_o_3__85_, fifo_data_o_3__84_, fifo_data_o_3__83_, fifo_data_o_3__82_, fifo_data_o_3__81_, fifo_data_o_3__80_, fifo_data_o_3__79_, fifo_data_o_3__78_, fifo_data_o_3__77_, fifo_data_o_3__76_, fifo_data_o_3__75_, fifo_data_o_3__74_, fifo_data_o_3__73_, fifo_data_o_3__72_, fifo_data_o_3__71_, fifo_data_o_3__70_, fifo_data_o_3__69_, fifo_data_o_3__68_, fifo_data_o_3__67_, fifo_data_o_3__66_, fifo_data_o_3__65_, fifo_data_o_3__64_, fifo_data_o_3__63_, fifo_data_o_3__62_, fifo_data_o_3__61_, fifo_data_o_3__60_, fifo_data_o_3__59_, fifo_data_o_3__58_, fifo_data_o_3__57_, fifo_data_o_3__56_, fifo_data_o_3__55_, fifo_data_o_3__54_, fifo_data_o_3__53_, fifo_data_o_3__52_, fifo_data_o_3__51_, fifo_data_o_3__50_, fifo_data_o_3__49_, fifo_data_o_3__48_, fifo_data_o_3__47_, fifo_data_o_3__46_, fifo_data_o_3__45_, fifo_data_o_3__44_, fifo_data_o_3__43_, fifo_data_o_3__42_, fifo_data_o_3__41_, fifo_data_o_3__40_, fifo_data_o_3__39_, fifo_data_o_3__38_, fifo_data_o_3__37_, fifo_data_o_3__36_, fifo_data_o_3__35_, fifo_data_o_3__34_, fifo_data_o_3__33_, fifo_data_o_3__32_, fifo_data_o_3__31_, fifo_data_o_3__30_, fifo_data_o_3__29_, fifo_data_o_3__28_, fifo_data_o_3__27_, fifo_data_o_3__26_, fifo_data_o_3__25_, fifo_data_o_3__24_, fifo_data_o_3__23_, fifo_data_o_3__22_, fifo_data_o_3__21_, fifo_data_o_3__20_, fifo_data_o_3__19_, fifo_data_o_3__18_, fifo_data_o_3__17_, fifo_data_o_3__16_, fifo_data_o_3__15_, fifo_data_o_3__14_, fifo_data_o_3__13_, fifo_data_o_3__12_, fifo_data_o_3__11_, fifo_data_o_3__10_, fifo_data_o_3__9_, fifo_data_o_3__8_, fifo_data_o_3__7_, fifo_data_o_3__6_, fifo_data_o_3__5_, fifo_data_o_3__4_, fifo_data_o_3__3_, fifo_data_o_3__2_, fifo_data_o_3__1_, fifo_data_o_3__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, fifo_data_o_1__130_, fifo_data_o_1__129_, fifo_data_o_1__128_, fifo_data_o_1__127_, fifo_data_o_1__126_, fifo_data_o_1__125_, fifo_data_o_1__124_, fifo_data_o_1__123_, fifo_data_o_1__122_, fifo_data_o_1__121_, fifo_data_o_1__120_, fifo_data_o_1__119_, fifo_data_o_1__118_, fifo_data_o_1__117_, fifo_data_o_1__116_, fifo_data_o_1__115_, fifo_data_o_1__114_, fifo_data_o_1__113_, fifo_data_o_1__112_, fifo_data_o_1__111_, fifo_data_o_1__110_, fifo_data_o_1__109_, fifo_data_o_1__108_, fifo_data_o_1__107_, fifo_data_o_1__106_, fifo_data_o_1__105_, fifo_data_o_1__104_, fifo_data_o_1__103_, fifo_data_o_1__102_, fifo_data_o_1__101_, fifo_data_o_1__100_, fifo_data_o_1__99_, fifo_data_o_1__98_, fifo_data_o_1__97_, fifo_data_o_1__96_, fifo_data_o_1__95_, fifo_data_o_1__94_, fifo_data_o_1__93_, fifo_data_o_1__92_, fifo_data_o_1__91_, fifo_data_o_1__90_, fifo_data_o_1__89_, fifo_data_o_1__88_, fifo_data_o_1__87_, fifo_data_o_1__86_, fifo_data_o_1__85_, fifo_data_o_1__84_, fifo_data_o_1__83_, fifo_data_o_1__82_, fifo_data_o_1__81_, fifo_data_o_1__80_, fifo_data_o_1__79_, fifo_data_o_1__78_, fifo_data_o_1__77_, fifo_data_o_1__76_, fifo_data_o_1__75_, fifo_data_o_1__74_, fifo_data_o_1__73_, fifo_data_o_1__72_, fifo_data_o_1__71_, fifo_data_o_1__70_, fifo_data_o_1__69_, fifo_data_o_1__68_, fifo_data_o_1__67_, fifo_data_o_1__66_, fifo_data_o_1__65_, fifo_data_o_1__64_, fifo_data_o_1__63_, fifo_data_o_1__62_, fifo_data_o_1__61_, fifo_data_o_1__60_, fifo_data_o_1__59_, fifo_data_o_1__58_, fifo_data_o_1__57_, fifo_data_o_1__56_, fifo_data_o_1__55_, fifo_data_o_1__54_, fifo_data_o_1__53_, fifo_data_o_1__52_, fifo_data_o_1__51_, fifo_data_o_1__50_, fifo_data_o_1__49_, fifo_data_o_1__48_, fifo_data_o_1__47_, fifo_data_o_1__46_, fifo_data_o_1__45_, fifo_data_o_1__44_, fifo_data_o_1__43_, fifo_data_o_1__42_, fifo_data_o_1__41_, fifo_data_o_1__40_, fifo_data_o_1__39_, fifo_data_o_1__38_, fifo_data_o_1__37_, fifo_data_o_1__36_, fifo_data_o_1__35_, fifo_data_o_1__34_, fifo_data_o_1__33_, fifo_data_o_1__32_, fifo_data_o_1__31_, fifo_data_o_1__30_, fifo_data_o_1__29_, fifo_data_o_1__28_, fifo_data_o_1__27_, fifo_data_o_1__26_, fifo_data_o_1__25_, fifo_data_o_1__24_, fifo_data_o_1__23_, fifo_data_o_1__22_, fifo_data_o_1__21_, fifo_data_o_1__20_, fifo_data_o_1__19_, fifo_data_o_1__18_, fifo_data_o_1__17_, fifo_data_o_1__16_, fifo_data_o_1__15_, fifo_data_o_1__14_, fifo_data_o_1__13_, fifo_data_o_1__12_, fifo_data_o_1__11_, fifo_data_o_1__10_, fifo_data_o_1__9_, fifo_data_o_1__8_, fifo_data_o_1__7_, fifo_data_o_1__6_, fifo_data_o_1__5_, fifo_data_o_1__4_, fifo_data_o_1__3_, fifo_data_o_1__2_, fifo_data_o_1__1_, fifo_data_o_1__0_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }),
    .sel_one_hot_i({ arb_sel_o_0__4_, arb_sel_o_0__3_, arb_sel_o_0__2_, arb_sel_o_0__1_, arb_sel_o_0__0_ }),
    .data_o(data_o[130:0])
  );

  assign N278 = N0 & local_x_cord_i[0];
  assign N0 = ~1'b0;
  assign N279 = 1'b0 & N1;
  assign N1 = ~local_x_cord_i[0];
  assign N283 = N2 & local_y_cord_i[0];
  assign N2 = ~1'b0;
  assign N284 = 1'b0 & N3;
  assign N3 = ~local_y_cord_i[0];
  assign N4 = fifo_data_o_1__1_ ^ local_y_cord_i[0];
  assign N285 = ~N4;
  assign N5 = fifo_data_o_1__0_ ^ local_x_cord_i[0];
  assign N287 = ~N5;
  assign N288 = fifo_data_o_1__0_ & N6;
  assign N6 = ~local_x_cord_i[0];
  assign N291 = N7 & local_y_cord_i[0];
  assign N7 = ~fifo_data_o_1__1_;
  assign N292 = fifo_data_o_1__1_ & N8;
  assign N8 = ~local_y_cord_i[0];
  assign N9 = fifo_data_o_3__1_ ^ local_y_cord_i[0];
  assign N293 = ~N9;
  assign N10 = fifo_data_o_3__0_ ^ local_x_cord_i[0];
  assign N295 = ~N10;
  assign N296 = N11 & local_x_cord_i[0];
  assign N11 = ~fifo_data_o_3__0_;
  assign N297 = fifo_data_o_3__0_ & N12;
  assign N12 = ~local_x_cord_i[0];
  assign N301 = fifo_data_o_3__1_ & N13;
  assign N13 = ~local_y_cord_i[0];
  assign N323 = out_count_r[2] | out_count_r[3];
  assign N324 = ~N323;
  assign N325 = out_count_r[2] | out_count_r[3];
  assign N326 = ~N325;
  assign N327 = out_count_r[2] | out_count_r[3];
  assign N328 = ~N327;
  assign N329 = out_count_r[2] | out_count_r[3];
  assign N330 = ~N329;
  assign N331 = out_count_r[4] | out_count_r[5];
  assign N332 = ~N331;
  assign N333 = out_count_r[4] | out_count_r[5];
  assign N334 = ~N333;
  assign N335 = out_count_r[4] | out_count_r[5];
  assign N336 = ~N335;
  assign N337 = out_count_r[4] | out_count_r[5];
  assign N338 = ~N337;
  assign N339 = out_count_r[6] | out_count_r[7];
  assign N340 = ~N339;
  assign N341 = out_count_r[6] | out_count_r[7];
  assign N342 = ~N341;
  assign N343 = out_count_r[6] | out_count_r[7];
  assign N344 = ~N343;
  assign N345 = out_count_r[6] | out_count_r[7];
  assign N346 = ~N345;
  assign N347 = out_count_r[8] | out_count_r[9];
  assign N348 = ~N347;
  assign N349 = out_count_r[8] | out_count_r[9];
  assign N350 = ~N349;
  assign N351 = out_count_r[8] | out_count_r[9];
  assign N352 = ~N351;
  assign N353 = out_count_r[8] | out_count_r[9];
  assign N354 = ~N353;
  assign N355 = out_count_r[0] | out_count_r[1];
  assign N356 = ~N355;
  assign N357 = out_count_r[0] | out_count_r[1];
  assign N358 = ~N357;
  assign N359 = out_count_r[0] | out_count_r[1];
  assign N360 = ~N359;
  assign N361 = out_count_r[0] | out_count_r[1];
  assign N362 = ~N361;
  assign N363 = out_count_r[0] | out_count_r[1];
  assign N364 = ~N363;
  assign N365 = out_count_r[0] | out_count_r[1];
  assign N366 = out_count_r[2] | out_count_r[3];
  assign N367 = out_count_r[4] | out_count_r[5];
  assign N368 = out_count_r[6] | out_count_r[7];
  assign N369 = out_count_r[8] | out_count_r[9];
  assign N370 = out_count_r[0] | out_count_r[1];
  assign N371 = out_count_r[4] | out_count_r[5];
  assign N372 = out_count_r[6] | out_count_r[7];
  assign N373 = out_count_r[8] | out_count_r[9];
  assign N374 = out_count_r[0] | out_count_r[1];
  assign N375 = out_count_r[2] | out_count_r[3];
  assign N376 = out_count_r[6] | out_count_r[7];
  assign N377 = out_count_r[8] | out_count_r[9];
  assign N378 = out_count_r[0] | out_count_r[1];
  assign N379 = out_count_r[2] | out_count_r[3];
  assign N380 = out_count_r[4] | out_count_r[5];
  assign N381 = out_count_r[8] | out_count_r[9];
  assign N382 = out_count_r[0] | out_count_r[1];
  assign N383 = out_count_r[2] | out_count_r[3];
  assign N384 = out_count_r[4] | out_count_r[5];
  assign N385 = out_count_r[6] | out_count_r[7];
  assign N386 = count_r[8] | count_r[9];
  assign N387 = ~N386;
  assign N388 = count_r[6] | count_r[7];
  assign N389 = ~N388;
  assign N390 = count_r[4] | count_r[5];
  assign N391 = ~N390;
  assign N392 = count_r[2] | count_r[3];
  assign N393 = ~N392;
  assign N394 = count_r[0] | count_r[1];
  assign N395 = ~N394;
  assign N396 = ~local_y_cord_i[0];
  assign N397 = ~local_x_cord_i[0];
  assign N398 = count_r[0] | count_r[1];
  assign N399 = ~N398;
  assign N400 = count_r[2] | count_r[3];
  assign N401 = ~N400;
  assign N402 = count_r[4] | count_r[5];
  assign N403 = ~N402;
  assign N404 = count_r[6] | count_r[7];
  assign N405 = ~N404;
  assign N406 = count_r[8] | count_r[9];
  assign N407 = ~N406;
  assign N408 = out_count_r[0] | out_count_r[1];
  assign N409 = ~N408;
  assign N410 = out_count_r[2] | out_count_r[3];
  assign N411 = ~N410;
  assign N412 = out_count_r[4] | out_count_r[5];
  assign N413 = ~N412;
  assign N414 = out_count_r[6] | out_count_r[7];
  assign N415 = ~N414;
  assign N416 = out_count_r[8] | out_count_r[9];
  assign N417 = ~N416;
  assign { N126, N125 } = count_r[1:0] - 1'b1;
  assign { N140, N139 } = count_r[3:2] - 1'b1;
  assign { N153, N152 } = count_r[5:4] - 1'b1;
  assign { N167, N166 } = count_r[7:6] - 1'b1;
  assign { N180, N179 } = count_r[9:8] - 1'b1;
  assign { N194, N193 } = out_count_r[1:0] - 1'b1;
  assign { N208, N207 } = out_count_r[3:2] - 1'b1;
  assign { N222, N221 } = out_count_r[5:4] - 1'b1;
  assign { N236, N235 } = out_count_r[7:6] - 1'b1;
  assign { N250, N249 } = out_count_r[9:8] - 1'b1;
  assign { N128, N127 } = (N14)? { 1'b0, 1'b0 } :
                          (N15)? { N126, N125 } : 1'b0;
  assign N14 = N399;
  assign N15 = N398;
  assign { N130, N129 } = (N16)? { N128, N127 } :
                          (N123)? count_r[1:0] : 1'b0;
  assign N16 = fifo_yumi_i[0];
  assign { N132, N131 } = (N17)? { 1'b0, 1'b0 } :
                          (N18)? { N130, N129 } : 1'b0;
  assign N17 = N121;
  assign N18 = N120;
  assign { N142, N141 } = (N19)? { fifo_data_o_1__3_, fifo_data_o_1__2_ } :
                          (N20)? { N140, N139 } : 1'b0;
  assign N19 = N401;
  assign N20 = N400;
  assign { N144, N143 } = (N21)? { N142, N141 } :
                          (N137)? count_r[3:2] : 1'b0;
  assign N21 = N136;
  assign { N146, N145 } = (N22)? { 1'b0, 1'b0 } :
                          (N23)? { N144, N143 } : 1'b0;
  assign N22 = N134;
  assign N23 = N133;
  assign { N155, N154 } = (N24)? { 1'b0, 1'b0 } :
                          (N25)? { N153, N152 } : 1'b0;
  assign N24 = N403;
  assign N25 = N402;
  assign { N157, N156 } = (N26)? { N155, N154 } :
                          (N150)? count_r[5:4] : 1'b0;
  assign N26 = fifo_yumi_i[2];
  assign { N159, N158 } = (N27)? { 1'b0, 1'b0 } :
                          (N28)? { N157, N156 } : 1'b0;
  assign N27 = N148;
  assign N28 = N147;
  assign { N169, N168 } = (N29)? { fifo_data_o_3__3_, fifo_data_o_3__2_ } :
                          (N30)? { N167, N166 } : 1'b0;
  assign N29 = N405;
  assign N30 = N404;
  assign { N171, N170 } = (N31)? { N169, N168 } :
                          (N164)? count_r[7:6] : 1'b0;
  assign N31 = N163;
  assign { N173, N172 } = (N32)? { 1'b0, 1'b0 } :
                          (N33)? { N171, N170 } : 1'b0;
  assign N32 = N161;
  assign N33 = N160;
  assign { N182, N181 } = (N34)? { 1'b0, 1'b0 } :
                          (N35)? { N180, N179 } : 1'b0;
  assign N34 = N407;
  assign N35 = N406;
  assign { N184, N183 } = (N36)? { N182, N181 } :
                          (N177)? count_r[9:8] : 1'b0;
  assign N36 = fifo_yumi_i[4];
  assign { N186, N185 } = (N37)? { 1'b0, 1'b0 } :
                          (N38)? { N184, N183 } : 1'b0;
  assign N37 = N175;
  assign N38 = N174;
  assign { N196, N195 } = (N39)? data_o[3:2] :
                          (N40)? { N194, N193 } : 1'b0;
  assign N39 = N409;
  assign N40 = N408;
  assign { N198, N197 } = (N41)? { N196, N195 } :
                          (N191)? out_count_r[1:0] : 1'b0;
  assign N41 = N190;
  assign { N200, N199 } = (N42)? { 1'b0, 1'b0 } :
                          (N43)? { N198, N197 } : 1'b0;
  assign N42 = N188;
  assign N43 = N187;
  assign { N210, N209 } = (N44)? data_o[134:133] :
                          (N45)? { N208, N207 } : 1'b0;
  assign N44 = N411;
  assign N45 = N410;
  assign { N212, N211 } = (N46)? { N210, N209 } :
                          (N205)? out_count_r[3:2] : 1'b0;
  assign N46 = N204;
  assign { N214, N213 } = (N47)? { 1'b0, 1'b0 } :
                          (N48)? { N212, N211 } : 1'b0;
  assign N47 = N202;
  assign N48 = N201;
  assign { N224, N223 } = (N49)? data_o[265:264] :
                          (N50)? { N222, N221 } : 1'b0;
  assign N49 = N413;
  assign N50 = N412;
  assign { N226, N225 } = (N51)? { N224, N223 } :
                          (N219)? out_count_r[5:4] : 1'b0;
  assign N51 = N218;
  assign { N228, N227 } = (N52)? { 1'b0, 1'b0 } :
                          (N53)? { N226, N225 } : 1'b0;
  assign N52 = N216;
  assign N53 = N215;
  assign { N238, N237 } = (N54)? data_o[396:395] :
                          (N55)? { N236, N235 } : 1'b0;
  assign N54 = N415;
  assign N55 = N414;
  assign { N240, N239 } = (N56)? { N238, N237 } :
                          (N233)? out_count_r[7:6] : 1'b0;
  assign N56 = N232;
  assign { N242, N241 } = (N57)? { 1'b0, 1'b0 } :
                          (N58)? { N240, N239 } : 1'b0;
  assign N57 = N230;
  assign N58 = N229;
  assign { N252, N251 } = (N59)? data_o[527:526] :
                          (N60)? { N250, N249 } : 1'b0;
  assign N59 = N417;
  assign N60 = N416;
  assign { N254, N253 } = (N61)? { N252, N251 } :
                          (N247)? out_count_r[9:8] : 1'b0;
  assign N61 = N246;
  assign { N256, N255 } = (N62)? { 1'b0, 1'b0 } :
                          (N63)? { N254, N253 } : 1'b0;
  assign N62 = N244;
  assign N63 = N243;
  assign arb_valid_0__0_ = (N64)? new_valid_0__0_ :
                           (N65)? N257 : 1'b0;
  assign N64 = N364;
  assign N65 = N363;
  assign arb_valid_0__1_ = (N66)? new_valid_0__1_ :
                           (N67)? N258 : 1'b0;
  assign N66 = N330;
  assign N67 = N329;
  assign arb_valid_0__2_ = (N68)? new_valid_0__2_ :
                           (N69)? N259 : 1'b0;
  assign N68 = N338;
  assign N69 = N337;
  assign arb_valid_0__3_ = (N70)? new_valid_0__3_ :
                           (N71)? N260 : 1'b0;
  assign N70 = N346;
  assign N71 = N345;
  assign arb_valid_0__4_ = (N72)? new_valid_0__4_ :
                           (N73)? N261 : 1'b0;
  assign N72 = N354;
  assign N73 = N353;
  assign arb_valid_1__0_ = (N74)? new_valid_1__0_ :
                           (N75)? N262 : 1'b0;
  assign N74 = N362;
  assign N75 = N361;
  assign arb_valid_1__2_ = (N76)? new_valid_1__2_ :
                           (N77)? N263 : 1'b0;
  assign N76 = N336;
  assign N77 = N335;
  assign arb_valid_1__3_ = (N78)? new_valid_1__3_ :
                           (N79)? N264 : 1'b0;
  assign N78 = N344;
  assign N79 = N343;
  assign arb_valid_1__4_ = (N80)? new_valid_1__4_ :
                           (N81)? N265 : 1'b0;
  assign N80 = N352;
  assign N81 = N351;
  assign arb_valid_2__0_ = (N82)? new_valid_2__0_ :
                           (N83)? N266 : 1'b0;
  assign N82 = N360;
  assign N83 = N359;
  assign arb_valid_2__1_ = (N84)? new_valid_2__1_ :
                           (N85)? N267 : 1'b0;
  assign N84 = N328;
  assign N85 = N327;
  assign arb_valid_2__3_ = (N86)? new_valid_2__3_ :
                           (N87)? N268 : 1'b0;
  assign N86 = N342;
  assign N87 = N341;
  assign arb_valid_2__4_ = (N88)? new_valid_2__4_ :
                           (N89)? N269 : 1'b0;
  assign N88 = N350;
  assign N89 = N349;
  assign arb_valid_3__0_ = (N90)? new_valid_3__0_ :
                           (N91)? N270 : 1'b0;
  assign N90 = N358;
  assign N91 = N357;
  assign arb_valid_3__1_ = (N92)? new_valid_3__1_ :
                           (N93)? N271 : 1'b0;
  assign N92 = N326;
  assign N93 = N325;
  assign arb_valid_3__2_ = (N94)? new_valid_3__2_ :
                           (N95)? N272 : 1'b0;
  assign N94 = N334;
  assign N95 = N333;
  assign arb_valid_3__4_ = (N96)? new_valid_3__4_ :
                           (N97)? N273 : 1'b0;
  assign N96 = N348;
  assign N97 = N347;
  assign arb_valid_4__0_ = (N98)? new_valid_4__0_ :
                           (N99)? N274 : 1'b0;
  assign N98 = N356;
  assign N99 = N355;
  assign arb_valid_4__1_ = (N100)? new_valid_4__1_ :
                           (N101)? N275 : 1'b0;
  assign N100 = N324;
  assign N101 = N323;
  assign arb_valid_4__2_ = (N102)? new_valid_4__2_ :
                           (N103)? N276 : 1'b0;
  assign N102 = N332;
  assign N103 = N331;
  assign arb_valid_4__3_ = (N104)? new_valid_4__3_ :
                           (N105)? N277 : 1'b0;
  assign N104 = N340;
  assign N105 = N339;
  assign { N282, N281, N280 } = (N106)? { N279, N278, N397 } :
                                (N107)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N106 = N396;
  assign N107 = local_y_cord_i[0];
  assign { dest_n_0__4_, dest_n_0__3_, dest_n_0__2_, dest_n_0__1_, dest_n_0__0_ } = (N108)? { N284, N283, N282, N281, N280 } :
                                                                                    (N109)? { dest_r_0__4_, dest_r_0__3_, dest_r_0__2_, dest_r_0__1_, dest_r_0__0_ } : 1'b0;
  assign N108 = N395;
  assign N109 = N394;
  assign { N290, N289 } = (N110)? { N288, N287 } :
                          (N286)? { 1'b0, 1'b0 } : 1'b0;
  assign N110 = N285;
  assign { dest_n_1__4_, dest_n_1__3_, dest_n_1__2_, dest_n_1__0_ } = (N111)? { N292, N291, N290, N289 } :
                                                                      (N112)? { dest_r_1__4_, dest_r_1__3_, dest_r_1__2_, dest_r_1__0_ } : 1'b0;
  assign N111 = N393;
  assign N112 = N392;
  assign { dest_n_2__4_, dest_n_2__3_, dest_n_2__1_, dest_n_2__0_ } = (N113)? { N284, N283, N281, N280 } :
                                                                      (N114)? { dest_r_2__4_, dest_r_2__3_, dest_r_2__1_, dest_r_2__0_ } : 1'b0;
  assign N113 = N391;
  assign N114 = N390;
  assign { N300, N299, N298 } = (N115)? { N297, N296, N295 } :
                                (N294)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N115 = N293;
  assign { dest_n_3__4_, dest_n_3__2_, dest_n_3__1_, dest_n_3__0_ } = (N116)? { N301, N300, N299, N298 } :
                                                                      (N117)? { dest_r_3__4_, dest_r_3__2_, dest_r_3__1_, dest_r_3__0_ } : 1'b0;
  assign N116 = N389;
  assign N117 = N388;
  assign { dest_n_4__3_, dest_n_4__2_, dest_n_4__1_, dest_n_4__0_ } = (N118)? { N283, N282, N281, N280 } :
                                                                      (N119)? { dest_r_4__3_, dest_r_4__2_, dest_r_4__1_, dest_r_4__0_ } : 1'b0;
  assign N118 = N387;
  assign N119 = N386;
  assign N120 = ~reset_i;
  assign N121 = reset_i;
  assign N122 = N120;
  assign N123 = ~fifo_yumi_i[0];
  assign N124 = N122 & fifo_yumi_i[0];
  assign N133 = ~reset_i;
  assign N134 = reset_i;
  assign N135 = N133;
  assign N136 = fifo_yumi_i[1];
  assign N137 = ~N136;
  assign N138 = N135 & N136;
  assign N147 = ~reset_i;
  assign N148 = reset_i;
  assign N149 = N147;
  assign N150 = ~fifo_yumi_i[2];
  assign N151 = N149 & fifo_yumi_i[2];
  assign N160 = ~reset_i;
  assign N161 = reset_i;
  assign N162 = N160;
  assign N163 = fifo_yumi_i[3];
  assign N164 = ~N163;
  assign N165 = N162 & N163;
  assign N174 = ~reset_i;
  assign N175 = reset_i;
  assign N176 = N174;
  assign N177 = ~fifo_yumi_i[4];
  assign N178 = N176 & fifo_yumi_i[4];
  assign new_valid_0__0_ = 1'b0 & dest_n_0__0_;
  assign new_valid_0__1_ = 1'b0 & dest_n_0__1_;
  assign new_valid_0__2_ = 1'b0 & dest_n_0__2_;
  assign new_valid_0__3_ = 1'b0 & dest_n_0__3_;
  assign new_valid_0__4_ = 1'b0 & dest_n_0__4_;
  assign new_valid_1__0_ = fifo_valid_o_1 & dest_n_1__0_;
  assign new_valid_1__2_ = fifo_valid_o_1 & dest_n_1__2_;
  assign new_valid_1__3_ = fifo_valid_o_1 & dest_n_1__3_;
  assign new_valid_1__4_ = fifo_valid_o_1 & dest_n_1__4_;
  assign new_valid_2__0_ = 1'b0 & dest_n_2__0_;
  assign new_valid_2__1_ = 1'b0 & dest_n_2__1_;
  assign new_valid_2__3_ = 1'b0 & dest_n_2__3_;
  assign new_valid_2__4_ = 1'b0 & dest_n_2__4_;
  assign new_valid_3__0_ = fifo_valid_o[3] & dest_n_3__0_;
  assign new_valid_3__1_ = fifo_valid_o[3] & dest_n_3__1_;
  assign new_valid_3__2_ = fifo_valid_o[3] & dest_n_3__2_;
  assign new_valid_3__4_ = fifo_valid_o[3] & dest_n_3__4_;
  assign new_valid_4__0_ = 1'b0 & dest_n_4__0_;
  assign new_valid_4__1_ = 1'b0 & dest_n_4__1_;
  assign new_valid_4__2_ = 1'b0 & dest_n_4__2_;
  assign new_valid_4__3_ = 1'b0 & dest_n_4__3_;
  assign fifo_yumi_i[0] = N420 | arb_grants_o_0__0_;
  assign N420 = N419 | arb_grants_o_0__1_;
  assign N419 = N418 | arb_grants_o_0__2_;
  assign N418 = arb_grants_o_0__4_ | arb_grants_o_0__3_;
  assign fifo_yumi_i[1] = N423 | arb_grants_o_1__0_;
  assign N423 = N422 | 1'b0;
  assign N422 = N421 | arb_grants_o_1__2_;
  assign N421 = arb_grants_o_1__4_ | arb_grants_o_1__3_;
  assign fifo_yumi_i[2] = N426 | arb_grants_o_2__0_;
  assign N426 = N425 | arb_grants_o_2__1_;
  assign N425 = N424 | 1'b0;
  assign N424 = arb_grants_o_2__4_ | arb_grants_o_2__3_;
  assign fifo_yumi_i[3] = N429 | arb_grants_o_3__0_;
  assign N429 = N428 | arb_grants_o_3__1_;
  assign N428 = N427 | arb_grants_o_3__2_;
  assign N427 = arb_grants_o_3__4_ | 1'b0;
  assign fifo_yumi_i[4] = N432 | arb_grants_o_4__0_;
  assign N432 = N431 | arb_grants_o_4__1_;
  assign N431 = N430 | arb_grants_o_4__2_;
  assign N430 = 1'b0 | arb_grants_o_4__3_;
  assign N187 = ~reset_i;
  assign N188 = reset_i;
  assign N189 = N187;
  assign N190 = valid_o[0] & ready_i[0];
  assign N191 = ~N190;
  assign N192 = N189 & N190;
  assign N201 = ~reset_i;
  assign N202 = reset_i;
  assign N203 = N201;
  assign N204 = valid_o[1] & ready_i[1];
  assign N205 = ~N204;
  assign N206 = N203 & N204;
  assign N215 = ~reset_i;
  assign N216 = reset_i;
  assign N217 = N215;
  assign N218 = valid_o[2] & 1'b1;
  assign N219 = ~N218;
  assign N220 = N217 & N218;
  assign N229 = ~reset_i;
  assign N230 = reset_i;
  assign N231 = N229;
  assign N232 = valid_o[3] & 1'b1;
  assign N233 = ~N232;
  assign N234 = N231 & N232;
  assign N243 = ~reset_i;
  assign N244 = reset_i;
  assign N245 = N243;
  assign N246 = valid_o[4] & 1'b1;
  assign N247 = ~N246;
  assign N248 = N245 & N246;
  assign N257 = new_valid_0__0_ & arb_grants_r_0__0_;
  assign N258 = new_valid_0__1_ & arb_grants_r_0__1_;
  assign N259 = new_valid_0__2_ & arb_grants_r_0__2_;
  assign N260 = new_valid_0__3_ & arb_grants_r_0__3_;
  assign N261 = new_valid_0__4_ & arb_grants_r_0__4_;
  assign N262 = new_valid_1__0_ & arb_grants_r_1__0_;
  assign N263 = new_valid_1__2_ & arb_grants_r_1__2_;
  assign N264 = new_valid_1__3_ & arb_grants_r_1__3_;
  assign N265 = new_valid_1__4_ & arb_grants_r_1__4_;
  assign N266 = new_valid_2__0_ & arb_grants_r_2__0_;
  assign N267 = new_valid_2__1_ & arb_grants_r_2__1_;
  assign N268 = new_valid_2__3_ & arb_grants_r_2__3_;
  assign N269 = new_valid_2__4_ & arb_grants_r_2__4_;
  assign N270 = new_valid_3__0_ & arb_grants_r_3__0_;
  assign N271 = new_valid_3__1_ & arb_grants_r_3__1_;
  assign N272 = new_valid_3__2_ & arb_grants_r_3__2_;
  assign N273 = new_valid_3__4_ & arb_grants_r_3__4_;
  assign N274 = new_valid_4__0_ & arb_grants_r_4__0_;
  assign N275 = new_valid_4__1_ & arb_grants_r_4__1_;
  assign N276 = new_valid_4__2_ & arb_grants_r_4__2_;
  assign N277 = new_valid_4__3_ & arb_grants_r_4__3_;
  assign n_3_net_ = valid_o[1] & ready_i[1];
  assign n_9_net_ = valid_o[2] & 1'b1;
  assign n_15_net_ = valid_o[3] & 1'b1;
  assign n_21_net_ = valid_o[4] & 1'b1;
  assign n_27_net_ = valid_o[0] & ready_i[0];
  assign N286 = ~N285;
  assign N294 = ~N293;
  assign N302 = ~N365;
  assign N303 = ~N366;
  assign N304 = ~N367;
  assign N305 = ~N368;
  assign N306 = ~N369;
  assign N307 = ~N370;
  assign N308 = ~N371;
  assign N309 = ~N372;
  assign N310 = ~N373;
  assign N311 = ~N374;
  assign N312 = ~N375;
  assign N313 = ~N376;
  assign N314 = ~N377;
  assign N315 = ~N378;
  assign N316 = ~N379;
  assign N317 = ~N380;
  assign N318 = ~N381;
  assign N319 = ~N382;
  assign N320 = ~N383;
  assign N321 = ~N384;
  assign N322 = ~N385;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { count_r[9:0] } <= { N186, N185, N173, N172, N159, N158, N146, N145, N132, N131 };
      dest_r_0__4_ <= dest_n_0__4_;
      dest_r_0__3_ <= dest_n_0__3_;
      dest_r_0__2_ <= dest_n_0__2_;
      dest_r_0__1_ <= dest_n_0__1_;
      dest_r_0__0_ <= dest_n_0__0_;
      dest_r_1__4_ <= dest_n_1__4_;
      dest_r_1__3_ <= dest_n_1__3_;
      dest_r_1__2_ <= dest_n_1__2_;
      dest_r_1__0_ <= dest_n_1__0_;
      dest_r_2__4_ <= dest_n_2__4_;
      dest_r_2__3_ <= dest_n_2__3_;
      dest_r_2__1_ <= dest_n_2__1_;
      dest_r_2__0_ <= dest_n_2__0_;
      dest_r_3__4_ <= dest_n_3__4_;
      dest_r_3__2_ <= dest_n_3__2_;
      dest_r_3__1_ <= dest_n_3__1_;
      dest_r_3__0_ <= dest_n_3__0_;
      dest_r_4__3_ <= dest_n_4__3_;
      dest_r_4__2_ <= dest_n_4__2_;
      dest_r_4__1_ <= dest_n_4__1_;
      dest_r_4__0_ <= dest_n_4__0_;
      { out_count_r[9:0] } <= { N256, N255, N242, N241, N228, N227, N214, N213, N200, N199 };
    end
    if(N302) begin
      arb_grants_r_0__0_ <= arb_grants_o_0__0_;
    end
    if(N303) begin
      arb_grants_r_0__1_ <= arb_grants_o_0__1_;
    end
    if(N304) begin
      arb_grants_r_0__2_ <= arb_grants_o_0__2_;
    end
    if(N305) begin
      arb_grants_r_0__3_ <= arb_grants_o_0__3_;
    end
    if(N306) begin
      arb_grants_r_0__4_ <= arb_grants_o_0__4_;
    end
    if(N307) begin
      arb_grants_r_1__0_ <= arb_grants_o_1__0_;
    end
    if(N308) begin
      arb_grants_r_1__2_ <= arb_grants_o_1__2_;
    end
    if(N309) begin
      arb_grants_r_1__3_ <= arb_grants_o_1__3_;
    end
    if(N310) begin
      arb_grants_r_1__4_ <= arb_grants_o_1__4_;
    end
    if(N311) begin
      arb_grants_r_2__0_ <= arb_grants_o_2__0_;
    end
    if(N312) begin
      arb_grants_r_2__1_ <= arb_grants_o_2__1_;
    end
    if(N313) begin
      arb_grants_r_2__3_ <= arb_grants_o_2__3_;
    end
    if(N314) begin
      arb_grants_r_2__4_ <= arb_grants_o_2__4_;
    end
    if(N315) begin
      arb_grants_r_3__0_ <= arb_grants_o_3__0_;
    end
    if(N316) begin
      arb_grants_r_3__1_ <= arb_grants_o_3__1_;
    end
    if(N317) begin
      arb_grants_r_3__2_ <= arb_grants_o_3__2_;
    end
    if(N318) begin
      arb_grants_r_3__4_ <= arb_grants_o_3__4_;
    end
    if(N319) begin
      arb_grants_r_4__0_ <= arb_grants_o_4__0_;
    end
    if(N320) begin
      arb_grants_r_4__1_ <= arb_grants_o_4__1_;
    end
    if(N321) begin
      arb_grants_r_4__2_ <= arb_grants_o_4__2_;
    end
    if(N322) begin
      arb_grants_r_4__3_ <= arb_grants_o_4__3_;
    end
  end


endmodule



module bp_me_network_pkt_encode_data_cmd_num_lce_p2_lce_assoc_p8_block_size_in_bits_p512_max_num_flit_p4_x_cord_width_p1_y_cord_width_p1
(
  payload_i,
  packet_o
);

  input [517:0] payload_i;
  output [521:0] packet_o;
  wire [521:0] packet_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11;
  assign packet_o[1] = 1'b1;
  assign packet_o[521] = payload_i[517];
  assign packet_o[520] = payload_i[516];
  assign packet_o[519] = payload_i[515];
  assign packet_o[518] = payload_i[514];
  assign packet_o[517] = payload_i[513];
  assign packet_o[516] = payload_i[512];
  assign packet_o[515] = payload_i[511];
  assign packet_o[514] = payload_i[510];
  assign packet_o[513] = payload_i[509];
  assign packet_o[512] = payload_i[508];
  assign packet_o[511] = payload_i[507];
  assign packet_o[510] = payload_i[506];
  assign packet_o[509] = payload_i[505];
  assign packet_o[508] = payload_i[504];
  assign packet_o[507] = payload_i[503];
  assign packet_o[506] = payload_i[502];
  assign packet_o[505] = payload_i[501];
  assign packet_o[504] = payload_i[500];
  assign packet_o[503] = payload_i[499];
  assign packet_o[502] = payload_i[498];
  assign packet_o[501] = payload_i[497];
  assign packet_o[500] = payload_i[496];
  assign packet_o[499] = payload_i[495];
  assign packet_o[498] = payload_i[494];
  assign packet_o[497] = payload_i[493];
  assign packet_o[496] = payload_i[492];
  assign packet_o[495] = payload_i[491];
  assign packet_o[494] = payload_i[490];
  assign packet_o[493] = payload_i[489];
  assign packet_o[492] = payload_i[488];
  assign packet_o[491] = payload_i[487];
  assign packet_o[490] = payload_i[486];
  assign packet_o[489] = payload_i[485];
  assign packet_o[488] = payload_i[484];
  assign packet_o[487] = payload_i[483];
  assign packet_o[486] = payload_i[482];
  assign packet_o[485] = payload_i[481];
  assign packet_o[484] = payload_i[480];
  assign packet_o[483] = payload_i[479];
  assign packet_o[482] = payload_i[478];
  assign packet_o[481] = payload_i[477];
  assign packet_o[480] = payload_i[476];
  assign packet_o[479] = payload_i[475];
  assign packet_o[478] = payload_i[474];
  assign packet_o[477] = payload_i[473];
  assign packet_o[476] = payload_i[472];
  assign packet_o[475] = payload_i[471];
  assign packet_o[474] = payload_i[470];
  assign packet_o[473] = payload_i[469];
  assign packet_o[472] = payload_i[468];
  assign packet_o[471] = payload_i[467];
  assign packet_o[470] = payload_i[466];
  assign packet_o[469] = payload_i[465];
  assign packet_o[468] = payload_i[464];
  assign packet_o[467] = payload_i[463];
  assign packet_o[466] = payload_i[462];
  assign packet_o[465] = payload_i[461];
  assign packet_o[464] = payload_i[460];
  assign packet_o[463] = payload_i[459];
  assign packet_o[462] = payload_i[458];
  assign packet_o[461] = payload_i[457];
  assign packet_o[460] = payload_i[456];
  assign packet_o[459] = payload_i[455];
  assign packet_o[458] = payload_i[454];
  assign packet_o[457] = payload_i[453];
  assign packet_o[456] = payload_i[452];
  assign packet_o[455] = payload_i[451];
  assign packet_o[454] = payload_i[450];
  assign packet_o[453] = payload_i[449];
  assign packet_o[452] = payload_i[448];
  assign packet_o[451] = payload_i[447];
  assign packet_o[450] = payload_i[446];
  assign packet_o[449] = payload_i[445];
  assign packet_o[448] = payload_i[444];
  assign packet_o[447] = payload_i[443];
  assign packet_o[446] = payload_i[442];
  assign packet_o[445] = payload_i[441];
  assign packet_o[444] = payload_i[440];
  assign packet_o[443] = payload_i[439];
  assign packet_o[442] = payload_i[438];
  assign packet_o[441] = payload_i[437];
  assign packet_o[440] = payload_i[436];
  assign packet_o[439] = payload_i[435];
  assign packet_o[438] = payload_i[434];
  assign packet_o[437] = payload_i[433];
  assign packet_o[436] = payload_i[432];
  assign packet_o[435] = payload_i[431];
  assign packet_o[434] = payload_i[430];
  assign packet_o[433] = payload_i[429];
  assign packet_o[432] = payload_i[428];
  assign packet_o[431] = payload_i[427];
  assign packet_o[430] = payload_i[426];
  assign packet_o[429] = payload_i[425];
  assign packet_o[428] = payload_i[424];
  assign packet_o[427] = payload_i[423];
  assign packet_o[426] = payload_i[422];
  assign packet_o[425] = payload_i[421];
  assign packet_o[424] = payload_i[420];
  assign packet_o[423] = payload_i[419];
  assign packet_o[422] = payload_i[418];
  assign packet_o[421] = payload_i[417];
  assign packet_o[420] = payload_i[416];
  assign packet_o[419] = payload_i[415];
  assign packet_o[418] = payload_i[414];
  assign packet_o[417] = payload_i[413];
  assign packet_o[416] = payload_i[412];
  assign packet_o[415] = payload_i[411];
  assign packet_o[414] = payload_i[410];
  assign packet_o[413] = payload_i[409];
  assign packet_o[412] = payload_i[408];
  assign packet_o[411] = payload_i[407];
  assign packet_o[410] = payload_i[406];
  assign packet_o[409] = payload_i[405];
  assign packet_o[408] = payload_i[404];
  assign packet_o[407] = payload_i[403];
  assign packet_o[406] = payload_i[402];
  assign packet_o[405] = payload_i[401];
  assign packet_o[404] = payload_i[400];
  assign packet_o[403] = payload_i[399];
  assign packet_o[402] = payload_i[398];
  assign packet_o[401] = payload_i[397];
  assign packet_o[400] = payload_i[396];
  assign packet_o[399] = payload_i[395];
  assign packet_o[398] = payload_i[394];
  assign packet_o[397] = payload_i[393];
  assign packet_o[396] = payload_i[392];
  assign packet_o[395] = payload_i[391];
  assign packet_o[394] = payload_i[390];
  assign packet_o[393] = payload_i[389];
  assign packet_o[392] = payload_i[388];
  assign packet_o[391] = payload_i[387];
  assign packet_o[390] = payload_i[386];
  assign packet_o[389] = payload_i[385];
  assign packet_o[388] = payload_i[384];
  assign packet_o[387] = payload_i[383];
  assign packet_o[386] = payload_i[382];
  assign packet_o[385] = payload_i[381];
  assign packet_o[384] = payload_i[380];
  assign packet_o[383] = payload_i[379];
  assign packet_o[382] = payload_i[378];
  assign packet_o[381] = payload_i[377];
  assign packet_o[380] = payload_i[376];
  assign packet_o[379] = payload_i[375];
  assign packet_o[378] = payload_i[374];
  assign packet_o[377] = payload_i[373];
  assign packet_o[376] = payload_i[372];
  assign packet_o[375] = payload_i[371];
  assign packet_o[374] = payload_i[370];
  assign packet_o[373] = payload_i[369];
  assign packet_o[372] = payload_i[368];
  assign packet_o[371] = payload_i[367];
  assign packet_o[370] = payload_i[366];
  assign packet_o[369] = payload_i[365];
  assign packet_o[368] = payload_i[364];
  assign packet_o[367] = payload_i[363];
  assign packet_o[366] = payload_i[362];
  assign packet_o[365] = payload_i[361];
  assign packet_o[364] = payload_i[360];
  assign packet_o[363] = payload_i[359];
  assign packet_o[362] = payload_i[358];
  assign packet_o[361] = payload_i[357];
  assign packet_o[360] = payload_i[356];
  assign packet_o[359] = payload_i[355];
  assign packet_o[358] = payload_i[354];
  assign packet_o[357] = payload_i[353];
  assign packet_o[356] = payload_i[352];
  assign packet_o[355] = payload_i[351];
  assign packet_o[354] = payload_i[350];
  assign packet_o[353] = payload_i[349];
  assign packet_o[352] = payload_i[348];
  assign packet_o[351] = payload_i[347];
  assign packet_o[350] = payload_i[346];
  assign packet_o[349] = payload_i[345];
  assign packet_o[348] = payload_i[344];
  assign packet_o[347] = payload_i[343];
  assign packet_o[346] = payload_i[342];
  assign packet_o[345] = payload_i[341];
  assign packet_o[344] = payload_i[340];
  assign packet_o[343] = payload_i[339];
  assign packet_o[342] = payload_i[338];
  assign packet_o[341] = payload_i[337];
  assign packet_o[340] = payload_i[336];
  assign packet_o[339] = payload_i[335];
  assign packet_o[338] = payload_i[334];
  assign packet_o[337] = payload_i[333];
  assign packet_o[336] = payload_i[332];
  assign packet_o[335] = payload_i[331];
  assign packet_o[334] = payload_i[330];
  assign packet_o[333] = payload_i[329];
  assign packet_o[332] = payload_i[328];
  assign packet_o[331] = payload_i[327];
  assign packet_o[330] = payload_i[326];
  assign packet_o[329] = payload_i[325];
  assign packet_o[328] = payload_i[324];
  assign packet_o[327] = payload_i[323];
  assign packet_o[326] = payload_i[322];
  assign packet_o[325] = payload_i[321];
  assign packet_o[324] = payload_i[320];
  assign packet_o[323] = payload_i[319];
  assign packet_o[322] = payload_i[318];
  assign packet_o[321] = payload_i[317];
  assign packet_o[320] = payload_i[316];
  assign packet_o[319] = payload_i[315];
  assign packet_o[318] = payload_i[314];
  assign packet_o[317] = payload_i[313];
  assign packet_o[316] = payload_i[312];
  assign packet_o[315] = payload_i[311];
  assign packet_o[314] = payload_i[310];
  assign packet_o[313] = payload_i[309];
  assign packet_o[312] = payload_i[308];
  assign packet_o[311] = payload_i[307];
  assign packet_o[310] = payload_i[306];
  assign packet_o[309] = payload_i[305];
  assign packet_o[308] = payload_i[304];
  assign packet_o[307] = payload_i[303];
  assign packet_o[306] = payload_i[302];
  assign packet_o[305] = payload_i[301];
  assign packet_o[304] = payload_i[300];
  assign packet_o[303] = payload_i[299];
  assign packet_o[302] = payload_i[298];
  assign packet_o[301] = payload_i[297];
  assign packet_o[300] = payload_i[296];
  assign packet_o[299] = payload_i[295];
  assign packet_o[298] = payload_i[294];
  assign packet_o[297] = payload_i[293];
  assign packet_o[296] = payload_i[292];
  assign packet_o[295] = payload_i[291];
  assign packet_o[294] = payload_i[290];
  assign packet_o[293] = payload_i[289];
  assign packet_o[292] = payload_i[288];
  assign packet_o[291] = payload_i[287];
  assign packet_o[290] = payload_i[286];
  assign packet_o[289] = payload_i[285];
  assign packet_o[288] = payload_i[284];
  assign packet_o[287] = payload_i[283];
  assign packet_o[286] = payload_i[282];
  assign packet_o[285] = payload_i[281];
  assign packet_o[284] = payload_i[280];
  assign packet_o[283] = payload_i[279];
  assign packet_o[282] = payload_i[278];
  assign packet_o[281] = payload_i[277];
  assign packet_o[280] = payload_i[276];
  assign packet_o[279] = payload_i[275];
  assign packet_o[278] = payload_i[274];
  assign packet_o[277] = payload_i[273];
  assign packet_o[276] = payload_i[272];
  assign packet_o[275] = payload_i[271];
  assign packet_o[274] = payload_i[270];
  assign packet_o[273] = payload_i[269];
  assign packet_o[272] = payload_i[268];
  assign packet_o[271] = payload_i[267];
  assign packet_o[270] = payload_i[266];
  assign packet_o[269] = payload_i[265];
  assign packet_o[268] = payload_i[264];
  assign packet_o[267] = payload_i[263];
  assign packet_o[266] = payload_i[262];
  assign packet_o[265] = payload_i[261];
  assign packet_o[264] = payload_i[260];
  assign packet_o[263] = payload_i[259];
  assign packet_o[262] = payload_i[258];
  assign packet_o[261] = payload_i[257];
  assign packet_o[260] = payload_i[256];
  assign packet_o[259] = payload_i[255];
  assign packet_o[258] = payload_i[254];
  assign packet_o[257] = payload_i[253];
  assign packet_o[256] = payload_i[252];
  assign packet_o[255] = payload_i[251];
  assign packet_o[254] = payload_i[250];
  assign packet_o[253] = payload_i[249];
  assign packet_o[252] = payload_i[248];
  assign packet_o[251] = payload_i[247];
  assign packet_o[250] = payload_i[246];
  assign packet_o[249] = payload_i[245];
  assign packet_o[248] = payload_i[244];
  assign packet_o[247] = payload_i[243];
  assign packet_o[246] = payload_i[242];
  assign packet_o[245] = payload_i[241];
  assign packet_o[244] = payload_i[240];
  assign packet_o[243] = payload_i[239];
  assign packet_o[242] = payload_i[238];
  assign packet_o[241] = payload_i[237];
  assign packet_o[240] = payload_i[236];
  assign packet_o[239] = payload_i[235];
  assign packet_o[238] = payload_i[234];
  assign packet_o[237] = payload_i[233];
  assign packet_o[236] = payload_i[232];
  assign packet_o[235] = payload_i[231];
  assign packet_o[234] = payload_i[230];
  assign packet_o[233] = payload_i[229];
  assign packet_o[232] = payload_i[228];
  assign packet_o[231] = payload_i[227];
  assign packet_o[230] = payload_i[226];
  assign packet_o[229] = payload_i[225];
  assign packet_o[228] = payload_i[224];
  assign packet_o[227] = payload_i[223];
  assign packet_o[226] = payload_i[222];
  assign packet_o[225] = payload_i[221];
  assign packet_o[224] = payload_i[220];
  assign packet_o[223] = payload_i[219];
  assign packet_o[222] = payload_i[218];
  assign packet_o[221] = payload_i[217];
  assign packet_o[220] = payload_i[216];
  assign packet_o[219] = payload_i[215];
  assign packet_o[218] = payload_i[214];
  assign packet_o[217] = payload_i[213];
  assign packet_o[216] = payload_i[212];
  assign packet_o[215] = payload_i[211];
  assign packet_o[214] = payload_i[210];
  assign packet_o[213] = payload_i[209];
  assign packet_o[212] = payload_i[208];
  assign packet_o[211] = payload_i[207];
  assign packet_o[210] = payload_i[206];
  assign packet_o[209] = payload_i[205];
  assign packet_o[208] = payload_i[204];
  assign packet_o[207] = payload_i[203];
  assign packet_o[206] = payload_i[202];
  assign packet_o[205] = payload_i[201];
  assign packet_o[204] = payload_i[200];
  assign packet_o[203] = payload_i[199];
  assign packet_o[202] = payload_i[198];
  assign packet_o[201] = payload_i[197];
  assign packet_o[200] = payload_i[196];
  assign packet_o[199] = payload_i[195];
  assign packet_o[198] = payload_i[194];
  assign packet_o[197] = payload_i[193];
  assign packet_o[196] = payload_i[192];
  assign packet_o[195] = payload_i[191];
  assign packet_o[194] = payload_i[190];
  assign packet_o[193] = payload_i[189];
  assign packet_o[192] = payload_i[188];
  assign packet_o[191] = payload_i[187];
  assign packet_o[190] = payload_i[186];
  assign packet_o[189] = payload_i[185];
  assign packet_o[188] = payload_i[184];
  assign packet_o[187] = payload_i[183];
  assign packet_o[186] = payload_i[182];
  assign packet_o[185] = payload_i[181];
  assign packet_o[184] = payload_i[180];
  assign packet_o[183] = payload_i[179];
  assign packet_o[182] = payload_i[178];
  assign packet_o[181] = payload_i[177];
  assign packet_o[180] = payload_i[176];
  assign packet_o[179] = payload_i[175];
  assign packet_o[178] = payload_i[174];
  assign packet_o[177] = payload_i[173];
  assign packet_o[176] = payload_i[172];
  assign packet_o[175] = payload_i[171];
  assign packet_o[174] = payload_i[170];
  assign packet_o[173] = payload_i[169];
  assign packet_o[172] = payload_i[168];
  assign packet_o[171] = payload_i[167];
  assign packet_o[170] = payload_i[166];
  assign packet_o[169] = payload_i[165];
  assign packet_o[168] = payload_i[164];
  assign packet_o[167] = payload_i[163];
  assign packet_o[166] = payload_i[162];
  assign packet_o[165] = payload_i[161];
  assign packet_o[164] = payload_i[160];
  assign packet_o[163] = payload_i[159];
  assign packet_o[162] = payload_i[158];
  assign packet_o[161] = payload_i[157];
  assign packet_o[160] = payload_i[156];
  assign packet_o[159] = payload_i[155];
  assign packet_o[158] = payload_i[154];
  assign packet_o[157] = payload_i[153];
  assign packet_o[156] = payload_i[152];
  assign packet_o[155] = payload_i[151];
  assign packet_o[154] = payload_i[150];
  assign packet_o[153] = payload_i[149];
  assign packet_o[152] = payload_i[148];
  assign packet_o[151] = payload_i[147];
  assign packet_o[150] = payload_i[146];
  assign packet_o[149] = payload_i[145];
  assign packet_o[148] = payload_i[144];
  assign packet_o[147] = payload_i[143];
  assign packet_o[146] = payload_i[142];
  assign packet_o[145] = payload_i[141];
  assign packet_o[144] = payload_i[140];
  assign packet_o[143] = payload_i[139];
  assign packet_o[142] = payload_i[138];
  assign packet_o[141] = payload_i[137];
  assign packet_o[140] = payload_i[136];
  assign packet_o[139] = payload_i[135];
  assign packet_o[138] = payload_i[134];
  assign packet_o[137] = payload_i[133];
  assign packet_o[136] = payload_i[132];
  assign packet_o[135] = payload_i[131];
  assign packet_o[134] = payload_i[130];
  assign packet_o[133] = payload_i[129];
  assign packet_o[132] = payload_i[128];
  assign packet_o[131] = payload_i[127];
  assign packet_o[130] = payload_i[126];
  assign packet_o[129] = payload_i[125];
  assign packet_o[128] = payload_i[124];
  assign packet_o[127] = payload_i[123];
  assign packet_o[126] = payload_i[122];
  assign packet_o[125] = payload_i[121];
  assign packet_o[124] = payload_i[120];
  assign packet_o[123] = payload_i[119];
  assign packet_o[122] = payload_i[118];
  assign packet_o[121] = payload_i[117];
  assign packet_o[120] = payload_i[116];
  assign packet_o[119] = payload_i[115];
  assign packet_o[118] = payload_i[114];
  assign packet_o[117] = payload_i[113];
  assign packet_o[116] = payload_i[112];
  assign packet_o[115] = payload_i[111];
  assign packet_o[114] = payload_i[110];
  assign packet_o[113] = payload_i[109];
  assign packet_o[112] = payload_i[108];
  assign packet_o[111] = payload_i[107];
  assign packet_o[110] = payload_i[106];
  assign packet_o[109] = payload_i[105];
  assign packet_o[108] = payload_i[104];
  assign packet_o[107] = payload_i[103];
  assign packet_o[106] = payload_i[102];
  assign packet_o[105] = payload_i[101];
  assign packet_o[104] = payload_i[100];
  assign packet_o[103] = payload_i[99];
  assign packet_o[102] = payload_i[98];
  assign packet_o[101] = payload_i[97];
  assign packet_o[100] = payload_i[96];
  assign packet_o[99] = payload_i[95];
  assign packet_o[98] = payload_i[94];
  assign packet_o[97] = payload_i[93];
  assign packet_o[96] = payload_i[92];
  assign packet_o[95] = payload_i[91];
  assign packet_o[94] = payload_i[90];
  assign packet_o[93] = payload_i[89];
  assign packet_o[92] = payload_i[88];
  assign packet_o[91] = payload_i[87];
  assign packet_o[90] = payload_i[86];
  assign packet_o[89] = payload_i[85];
  assign packet_o[88] = payload_i[84];
  assign packet_o[87] = payload_i[83];
  assign packet_o[86] = payload_i[82];
  assign packet_o[85] = payload_i[81];
  assign packet_o[84] = payload_i[80];
  assign packet_o[83] = payload_i[79];
  assign packet_o[82] = payload_i[78];
  assign packet_o[81] = payload_i[77];
  assign packet_o[80] = payload_i[76];
  assign packet_o[79] = payload_i[75];
  assign packet_o[78] = payload_i[74];
  assign packet_o[77] = payload_i[73];
  assign packet_o[76] = payload_i[72];
  assign packet_o[75] = payload_i[71];
  assign packet_o[74] = payload_i[70];
  assign packet_o[73] = payload_i[69];
  assign packet_o[72] = payload_i[68];
  assign packet_o[71] = payload_i[67];
  assign packet_o[70] = payload_i[66];
  assign packet_o[69] = payload_i[65];
  assign packet_o[68] = payload_i[64];
  assign packet_o[67] = payload_i[63];
  assign packet_o[66] = payload_i[62];
  assign packet_o[65] = payload_i[61];
  assign packet_o[64] = payload_i[60];
  assign packet_o[63] = payload_i[59];
  assign packet_o[62] = payload_i[58];
  assign packet_o[61] = payload_i[57];
  assign packet_o[60] = payload_i[56];
  assign packet_o[59] = payload_i[55];
  assign packet_o[58] = payload_i[54];
  assign packet_o[57] = payload_i[53];
  assign packet_o[56] = payload_i[52];
  assign packet_o[55] = payload_i[51];
  assign packet_o[54] = payload_i[50];
  assign packet_o[53] = payload_i[49];
  assign packet_o[52] = payload_i[48];
  assign packet_o[51] = payload_i[47];
  assign packet_o[50] = payload_i[46];
  assign packet_o[49] = payload_i[45];
  assign packet_o[48] = payload_i[44];
  assign packet_o[47] = payload_i[43];
  assign packet_o[46] = payload_i[42];
  assign packet_o[45] = payload_i[41];
  assign packet_o[44] = payload_i[40];
  assign packet_o[43] = payload_i[39];
  assign packet_o[42] = payload_i[38];
  assign packet_o[41] = payload_i[37];
  assign packet_o[40] = payload_i[36];
  assign packet_o[39] = payload_i[35];
  assign packet_o[38] = payload_i[34];
  assign packet_o[37] = payload_i[33];
  assign packet_o[36] = payload_i[32];
  assign packet_o[35] = payload_i[31];
  assign packet_o[34] = payload_i[30];
  assign packet_o[33] = payload_i[29];
  assign packet_o[32] = payload_i[28];
  assign packet_o[31] = payload_i[27];
  assign packet_o[30] = payload_i[26];
  assign packet_o[29] = payload_i[25];
  assign packet_o[28] = payload_i[24];
  assign packet_o[27] = payload_i[23];
  assign packet_o[26] = payload_i[22];
  assign packet_o[25] = payload_i[21];
  assign packet_o[24] = payload_i[20];
  assign packet_o[23] = payload_i[19];
  assign packet_o[22] = payload_i[18];
  assign packet_o[21] = payload_i[17];
  assign packet_o[20] = payload_i[16];
  assign packet_o[19] = payload_i[15];
  assign packet_o[18] = payload_i[14];
  assign packet_o[17] = payload_i[13];
  assign packet_o[16] = payload_i[12];
  assign packet_o[15] = payload_i[11];
  assign packet_o[14] = payload_i[10];
  assign packet_o[13] = payload_i[9];
  assign packet_o[12] = payload_i[8];
  assign packet_o[11] = payload_i[7];
  assign packet_o[10] = payload_i[6];
  assign packet_o[0] = payload_i[5];
  assign packet_o[9] = payload_i[5];
  assign packet_o[8] = payload_i[4];
  assign packet_o[7] = payload_i[3];
  assign packet_o[6] = payload_i[2];
  assign packet_o[5] = payload_i[1];
  assign packet_o[4] = payload_i[0];
  assign N6 = N4 & N5;
  assign N7 = payload_i[4] | N5;
  assign N9 = N4 | payload_i[3];
  assign N11 = payload_i[4] & payload_i[3];
  assign packet_o[3:2] = (N0)? { 1'b1, 1'b1 } :
                         (N1)? { 1'b1, 1'b1 } :
                         (N2)? { 1'b0, 1'b0 } :
                         (N3)? { 1'b0, 1'b0 } : 1'b0;
  assign N0 = N6;
  assign N1 = N8;
  assign N2 = N10;
  assign N3 = N11;
  assign N4 = ~payload_i[4];
  assign N5 = ~payload_i[3];
  assign N8 = ~N7;
  assign N10 = ~N9;

endmodule



module bsg_mux_width_p131_els_p4
(
  data_i,
  sel_i,
  data_o
);

  input [523:0] data_i;
  input [1:0] sel_i;
  output [130:0] data_o;
  wire [130:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[130] = (N2)? data_i[130] :
                       (N4)? data_i[261] :
                       (N3)? data_i[392] :
                       (N5)? data_i[523] : 1'b0;
  assign data_o[129] = (N2)? data_i[129] :
                       (N4)? data_i[260] :
                       (N3)? data_i[391] :
                       (N5)? data_i[522] : 1'b0;
  assign data_o[128] = (N2)? data_i[128] :
                       (N4)? data_i[259] :
                       (N3)? data_i[390] :
                       (N5)? data_i[521] : 1'b0;
  assign data_o[127] = (N2)? data_i[127] :
                       (N4)? data_i[258] :
                       (N3)? data_i[389] :
                       (N5)? data_i[520] : 1'b0;
  assign data_o[126] = (N2)? data_i[126] :
                       (N4)? data_i[257] :
                       (N3)? data_i[388] :
                       (N5)? data_i[519] : 1'b0;
  assign data_o[125] = (N2)? data_i[125] :
                       (N4)? data_i[256] :
                       (N3)? data_i[387] :
                       (N5)? data_i[518] : 1'b0;
  assign data_o[124] = (N2)? data_i[124] :
                       (N4)? data_i[255] :
                       (N3)? data_i[386] :
                       (N5)? data_i[517] : 1'b0;
  assign data_o[123] = (N2)? data_i[123] :
                       (N4)? data_i[254] :
                       (N3)? data_i[385] :
                       (N5)? data_i[516] : 1'b0;
  assign data_o[122] = (N2)? data_i[122] :
                       (N4)? data_i[253] :
                       (N3)? data_i[384] :
                       (N5)? data_i[515] : 1'b0;
  assign data_o[121] = (N2)? data_i[121] :
                       (N4)? data_i[252] :
                       (N3)? data_i[383] :
                       (N5)? data_i[514] : 1'b0;
  assign data_o[120] = (N2)? data_i[120] :
                       (N4)? data_i[251] :
                       (N3)? data_i[382] :
                       (N5)? data_i[513] : 1'b0;
  assign data_o[119] = (N2)? data_i[119] :
                       (N4)? data_i[250] :
                       (N3)? data_i[381] :
                       (N5)? data_i[512] : 1'b0;
  assign data_o[118] = (N2)? data_i[118] :
                       (N4)? data_i[249] :
                       (N3)? data_i[380] :
                       (N5)? data_i[511] : 1'b0;
  assign data_o[117] = (N2)? data_i[117] :
                       (N4)? data_i[248] :
                       (N3)? data_i[379] :
                       (N5)? data_i[510] : 1'b0;
  assign data_o[116] = (N2)? data_i[116] :
                       (N4)? data_i[247] :
                       (N3)? data_i[378] :
                       (N5)? data_i[509] : 1'b0;
  assign data_o[115] = (N2)? data_i[115] :
                       (N4)? data_i[246] :
                       (N3)? data_i[377] :
                       (N5)? data_i[508] : 1'b0;
  assign data_o[114] = (N2)? data_i[114] :
                       (N4)? data_i[245] :
                       (N3)? data_i[376] :
                       (N5)? data_i[507] : 1'b0;
  assign data_o[113] = (N2)? data_i[113] :
                       (N4)? data_i[244] :
                       (N3)? data_i[375] :
                       (N5)? data_i[506] : 1'b0;
  assign data_o[112] = (N2)? data_i[112] :
                       (N4)? data_i[243] :
                       (N3)? data_i[374] :
                       (N5)? data_i[505] : 1'b0;
  assign data_o[111] = (N2)? data_i[111] :
                       (N4)? data_i[242] :
                       (N3)? data_i[373] :
                       (N5)? data_i[504] : 1'b0;
  assign data_o[110] = (N2)? data_i[110] :
                       (N4)? data_i[241] :
                       (N3)? data_i[372] :
                       (N5)? data_i[503] : 1'b0;
  assign data_o[109] = (N2)? data_i[109] :
                       (N4)? data_i[240] :
                       (N3)? data_i[371] :
                       (N5)? data_i[502] : 1'b0;
  assign data_o[108] = (N2)? data_i[108] :
                       (N4)? data_i[239] :
                       (N3)? data_i[370] :
                       (N5)? data_i[501] : 1'b0;
  assign data_o[107] = (N2)? data_i[107] :
                       (N4)? data_i[238] :
                       (N3)? data_i[369] :
                       (N5)? data_i[500] : 1'b0;
  assign data_o[106] = (N2)? data_i[106] :
                       (N4)? data_i[237] :
                       (N3)? data_i[368] :
                       (N5)? data_i[499] : 1'b0;
  assign data_o[105] = (N2)? data_i[105] :
                       (N4)? data_i[236] :
                       (N3)? data_i[367] :
                       (N5)? data_i[498] : 1'b0;
  assign data_o[104] = (N2)? data_i[104] :
                       (N4)? data_i[235] :
                       (N3)? data_i[366] :
                       (N5)? data_i[497] : 1'b0;
  assign data_o[103] = (N2)? data_i[103] :
                       (N4)? data_i[234] :
                       (N3)? data_i[365] :
                       (N5)? data_i[496] : 1'b0;
  assign data_o[102] = (N2)? data_i[102] :
                       (N4)? data_i[233] :
                       (N3)? data_i[364] :
                       (N5)? data_i[495] : 1'b0;
  assign data_o[101] = (N2)? data_i[101] :
                       (N4)? data_i[232] :
                       (N3)? data_i[363] :
                       (N5)? data_i[494] : 1'b0;
  assign data_o[100] = (N2)? data_i[100] :
                       (N4)? data_i[231] :
                       (N3)? data_i[362] :
                       (N5)? data_i[493] : 1'b0;
  assign data_o[99] = (N2)? data_i[99] :
                      (N4)? data_i[230] :
                      (N3)? data_i[361] :
                      (N5)? data_i[492] : 1'b0;
  assign data_o[98] = (N2)? data_i[98] :
                      (N4)? data_i[229] :
                      (N3)? data_i[360] :
                      (N5)? data_i[491] : 1'b0;
  assign data_o[97] = (N2)? data_i[97] :
                      (N4)? data_i[228] :
                      (N3)? data_i[359] :
                      (N5)? data_i[490] : 1'b0;
  assign data_o[96] = (N2)? data_i[96] :
                      (N4)? data_i[227] :
                      (N3)? data_i[358] :
                      (N5)? data_i[489] : 1'b0;
  assign data_o[95] = (N2)? data_i[95] :
                      (N4)? data_i[226] :
                      (N3)? data_i[357] :
                      (N5)? data_i[488] : 1'b0;
  assign data_o[94] = (N2)? data_i[94] :
                      (N4)? data_i[225] :
                      (N3)? data_i[356] :
                      (N5)? data_i[487] : 1'b0;
  assign data_o[93] = (N2)? data_i[93] :
                      (N4)? data_i[224] :
                      (N3)? data_i[355] :
                      (N5)? data_i[486] : 1'b0;
  assign data_o[92] = (N2)? data_i[92] :
                      (N4)? data_i[223] :
                      (N3)? data_i[354] :
                      (N5)? data_i[485] : 1'b0;
  assign data_o[91] = (N2)? data_i[91] :
                      (N4)? data_i[222] :
                      (N3)? data_i[353] :
                      (N5)? data_i[484] : 1'b0;
  assign data_o[90] = (N2)? data_i[90] :
                      (N4)? data_i[221] :
                      (N3)? data_i[352] :
                      (N5)? data_i[483] : 1'b0;
  assign data_o[89] = (N2)? data_i[89] :
                      (N4)? data_i[220] :
                      (N3)? data_i[351] :
                      (N5)? data_i[482] : 1'b0;
  assign data_o[88] = (N2)? data_i[88] :
                      (N4)? data_i[219] :
                      (N3)? data_i[350] :
                      (N5)? data_i[481] : 1'b0;
  assign data_o[87] = (N2)? data_i[87] :
                      (N4)? data_i[218] :
                      (N3)? data_i[349] :
                      (N5)? data_i[480] : 1'b0;
  assign data_o[86] = (N2)? data_i[86] :
                      (N4)? data_i[217] :
                      (N3)? data_i[348] :
                      (N5)? data_i[479] : 1'b0;
  assign data_o[85] = (N2)? data_i[85] :
                      (N4)? data_i[216] :
                      (N3)? data_i[347] :
                      (N5)? data_i[478] : 1'b0;
  assign data_o[84] = (N2)? data_i[84] :
                      (N4)? data_i[215] :
                      (N3)? data_i[346] :
                      (N5)? data_i[477] : 1'b0;
  assign data_o[83] = (N2)? data_i[83] :
                      (N4)? data_i[214] :
                      (N3)? data_i[345] :
                      (N5)? data_i[476] : 1'b0;
  assign data_o[82] = (N2)? data_i[82] :
                      (N4)? data_i[213] :
                      (N3)? data_i[344] :
                      (N5)? data_i[475] : 1'b0;
  assign data_o[81] = (N2)? data_i[81] :
                      (N4)? data_i[212] :
                      (N3)? data_i[343] :
                      (N5)? data_i[474] : 1'b0;
  assign data_o[80] = (N2)? data_i[80] :
                      (N4)? data_i[211] :
                      (N3)? data_i[342] :
                      (N5)? data_i[473] : 1'b0;
  assign data_o[79] = (N2)? data_i[79] :
                      (N4)? data_i[210] :
                      (N3)? data_i[341] :
                      (N5)? data_i[472] : 1'b0;
  assign data_o[78] = (N2)? data_i[78] :
                      (N4)? data_i[209] :
                      (N3)? data_i[340] :
                      (N5)? data_i[471] : 1'b0;
  assign data_o[77] = (N2)? data_i[77] :
                      (N4)? data_i[208] :
                      (N3)? data_i[339] :
                      (N5)? data_i[470] : 1'b0;
  assign data_o[76] = (N2)? data_i[76] :
                      (N4)? data_i[207] :
                      (N3)? data_i[338] :
                      (N5)? data_i[469] : 1'b0;
  assign data_o[75] = (N2)? data_i[75] :
                      (N4)? data_i[206] :
                      (N3)? data_i[337] :
                      (N5)? data_i[468] : 1'b0;
  assign data_o[74] = (N2)? data_i[74] :
                      (N4)? data_i[205] :
                      (N3)? data_i[336] :
                      (N5)? data_i[467] : 1'b0;
  assign data_o[73] = (N2)? data_i[73] :
                      (N4)? data_i[204] :
                      (N3)? data_i[335] :
                      (N5)? data_i[466] : 1'b0;
  assign data_o[72] = (N2)? data_i[72] :
                      (N4)? data_i[203] :
                      (N3)? data_i[334] :
                      (N5)? data_i[465] : 1'b0;
  assign data_o[71] = (N2)? data_i[71] :
                      (N4)? data_i[202] :
                      (N3)? data_i[333] :
                      (N5)? data_i[464] : 1'b0;
  assign data_o[70] = (N2)? data_i[70] :
                      (N4)? data_i[201] :
                      (N3)? data_i[332] :
                      (N5)? data_i[463] : 1'b0;
  assign data_o[69] = (N2)? data_i[69] :
                      (N4)? data_i[200] :
                      (N3)? data_i[331] :
                      (N5)? data_i[462] : 1'b0;
  assign data_o[68] = (N2)? data_i[68] :
                      (N4)? data_i[199] :
                      (N3)? data_i[330] :
                      (N5)? data_i[461] : 1'b0;
  assign data_o[67] = (N2)? data_i[67] :
                      (N4)? data_i[198] :
                      (N3)? data_i[329] :
                      (N5)? data_i[460] : 1'b0;
  assign data_o[66] = (N2)? data_i[66] :
                      (N4)? data_i[197] :
                      (N3)? data_i[328] :
                      (N5)? data_i[459] : 1'b0;
  assign data_o[65] = (N2)? data_i[65] :
                      (N4)? data_i[196] :
                      (N3)? data_i[327] :
                      (N5)? data_i[458] : 1'b0;
  assign data_o[64] = (N2)? data_i[64] :
                      (N4)? data_i[195] :
                      (N3)? data_i[326] :
                      (N5)? data_i[457] : 1'b0;
  assign data_o[63] = (N2)? data_i[63] :
                      (N4)? data_i[194] :
                      (N3)? data_i[325] :
                      (N5)? data_i[456] : 1'b0;
  assign data_o[62] = (N2)? data_i[62] :
                      (N4)? data_i[193] :
                      (N3)? data_i[324] :
                      (N5)? data_i[455] : 1'b0;
  assign data_o[61] = (N2)? data_i[61] :
                      (N4)? data_i[192] :
                      (N3)? data_i[323] :
                      (N5)? data_i[454] : 1'b0;
  assign data_o[60] = (N2)? data_i[60] :
                      (N4)? data_i[191] :
                      (N3)? data_i[322] :
                      (N5)? data_i[453] : 1'b0;
  assign data_o[59] = (N2)? data_i[59] :
                      (N4)? data_i[190] :
                      (N3)? data_i[321] :
                      (N5)? data_i[452] : 1'b0;
  assign data_o[58] = (N2)? data_i[58] :
                      (N4)? data_i[189] :
                      (N3)? data_i[320] :
                      (N5)? data_i[451] : 1'b0;
  assign data_o[57] = (N2)? data_i[57] :
                      (N4)? data_i[188] :
                      (N3)? data_i[319] :
                      (N5)? data_i[450] : 1'b0;
  assign data_o[56] = (N2)? data_i[56] :
                      (N4)? data_i[187] :
                      (N3)? data_i[318] :
                      (N5)? data_i[449] : 1'b0;
  assign data_o[55] = (N2)? data_i[55] :
                      (N4)? data_i[186] :
                      (N3)? data_i[317] :
                      (N5)? data_i[448] : 1'b0;
  assign data_o[54] = (N2)? data_i[54] :
                      (N4)? data_i[185] :
                      (N3)? data_i[316] :
                      (N5)? data_i[447] : 1'b0;
  assign data_o[53] = (N2)? data_i[53] :
                      (N4)? data_i[184] :
                      (N3)? data_i[315] :
                      (N5)? data_i[446] : 1'b0;
  assign data_o[52] = (N2)? data_i[52] :
                      (N4)? data_i[183] :
                      (N3)? data_i[314] :
                      (N5)? data_i[445] : 1'b0;
  assign data_o[51] = (N2)? data_i[51] :
                      (N4)? data_i[182] :
                      (N3)? data_i[313] :
                      (N5)? data_i[444] : 1'b0;
  assign data_o[50] = (N2)? data_i[50] :
                      (N4)? data_i[181] :
                      (N3)? data_i[312] :
                      (N5)? data_i[443] : 1'b0;
  assign data_o[49] = (N2)? data_i[49] :
                      (N4)? data_i[180] :
                      (N3)? data_i[311] :
                      (N5)? data_i[442] : 1'b0;
  assign data_o[48] = (N2)? data_i[48] :
                      (N4)? data_i[179] :
                      (N3)? data_i[310] :
                      (N5)? data_i[441] : 1'b0;
  assign data_o[47] = (N2)? data_i[47] :
                      (N4)? data_i[178] :
                      (N3)? data_i[309] :
                      (N5)? data_i[440] : 1'b0;
  assign data_o[46] = (N2)? data_i[46] :
                      (N4)? data_i[177] :
                      (N3)? data_i[308] :
                      (N5)? data_i[439] : 1'b0;
  assign data_o[45] = (N2)? data_i[45] :
                      (N4)? data_i[176] :
                      (N3)? data_i[307] :
                      (N5)? data_i[438] : 1'b0;
  assign data_o[44] = (N2)? data_i[44] :
                      (N4)? data_i[175] :
                      (N3)? data_i[306] :
                      (N5)? data_i[437] : 1'b0;
  assign data_o[43] = (N2)? data_i[43] :
                      (N4)? data_i[174] :
                      (N3)? data_i[305] :
                      (N5)? data_i[436] : 1'b0;
  assign data_o[42] = (N2)? data_i[42] :
                      (N4)? data_i[173] :
                      (N3)? data_i[304] :
                      (N5)? data_i[435] : 1'b0;
  assign data_o[41] = (N2)? data_i[41] :
                      (N4)? data_i[172] :
                      (N3)? data_i[303] :
                      (N5)? data_i[434] : 1'b0;
  assign data_o[40] = (N2)? data_i[40] :
                      (N4)? data_i[171] :
                      (N3)? data_i[302] :
                      (N5)? data_i[433] : 1'b0;
  assign data_o[39] = (N2)? data_i[39] :
                      (N4)? data_i[170] :
                      (N3)? data_i[301] :
                      (N5)? data_i[432] : 1'b0;
  assign data_o[38] = (N2)? data_i[38] :
                      (N4)? data_i[169] :
                      (N3)? data_i[300] :
                      (N5)? data_i[431] : 1'b0;
  assign data_o[37] = (N2)? data_i[37] :
                      (N4)? data_i[168] :
                      (N3)? data_i[299] :
                      (N5)? data_i[430] : 1'b0;
  assign data_o[36] = (N2)? data_i[36] :
                      (N4)? data_i[167] :
                      (N3)? data_i[298] :
                      (N5)? data_i[429] : 1'b0;
  assign data_o[35] = (N2)? data_i[35] :
                      (N4)? data_i[166] :
                      (N3)? data_i[297] :
                      (N5)? data_i[428] : 1'b0;
  assign data_o[34] = (N2)? data_i[34] :
                      (N4)? data_i[165] :
                      (N3)? data_i[296] :
                      (N5)? data_i[427] : 1'b0;
  assign data_o[33] = (N2)? data_i[33] :
                      (N4)? data_i[164] :
                      (N3)? data_i[295] :
                      (N5)? data_i[426] : 1'b0;
  assign data_o[32] = (N2)? data_i[32] :
                      (N4)? data_i[163] :
                      (N3)? data_i[294] :
                      (N5)? data_i[425] : 1'b0;
  assign data_o[31] = (N2)? data_i[31] :
                      (N4)? data_i[162] :
                      (N3)? data_i[293] :
                      (N5)? data_i[424] : 1'b0;
  assign data_o[30] = (N2)? data_i[30] :
                      (N4)? data_i[161] :
                      (N3)? data_i[292] :
                      (N5)? data_i[423] : 1'b0;
  assign data_o[29] = (N2)? data_i[29] :
                      (N4)? data_i[160] :
                      (N3)? data_i[291] :
                      (N5)? data_i[422] : 1'b0;
  assign data_o[28] = (N2)? data_i[28] :
                      (N4)? data_i[159] :
                      (N3)? data_i[290] :
                      (N5)? data_i[421] : 1'b0;
  assign data_o[27] = (N2)? data_i[27] :
                      (N4)? data_i[158] :
                      (N3)? data_i[289] :
                      (N5)? data_i[420] : 1'b0;
  assign data_o[26] = (N2)? data_i[26] :
                      (N4)? data_i[157] :
                      (N3)? data_i[288] :
                      (N5)? data_i[419] : 1'b0;
  assign data_o[25] = (N2)? data_i[25] :
                      (N4)? data_i[156] :
                      (N3)? data_i[287] :
                      (N5)? data_i[418] : 1'b0;
  assign data_o[24] = (N2)? data_i[24] :
                      (N4)? data_i[155] :
                      (N3)? data_i[286] :
                      (N5)? data_i[417] : 1'b0;
  assign data_o[23] = (N2)? data_i[23] :
                      (N4)? data_i[154] :
                      (N3)? data_i[285] :
                      (N5)? data_i[416] : 1'b0;
  assign data_o[22] = (N2)? data_i[22] :
                      (N4)? data_i[153] :
                      (N3)? data_i[284] :
                      (N5)? data_i[415] : 1'b0;
  assign data_o[21] = (N2)? data_i[21] :
                      (N4)? data_i[152] :
                      (N3)? data_i[283] :
                      (N5)? data_i[414] : 1'b0;
  assign data_o[20] = (N2)? data_i[20] :
                      (N4)? data_i[151] :
                      (N3)? data_i[282] :
                      (N5)? data_i[413] : 1'b0;
  assign data_o[19] = (N2)? data_i[19] :
                      (N4)? data_i[150] :
                      (N3)? data_i[281] :
                      (N5)? data_i[412] : 1'b0;
  assign data_o[18] = (N2)? data_i[18] :
                      (N4)? data_i[149] :
                      (N3)? data_i[280] :
                      (N5)? data_i[411] : 1'b0;
  assign data_o[17] = (N2)? data_i[17] :
                      (N4)? data_i[148] :
                      (N3)? data_i[279] :
                      (N5)? data_i[410] : 1'b0;
  assign data_o[16] = (N2)? data_i[16] :
                      (N4)? data_i[147] :
                      (N3)? data_i[278] :
                      (N5)? data_i[409] : 1'b0;
  assign data_o[15] = (N2)? data_i[15] :
                      (N4)? data_i[146] :
                      (N3)? data_i[277] :
                      (N5)? data_i[408] : 1'b0;
  assign data_o[14] = (N2)? data_i[14] :
                      (N4)? data_i[145] :
                      (N3)? data_i[276] :
                      (N5)? data_i[407] : 1'b0;
  assign data_o[13] = (N2)? data_i[13] :
                      (N4)? data_i[144] :
                      (N3)? data_i[275] :
                      (N5)? data_i[406] : 1'b0;
  assign data_o[12] = (N2)? data_i[12] :
                      (N4)? data_i[143] :
                      (N3)? data_i[274] :
                      (N5)? data_i[405] : 1'b0;
  assign data_o[11] = (N2)? data_i[11] :
                      (N4)? data_i[142] :
                      (N3)? data_i[273] :
                      (N5)? data_i[404] : 1'b0;
  assign data_o[10] = (N2)? data_i[10] :
                      (N4)? data_i[141] :
                      (N3)? data_i[272] :
                      (N5)? data_i[403] : 1'b0;
  assign data_o[9] = (N2)? data_i[9] :
                     (N4)? data_i[140] :
                     (N3)? data_i[271] :
                     (N5)? data_i[402] : 1'b0;
  assign data_o[8] = (N2)? data_i[8] :
                     (N4)? data_i[139] :
                     (N3)? data_i[270] :
                     (N5)? data_i[401] : 1'b0;
  assign data_o[7] = (N2)? data_i[7] :
                     (N4)? data_i[138] :
                     (N3)? data_i[269] :
                     (N5)? data_i[400] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] :
                     (N4)? data_i[137] :
                     (N3)? data_i[268] :
                     (N5)? data_i[399] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] :
                     (N4)? data_i[136] :
                     (N3)? data_i[267] :
                     (N5)? data_i[398] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] :
                     (N4)? data_i[135] :
                     (N3)? data_i[266] :
                     (N5)? data_i[397] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] :
                     (N4)? data_i[134] :
                     (N3)? data_i[265] :
                     (N5)? data_i[396] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] :
                     (N4)? data_i[133] :
                     (N3)? data_i[264] :
                     (N5)? data_i[395] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] :
                     (N4)? data_i[132] :
                     (N3)? data_i[263] :
                     (N5)? data_i[394] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] :
                     (N4)? data_i[131] :
                     (N3)? data_i[262] :
                     (N5)? data_i[393] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_wormhole_router_adapter_in_max_num_flit_p4_max_payload_width_p518_x_cord_width_p1_y_cord_width_p1
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  ready_o,
  data_o,
  v_o,
  ready_i
);

  input [521:0] data_i;
  output [130:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input ready_i;
  output ready_o;
  output v_o;
  wire [130:0] data_o;
  wire ready_o,v_o,N0,N1,N2,N3,state_n,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24,N25;
  wire [1:0] count_n;
  reg [1:0] count_r;
  reg state_r;

  bsg_mux_width_p131_els_p4
  mux
  (
    .data_i({ 1'b0, 1'b0, data_i }),
    .sel_i(count_r),
    .data_o(data_o)
  );

  assign N10 = count_r == data_i[3:2];
  assign N12 = count_r == data_i[3:2];
  assign { N9, N8 } = count_r + 1'b1;
  assign N14 = ~N13;
  assign count_n = (N0)? { 1'b0, 1'b0 } :
                   (N1)? { N9, N8 } : 1'b0;
  assign N0 = N4;
  assign N1 = v_o;
  assign state_n = (N0)? 1'b1 :
                   (N1)? N14 : 1'b0;
  assign ready_o = (N0)? 1'b0 :
                   (N1)? N11 : 1'b0;
  assign N16 = (N2)? 1'b0 :
               (N3)? state_n : 1'b0;
  assign N2 = reset_i;
  assign N3 = N15;
  assign { N18, N17 } = (N2)? { 1'b0, 1'b0 } :
                        (N3)? count_n : 1'b0;
  assign N4 = ~state_r;
  assign v_o = state_r;
  assign N5 = ~v_i;
  assign N6 = v_o;
  assign N7 = ~ready_i;
  assign N11 = ready_i & N10;
  assign N13 = ready_i & N12;
  assign N15 = ~reset_i;
  assign N19 = N4 & N15;
  assign N20 = N5 & N19;
  assign N21 = v_o & N15;
  assign N22 = N7 & N21;
  assign N23 = N20 | N22;
  assign N24 = ~N23;
  assign N25 = ~N20;

  always @(posedge clk_i) begin
    if(N24) begin
      { count_r[1:0] } <= { N18, N17 };
    end
    if(N25) begin
      state_r <= N16;
    end
  end


endmodule



module bsg_wormhole_router_adapter_out_max_num_flit_p4_max_payload_width_p518_x_cord_width_p1_y_cord_width_p1
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  ready_o,
  data_o,
  v_o,
  ready_i
);

  input [130:0] data_i;
  output [521:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input ready_i;
  output ready_o;
  output v_o;
  wire ready_o,v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,we,clear,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,
  N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,
  N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,
  N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,
  N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,
  N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,
  N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,
  N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,
  N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211;
  wire [1:0] state_n,count_n;
  reg [521:0] data_o;
  reg [1:0] state_r,count_r;
  assign N16 = N14 & N15;
  assign N17 = state_r[1] | N15;
  assign N19 = N14 | state_r[0];
  assign N21 = state_r[1] & state_r[0];
  assign N29 = data_o[3:2] == count_r;
  assign N210 = data_i[2] | data_i[3];
  assign N211 = ~N210;
  assign { N25, N24 } = count_r + 1'b1;
  assign { N28, N27 } = count_r + 1'b1;
  assign N38 = count_r[0] & count_r[1];
  assign N37 = N0 & count_r[1];
  assign N0 = ~count_r[0];
  assign N36 = count_r[0] & N1;
  assign N1 = ~count_r[1];
  assign N35 = N2 & N3;
  assign N2 = ~count_r[0];
  assign N3 = ~count_r[1];
  assign N30 = ~N29;
  assign ready_o = (N4)? 1'b1 :
                   (N5)? 1'b1 :
                   (N6)? 1'b0 :
                   (N7)? 1'b0 : 1'b0;
  assign N4 = N16;
  assign N5 = N18;
  assign N6 = N20;
  assign N7 = N21;
  assign state_n = (N4)? { N211, N210 } :
                   (N5)? { N29, N30 } :
                   (N6)? { 1'b0, 1'b0 } :
                   (N7)? { 1'b0, 1'b0 } : 1'b0;
  assign we = (N4)? v_i :
              (N5)? v_i :
              (N6)? ready_i :
              (N7)? 1'b0 : 1'b0;
  assign count_n = (N4)? { N25, N24 } :
                   (N5)? { N28, N27 } :
                   (N6)? { 1'b0, 1'b0 } : 1'b0;
  assign v_o = (N4)? 1'b0 :
               (N5)? 1'b0 :
               (N6)? 1'b1 :
               (N7)? 1'b0 : 1'b0;
  assign clear = (N4)? 1'b0 :
                 (N5)? 1'b0 :
                 (N6)? ready_i :
                 (N7)? 1'b0 : 1'b0;
  assign { N177, N176, N175, N174, N173, N172, N41, N39 } = (N8)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } :
                                                            (N9)? { N38, N38, N37, N37, N36, N36, N35, N35 } : 1'b0;
  assign N8 = clear;
  assign N9 = N34;
  assign { N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N40 } = (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (N9)? data_i : 1'b0;
  assign { N185, N184, N183, N182, N181, N180, N179, N178 } = (N10)? { N177, N176, N175, N174, N173, N172, N41, N39 } :
                                                              (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = we;
  assign N11 = N33;
  assign { N187, N186 } = (N12)? { 1'b0, 1'b0 } :
                          (N13)? state_n : 1'b0;
  assign N12 = reset_i;
  assign N13 = N32;
  assign { N189, N188 } = (N12)? { 1'b0, 1'b0 } :
                          (N13)? count_n : 1'b0;
  assign { N197, N196, N195, N194, N193, N192, N191, N190 } = (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                              (N13)? { N185, N184, N183, N182, N181, N180, N179, N178 } : 1'b0;
  assign N14 = ~state_r[1];
  assign N15 = ~state_r[0];
  assign N18 = ~N17;
  assign N20 = ~N19;
  assign N22 = N16;
  assign N23 = ~v_i;
  assign N26 = N18;
  assign N31 = ~ready_i;
  assign N32 = ~reset_i;
  assign N33 = ~we;
  assign N34 = ~clear;
  assign N198 = N16 & N32;
  assign N199 = N23 & N198;
  assign N200 = N18 & N32;
  assign N201 = N23 & N200;
  assign N202 = N199 | N201;
  assign N203 = N20 & N32;
  assign N204 = N31 & N203;
  assign N205 = N202 | N204;
  assign N206 = ~N205;
  assign N207 = N21 & N32;
  assign N208 = N205 | N207;
  assign N209 = ~N208;

  always @(posedge clk_i) begin
    if(N196) begin
      { data_o[521:423], data_o[393:393] } <= { N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N40 };
    end
    if(N197) begin
      { data_o[422:394] } <= { N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42 };
    end
    if(N194) begin
      { data_o[392:294], data_o[262:262] } <= { N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N40 };
    end
    if(N195) begin
      { data_o[293:263] } <= { N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42 };
    end
    if(N192) begin
      { data_o[261:163], data_o[131:131] } <= { N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N40 };
    end
    if(N193) begin
      { data_o[162:132] } <= { N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42 };
    end
    if(N190) begin
      { data_o[130:32], data_o[0:0] } <= { N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N40 };
    end
    if(N191) begin
      { data_o[31:1] } <= { N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42 };
    end
    if(N206) begin
      { state_r[1:0] } <= { N187, N186 };
    end
    if(N209) begin
      { count_r[1:0] } <= { N189, N188 };
    end
  end


endmodule



module bp_me_network_channel_data_cmd_num_lce_p2_num_cce_p1_lce_assoc_p8_block_size_in_bits_p512_max_num_flit_p4
(
  clk_i,
  reset_i,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i,
  cce_lce_data_cmd_i,
  cce_lce_data_cmd_v_i,
  cce_lce_data_cmd_ready_o,
  lce_lce_data_cmd_i,
  lce_lce_data_cmd_v_i,
  lce_lce_data_cmd_ready_o
);

  output [1035:0] lce_data_cmd_o;
  output [1:0] lce_data_cmd_v_o;
  input [1:0] lce_data_cmd_ready_i;
  input [517:0] cce_lce_data_cmd_i;
  input [0:0] cce_lce_data_cmd_v_i;
  output [0:0] cce_lce_data_cmd_ready_o;
  input [1035:0] lce_lce_data_cmd_i;
  input [1:0] lce_lce_data_cmd_v_i;
  output [1:0] lce_lce_data_cmd_ready_o;
  input clk_i;
  input reset_i;
  wire [1035:0] lce_data_cmd_o;
  wire [1:0] lce_data_cmd_v_o,lce_lce_data_cmd_ready_o;
  wire [0:0] cce_lce_data_cmd_ready_o;
  wire valid_li_1__4_,valid_li_1__3_,valid_li_1__2_,valid_li_1__0_,valid_li_0__4_,
  valid_li_0__3_,valid_li_0__1_,valid_li_0__0_,data_li_1__0__130_,data_li_1__0__129_,
  data_li_1__0__128_,data_li_1__0__127_,data_li_1__0__126_,data_li_1__0__125_,
  data_li_1__0__124_,data_li_1__0__123_,data_li_1__0__122_,data_li_1__0__121_,
  data_li_1__0__120_,data_li_1__0__119_,data_li_1__0__118_,data_li_1__0__117_,
  data_li_1__0__116_,data_li_1__0__115_,data_li_1__0__114_,data_li_1__0__113_,
  data_li_1__0__112_,data_li_1__0__111_,data_li_1__0__110_,data_li_1__0__109_,data_li_1__0__108_,
  data_li_1__0__107_,data_li_1__0__106_,data_li_1__0__105_,data_li_1__0__104_,
  data_li_1__0__103_,data_li_1__0__102_,data_li_1__0__101_,data_li_1__0__100_,
  data_li_1__0__99_,data_li_1__0__98_,data_li_1__0__97_,data_li_1__0__96_,data_li_1__0__95_,
  data_li_1__0__94_,data_li_1__0__93_,data_li_1__0__92_,data_li_1__0__91_,
  data_li_1__0__90_,data_li_1__0__89_,data_li_1__0__88_,data_li_1__0__87_,
  data_li_1__0__86_,data_li_1__0__85_,data_li_1__0__84_,data_li_1__0__83_,data_li_1__0__82_,
  data_li_1__0__81_,data_li_1__0__80_,data_li_1__0__79_,data_li_1__0__78_,
  data_li_1__0__77_,data_li_1__0__76_,data_li_1__0__75_,data_li_1__0__74_,data_li_1__0__73_,
  data_li_1__0__72_,data_li_1__0__71_,data_li_1__0__70_,data_li_1__0__69_,
  data_li_1__0__68_,data_li_1__0__67_,data_li_1__0__66_,data_li_1__0__65_,data_li_1__0__64_,
  data_li_1__0__63_,data_li_1__0__62_,data_li_1__0__61_,data_li_1__0__60_,
  data_li_1__0__59_,data_li_1__0__58_,data_li_1__0__57_,data_li_1__0__56_,data_li_1__0__55_,
  data_li_1__0__54_,data_li_1__0__53_,data_li_1__0__52_,data_li_1__0__51_,
  data_li_1__0__50_,data_li_1__0__49_,data_li_1__0__48_,data_li_1__0__47_,
  data_li_1__0__46_,data_li_1__0__45_,data_li_1__0__44_,data_li_1__0__43_,data_li_1__0__42_,
  data_li_1__0__41_,data_li_1__0__40_,data_li_1__0__39_,data_li_1__0__38_,
  data_li_1__0__37_,data_li_1__0__36_,data_li_1__0__35_,data_li_1__0__34_,data_li_1__0__33_,
  data_li_1__0__32_,data_li_1__0__31_,data_li_1__0__30_,data_li_1__0__29_,
  data_li_1__0__28_,data_li_1__0__27_,data_li_1__0__26_,data_li_1__0__25_,data_li_1__0__24_,
  data_li_1__0__23_,data_li_1__0__22_,data_li_1__0__21_,data_li_1__0__20_,
  data_li_1__0__19_,data_li_1__0__18_,data_li_1__0__17_,data_li_1__0__16_,data_li_1__0__15_,
  data_li_1__0__14_,data_li_1__0__13_,data_li_1__0__12_,data_li_1__0__11_,
  data_li_1__0__10_,data_li_1__0__9_,data_li_1__0__8_,data_li_1__0__7_,data_li_1__0__6_,
  data_li_1__0__5_,data_li_1__0__4_,data_li_1__0__3_,data_li_1__0__2_,
  data_li_1__0__1_,data_li_1__0__0_,data_li_0__4__130_,data_li_0__4__129_,data_li_0__4__128_,
  data_li_0__4__127_,data_li_0__4__126_,data_li_0__4__125_,data_li_0__4__124_,
  data_li_0__4__123_,data_li_0__4__122_,data_li_0__4__121_,data_li_0__4__120_,
  data_li_0__4__119_,data_li_0__4__118_,data_li_0__4__117_,data_li_0__4__116_,
  data_li_0__4__115_,data_li_0__4__114_,data_li_0__4__113_,data_li_0__4__112_,data_li_0__4__111_,
  data_li_0__4__110_,data_li_0__4__109_,data_li_0__4__108_,data_li_0__4__107_,
  data_li_0__4__106_,data_li_0__4__105_,data_li_0__4__104_,data_li_0__4__103_,
  data_li_0__4__102_,data_li_0__4__101_,data_li_0__4__100_,data_li_0__4__99_,
  data_li_0__4__98_,data_li_0__4__97_,data_li_0__4__96_,data_li_0__4__95_,data_li_0__4__94_,
  data_li_0__4__93_,data_li_0__4__92_,data_li_0__4__91_,data_li_0__4__90_,
  data_li_0__4__89_,data_li_0__4__88_,data_li_0__4__87_,data_li_0__4__86_,data_li_0__4__85_,
  data_li_0__4__84_,data_li_0__4__83_,data_li_0__4__82_,data_li_0__4__81_,
  data_li_0__4__80_,data_li_0__4__79_,data_li_0__4__78_,data_li_0__4__77_,data_li_0__4__76_,
  data_li_0__4__75_,data_li_0__4__74_,data_li_0__4__73_,data_li_0__4__72_,
  data_li_0__4__71_,data_li_0__4__70_,data_li_0__4__69_,data_li_0__4__68_,
  data_li_0__4__67_,data_li_0__4__66_,data_li_0__4__65_,data_li_0__4__64_,data_li_0__4__63_,
  data_li_0__4__62_,data_li_0__4__61_,data_li_0__4__60_,data_li_0__4__59_,
  data_li_0__4__58_,data_li_0__4__57_,data_li_0__4__56_,data_li_0__4__55_,data_li_0__4__54_,
  data_li_0__4__53_,data_li_0__4__52_,data_li_0__4__51_,data_li_0__4__50_,
  data_li_0__4__49_,data_li_0__4__48_,data_li_0__4__47_,data_li_0__4__46_,data_li_0__4__45_,
  data_li_0__4__44_,data_li_0__4__43_,data_li_0__4__42_,data_li_0__4__41_,
  data_li_0__4__40_,data_li_0__4__39_,data_li_0__4__38_,data_li_0__4__37_,data_li_0__4__36_,
  data_li_0__4__35_,data_li_0__4__34_,data_li_0__4__33_,data_li_0__4__32_,
  data_li_0__4__31_,data_li_0__4__30_,data_li_0__4__29_,data_li_0__4__28_,
  data_li_0__4__27_,data_li_0__4__26_,data_li_0__4__25_,data_li_0__4__24_,data_li_0__4__23_,
  data_li_0__4__22_,data_li_0__4__21_,data_li_0__4__20_,data_li_0__4__19_,
  data_li_0__4__18_,data_li_0__4__17_,data_li_0__4__16_,data_li_0__4__15_,data_li_0__4__14_,
  data_li_0__4__13_,data_li_0__4__12_,data_li_0__4__11_,data_li_0__4__10_,
  data_li_0__4__9_,data_li_0__4__8_,data_li_0__4__7_,data_li_0__4__6_,data_li_0__4__5_,
  data_li_0__4__4_,data_li_0__4__3_,data_li_0__4__2_,data_li_0__4__1_,data_li_0__4__0_,
  data_li_0__3__130_,data_li_0__3__129_,data_li_0__3__128_,data_li_0__3__127_,
  data_li_0__3__126_,data_li_0__3__125_,data_li_0__3__124_,data_li_0__3__123_,
  data_li_0__3__122_,data_li_0__3__121_,data_li_0__3__120_,data_li_0__3__119_,
  data_li_0__3__118_,data_li_0__3__117_,data_li_0__3__116_,data_li_0__3__115_,
  data_li_0__3__114_,data_li_0__3__113_,data_li_0__3__112_,data_li_0__3__111_,data_li_0__3__110_,
  data_li_0__3__109_,data_li_0__3__108_,data_li_0__3__107_,data_li_0__3__106_,
  data_li_0__3__105_,data_li_0__3__104_,data_li_0__3__103_,data_li_0__3__102_,
  data_li_0__3__101_,data_li_0__3__100_,data_li_0__3__99_,data_li_0__3__98_,
  data_li_0__3__97_,data_li_0__3__96_,data_li_0__3__95_,data_li_0__3__94_,data_li_0__3__93_,
  data_li_0__3__92_,data_li_0__3__91_,data_li_0__3__90_,data_li_0__3__89_,
  data_li_0__3__88_,data_li_0__3__87_,data_li_0__3__86_,data_li_0__3__85_,data_li_0__3__84_,
  data_li_0__3__83_,data_li_0__3__82_,data_li_0__3__81_,data_li_0__3__80_,
  data_li_0__3__79_,data_li_0__3__78_,data_li_0__3__77_,data_li_0__3__76_,data_li_0__3__75_,
  data_li_0__3__74_,data_li_0__3__73_,data_li_0__3__72_,data_li_0__3__71_,
  data_li_0__3__70_,data_li_0__3__69_,data_li_0__3__68_,data_li_0__3__67_,data_li_0__3__66_,
  data_li_0__3__65_,data_li_0__3__64_,data_li_0__3__63_,data_li_0__3__62_,
  data_li_0__3__61_,data_li_0__3__60_,data_li_0__3__59_,data_li_0__3__58_,
  data_li_0__3__57_,data_li_0__3__56_,data_li_0__3__55_,data_li_0__3__54_,data_li_0__3__53_,
  data_li_0__3__52_,data_li_0__3__51_,data_li_0__3__50_,data_li_0__3__49_,
  data_li_0__3__48_,data_li_0__3__47_,data_li_0__3__46_,data_li_0__3__45_,data_li_0__3__44_,
  data_li_0__3__43_,data_li_0__3__42_,data_li_0__3__41_,data_li_0__3__40_,
  data_li_0__3__39_,data_li_0__3__38_,data_li_0__3__37_,data_li_0__3__36_,data_li_0__3__35_,
  data_li_0__3__34_,data_li_0__3__33_,data_li_0__3__32_,data_li_0__3__31_,
  data_li_0__3__30_,data_li_0__3__29_,data_li_0__3__28_,data_li_0__3__27_,data_li_0__3__26_,
  data_li_0__3__25_,data_li_0__3__24_,data_li_0__3__23_,data_li_0__3__22_,
  data_li_0__3__21_,data_li_0__3__20_,data_li_0__3__19_,data_li_0__3__18_,
  data_li_0__3__17_,data_li_0__3__16_,data_li_0__3__15_,data_li_0__3__14_,data_li_0__3__13_,
  data_li_0__3__12_,data_li_0__3__11_,data_li_0__3__10_,data_li_0__3__9_,
  data_li_0__3__8_,data_li_0__3__7_,data_li_0__3__6_,data_li_0__3__5_,data_li_0__3__4_,
  data_li_0__3__3_,data_li_0__3__2_,data_li_0__3__1_,data_li_0__3__0_,data_li_0__1__130_,
  data_li_0__1__129_,data_li_0__1__128_,data_li_0__1__127_,data_li_0__1__126_,
  data_li_0__1__125_,data_li_0__1__124_,data_li_0__1__123_,data_li_0__1__122_,
  data_li_0__1__121_,data_li_0__1__120_,data_li_0__1__119_,data_li_0__1__118_,
  data_li_0__1__117_,data_li_0__1__116_,data_li_0__1__115_,data_li_0__1__114_,data_li_0__1__113_,
  data_li_0__1__112_,data_li_0__1__111_,data_li_0__1__110_,data_li_0__1__109_,
  data_li_0__1__108_,data_li_0__1__107_,data_li_0__1__106_,data_li_0__1__105_,
  data_li_0__1__104_,data_li_0__1__103_,data_li_0__1__102_,data_li_0__1__101_,
  data_li_0__1__100_,data_li_0__1__99_,data_li_0__1__98_,data_li_0__1__97_,data_li_0__1__96_,
  data_li_0__1__95_,data_li_0__1__94_,data_li_0__1__93_,data_li_0__1__92_,
  data_li_0__1__91_,data_li_0__1__90_,data_li_0__1__89_,data_li_0__1__88_,data_li_0__1__87_,
  data_li_0__1__86_,data_li_0__1__85_,data_li_0__1__84_,data_li_0__1__83_,
  data_li_0__1__82_,data_li_0__1__81_,data_li_0__1__80_,data_li_0__1__79_,
  data_li_0__1__78_,data_li_0__1__77_,data_li_0__1__76_,data_li_0__1__75_,data_li_0__1__74_,
  data_li_0__1__73_,data_li_0__1__72_,data_li_0__1__71_,data_li_0__1__70_,
  data_li_0__1__69_,data_li_0__1__68_,data_li_0__1__67_,data_li_0__1__66_,data_li_0__1__65_,
  data_li_0__1__64_,data_li_0__1__63_,data_li_0__1__62_,data_li_0__1__61_,
  data_li_0__1__60_,data_li_0__1__59_,data_li_0__1__58_,data_li_0__1__57_,data_li_0__1__56_,
  data_li_0__1__55_,data_li_0__1__54_,data_li_0__1__53_,data_li_0__1__52_,
  data_li_0__1__51_,data_li_0__1__50_,data_li_0__1__49_,data_li_0__1__48_,data_li_0__1__47_,
  data_li_0__1__46_,data_li_0__1__45_,data_li_0__1__44_,data_li_0__1__43_,
  data_li_0__1__42_,data_li_0__1__41_,data_li_0__1__40_,data_li_0__1__39_,
  data_li_0__1__38_,data_li_0__1__37_,data_li_0__1__36_,data_li_0__1__35_,data_li_0__1__34_,
  data_li_0__1__33_,data_li_0__1__32_,data_li_0__1__31_,data_li_0__1__30_,
  data_li_0__1__29_,data_li_0__1__28_,data_li_0__1__27_,data_li_0__1__26_,data_li_0__1__25_,
  data_li_0__1__24_,data_li_0__1__23_,data_li_0__1__22_,data_li_0__1__21_,
  data_li_0__1__20_,data_li_0__1__19_,data_li_0__1__18_,data_li_0__1__17_,data_li_0__1__16_,
  data_li_0__1__15_,data_li_0__1__14_,data_li_0__1__13_,data_li_0__1__12_,
  data_li_0__1__11_,data_li_0__1__10_,data_li_0__1__9_,data_li_0__1__8_,data_li_0__1__7_,
  data_li_0__1__6_,data_li_0__1__5_,data_li_0__1__4_,data_li_0__1__3_,
  data_li_0__1__2_,data_li_0__1__1_,data_li_0__1__0_,data_li_0__0__130_,data_li_0__0__129_,
  data_li_0__0__128_,data_li_0__0__127_,data_li_0__0__126_,data_li_0__0__125_,
  data_li_0__0__124_,data_li_0__0__123_,data_li_0__0__122_,data_li_0__0__121_,
  data_li_0__0__120_,data_li_0__0__119_,data_li_0__0__118_,data_li_0__0__117_,
  data_li_0__0__116_,data_li_0__0__115_,data_li_0__0__114_,data_li_0__0__113_,data_li_0__0__112_,
  data_li_0__0__111_,data_li_0__0__110_,data_li_0__0__109_,data_li_0__0__108_,
  data_li_0__0__107_,data_li_0__0__106_,data_li_0__0__105_,data_li_0__0__104_,
  data_li_0__0__103_,data_li_0__0__102_,data_li_0__0__101_,data_li_0__0__100_,
  data_li_0__0__99_,data_li_0__0__98_,data_li_0__0__97_,data_li_0__0__96_,data_li_0__0__95_,
  data_li_0__0__94_,data_li_0__0__93_,data_li_0__0__92_,data_li_0__0__91_,
  data_li_0__0__90_,data_li_0__0__89_,data_li_0__0__88_,data_li_0__0__87_,data_li_0__0__86_,
  data_li_0__0__85_,data_li_0__0__84_,data_li_0__0__83_,data_li_0__0__82_,
  data_li_0__0__81_,data_li_0__0__80_,data_li_0__0__79_,data_li_0__0__78_,data_li_0__0__77_,
  data_li_0__0__76_,data_li_0__0__75_,data_li_0__0__74_,data_li_0__0__73_,
  data_li_0__0__72_,data_li_0__0__71_,data_li_0__0__70_,data_li_0__0__69_,
  data_li_0__0__68_,data_li_0__0__67_,data_li_0__0__66_,data_li_0__0__65_,data_li_0__0__64_,
  data_li_0__0__63_,data_li_0__0__62_,data_li_0__0__61_,data_li_0__0__60_,
  data_li_0__0__59_,data_li_0__0__58_,data_li_0__0__57_,data_li_0__0__56_,data_li_0__0__55_,
  data_li_0__0__54_,data_li_0__0__53_,data_li_0__0__52_,data_li_0__0__51_,
  data_li_0__0__50_,data_li_0__0__49_,data_li_0__0__48_,data_li_0__0__47_,data_li_0__0__46_,
  data_li_0__0__45_,data_li_0__0__44_,data_li_0__0__43_,data_li_0__0__42_,
  data_li_0__0__41_,data_li_0__0__40_,data_li_0__0__39_,data_li_0__0__38_,data_li_0__0__37_,
  data_li_0__0__36_,data_li_0__0__35_,data_li_0__0__34_,data_li_0__0__33_,
  data_li_0__0__32_,data_li_0__0__31_,data_li_0__0__30_,data_li_0__0__29_,
  data_li_0__0__28_,data_li_0__0__27_,data_li_0__0__26_,data_li_0__0__25_,data_li_0__0__24_,
  data_li_0__0__23_,data_li_0__0__22_,data_li_0__0__21_,data_li_0__0__20_,
  data_li_0__0__19_,data_li_0__0__18_,data_li_0__0__17_,data_li_0__0__16_,data_li_0__0__15_,
  data_li_0__0__14_,data_li_0__0__13_,data_li_0__0__12_,data_li_0__0__11_,
  data_li_0__0__10_,data_li_0__0__9_,data_li_0__0__8_,data_li_0__0__7_,data_li_0__0__6_,
  data_li_0__0__5_,data_li_0__0__4_,data_li_0__0__3_,data_li_0__0__2_,data_li_0__0__1_,
  data_li_0__0__0_,ready_li_1__4_,ready_li_1__3_,ready_li_1__2_,ready_li_1__0_,
  ready_li_0__4_,ready_li_0__3_,ready_li_0__1_,ready_li_0__0_,data_li_1__4__130_,
  data_li_1__4__129_,data_li_1__4__128_,data_li_1__4__127_,data_li_1__4__126_,
  data_li_1__4__125_,data_li_1__4__124_,data_li_1__4__123_,data_li_1__4__122_,
  data_li_1__4__121_,data_li_1__4__120_,data_li_1__4__119_,data_li_1__4__118_,
  data_li_1__4__117_,data_li_1__4__116_,data_li_1__4__115_,data_li_1__4__114_,data_li_1__4__113_,
  data_li_1__4__112_,data_li_1__4__111_,data_li_1__4__110_,data_li_1__4__109_,
  data_li_1__4__108_,data_li_1__4__107_,data_li_1__4__106_,data_li_1__4__105_,
  data_li_1__4__104_,data_li_1__4__103_,data_li_1__4__102_,data_li_1__4__101_,
  data_li_1__4__100_,data_li_1__4__99_,data_li_1__4__98_,data_li_1__4__97_,data_li_1__4__96_,
  data_li_1__4__95_,data_li_1__4__94_,data_li_1__4__93_,data_li_1__4__92_,
  data_li_1__4__91_,data_li_1__4__90_,data_li_1__4__89_,data_li_1__4__88_,data_li_1__4__87_,
  data_li_1__4__86_,data_li_1__4__85_,data_li_1__4__84_,data_li_1__4__83_,
  data_li_1__4__82_,data_li_1__4__81_,data_li_1__4__80_,data_li_1__4__79_,data_li_1__4__78_,
  data_li_1__4__77_,data_li_1__4__76_,data_li_1__4__75_,data_li_1__4__74_,
  data_li_1__4__73_,data_li_1__4__72_,data_li_1__4__71_,data_li_1__4__70_,
  data_li_1__4__69_,data_li_1__4__68_,data_li_1__4__67_,data_li_1__4__66_,data_li_1__4__65_,
  data_li_1__4__64_,data_li_1__4__63_,data_li_1__4__62_,data_li_1__4__61_,
  data_li_1__4__60_,data_li_1__4__59_,data_li_1__4__58_,data_li_1__4__57_,data_li_1__4__56_,
  data_li_1__4__55_,data_li_1__4__54_,data_li_1__4__53_,data_li_1__4__52_,
  data_li_1__4__51_,data_li_1__4__50_,data_li_1__4__49_,data_li_1__4__48_,data_li_1__4__47_,
  data_li_1__4__46_,data_li_1__4__45_,data_li_1__4__44_,data_li_1__4__43_,
  data_li_1__4__42_,data_li_1__4__41_,data_li_1__4__40_,data_li_1__4__39_,data_li_1__4__38_,
  data_li_1__4__37_,data_li_1__4__36_,data_li_1__4__35_,data_li_1__4__34_,
  data_li_1__4__33_,data_li_1__4__32_,data_li_1__4__31_,data_li_1__4__30_,
  data_li_1__4__29_,data_li_1__4__28_,data_li_1__4__27_,data_li_1__4__26_,data_li_1__4__25_,
  data_li_1__4__24_,data_li_1__4__23_,data_li_1__4__22_,data_li_1__4__21_,
  data_li_1__4__20_,data_li_1__4__19_,data_li_1__4__18_,data_li_1__4__17_,data_li_1__4__16_,
  data_li_1__4__15_,data_li_1__4__14_,data_li_1__4__13_,data_li_1__4__12_,
  data_li_1__4__11_,data_li_1__4__10_,data_li_1__4__9_,data_li_1__4__8_,data_li_1__4__7_,
  data_li_1__4__6_,data_li_1__4__5_,data_li_1__4__4_,data_li_1__4__3_,data_li_1__4__2_,
  data_li_1__4__1_,data_li_1__4__0_,data_li_1__3__130_,data_li_1__3__129_,
  data_li_1__3__128_,data_li_1__3__127_,data_li_1__3__126_,data_li_1__3__125_,
  data_li_1__3__124_,data_li_1__3__123_,data_li_1__3__122_,data_li_1__3__121_,
  data_li_1__3__120_,data_li_1__3__119_,data_li_1__3__118_,data_li_1__3__117_,data_li_1__3__116_,
  data_li_1__3__115_,data_li_1__3__114_,data_li_1__3__113_,data_li_1__3__112_,
  data_li_1__3__111_,data_li_1__3__110_,data_li_1__3__109_,data_li_1__3__108_,
  data_li_1__3__107_,data_li_1__3__106_,data_li_1__3__105_,data_li_1__3__104_,
  data_li_1__3__103_,data_li_1__3__102_,data_li_1__3__101_,data_li_1__3__100_,
  data_li_1__3__99_,data_li_1__3__98_,data_li_1__3__97_,data_li_1__3__96_,data_li_1__3__95_,
  data_li_1__3__94_,data_li_1__3__93_,data_li_1__3__92_,data_li_1__3__91_,
  data_li_1__3__90_,data_li_1__3__89_,data_li_1__3__88_,data_li_1__3__87_,data_li_1__3__86_,
  data_li_1__3__85_,data_li_1__3__84_,data_li_1__3__83_,data_li_1__3__82_,
  data_li_1__3__81_,data_li_1__3__80_,data_li_1__3__79_,data_li_1__3__78_,data_li_1__3__77_,
  data_li_1__3__76_,data_li_1__3__75_,data_li_1__3__74_,data_li_1__3__73_,
  data_li_1__3__72_,data_li_1__3__71_,data_li_1__3__70_,data_li_1__3__69_,data_li_1__3__68_,
  data_li_1__3__67_,data_li_1__3__66_,data_li_1__3__65_,data_li_1__3__64_,
  data_li_1__3__63_,data_li_1__3__62_,data_li_1__3__61_,data_li_1__3__60_,
  data_li_1__3__59_,data_li_1__3__58_,data_li_1__3__57_,data_li_1__3__56_,data_li_1__3__55_,
  data_li_1__3__54_,data_li_1__3__53_,data_li_1__3__52_,data_li_1__3__51_,
  data_li_1__3__50_,data_li_1__3__49_,data_li_1__3__48_,data_li_1__3__47_,data_li_1__3__46_,
  data_li_1__3__45_,data_li_1__3__44_,data_li_1__3__43_,data_li_1__3__42_,
  data_li_1__3__41_,data_li_1__3__40_,data_li_1__3__39_,data_li_1__3__38_,data_li_1__3__37_,
  data_li_1__3__36_,data_li_1__3__35_,data_li_1__3__34_,data_li_1__3__33_,
  data_li_1__3__32_,data_li_1__3__31_,data_li_1__3__30_,data_li_1__3__29_,data_li_1__3__28_,
  data_li_1__3__27_,data_li_1__3__26_,data_li_1__3__25_,data_li_1__3__24_,
  data_li_1__3__23_,data_li_1__3__22_,data_li_1__3__21_,data_li_1__3__20_,
  data_li_1__3__19_,data_li_1__3__18_,data_li_1__3__17_,data_li_1__3__16_,data_li_1__3__15_,
  data_li_1__3__14_,data_li_1__3__13_,data_li_1__3__12_,data_li_1__3__11_,
  data_li_1__3__10_,data_li_1__3__9_,data_li_1__3__8_,data_li_1__3__7_,data_li_1__3__6_,
  data_li_1__3__5_,data_li_1__3__4_,data_li_1__3__3_,data_li_1__3__2_,data_li_1__3__1_,
  data_li_1__3__0_,data_li_1__2__130_,data_li_1__2__129_,data_li_1__2__128_,
  data_li_1__2__127_,data_li_1__2__126_,data_li_1__2__125_,data_li_1__2__124_,
  data_li_1__2__123_,data_li_1__2__122_,data_li_1__2__121_,data_li_1__2__120_,
  data_li_1__2__119_,data_li_1__2__118_,data_li_1__2__117_,data_li_1__2__116_,data_li_1__2__115_,
  data_li_1__2__114_,data_li_1__2__113_,data_li_1__2__112_,data_li_1__2__111_,
  data_li_1__2__110_,data_li_1__2__109_,data_li_1__2__108_,data_li_1__2__107_,
  data_li_1__2__106_,data_li_1__2__105_,data_li_1__2__104_,data_li_1__2__103_,
  data_li_1__2__102_,data_li_1__2__101_,data_li_1__2__100_,data_li_1__2__99_,data_li_1__2__98_,
  data_li_1__2__97_,data_li_1__2__96_,data_li_1__2__95_,data_li_1__2__94_,
  data_li_1__2__93_,data_li_1__2__92_,data_li_1__2__91_,data_li_1__2__90_,data_li_1__2__89_,
  data_li_1__2__88_,data_li_1__2__87_,data_li_1__2__86_,data_li_1__2__85_,
  data_li_1__2__84_,data_li_1__2__83_,data_li_1__2__82_,data_li_1__2__81_,
  data_li_1__2__80_,data_li_1__2__79_,data_li_1__2__78_,data_li_1__2__77_,data_li_1__2__76_,
  data_li_1__2__75_,data_li_1__2__74_,data_li_1__2__73_,data_li_1__2__72_,
  data_li_1__2__71_,data_li_1__2__70_,data_li_1__2__69_,data_li_1__2__68_,data_li_1__2__67_,
  data_li_1__2__66_,data_li_1__2__65_,data_li_1__2__64_,data_li_1__2__63_,
  data_li_1__2__62_,data_li_1__2__61_,data_li_1__2__60_,data_li_1__2__59_,data_li_1__2__58_,
  data_li_1__2__57_,data_li_1__2__56_,data_li_1__2__55_,data_li_1__2__54_,
  data_li_1__2__53_,data_li_1__2__52_,data_li_1__2__51_,data_li_1__2__50_,data_li_1__2__49_,
  data_li_1__2__48_,data_li_1__2__47_,data_li_1__2__46_,data_li_1__2__45_,
  data_li_1__2__44_,data_li_1__2__43_,data_li_1__2__42_,data_li_1__2__41_,
  data_li_1__2__40_,data_li_1__2__39_,data_li_1__2__38_,data_li_1__2__37_,data_li_1__2__36_,
  data_li_1__2__35_,data_li_1__2__34_,data_li_1__2__33_,data_li_1__2__32_,
  data_li_1__2__31_,data_li_1__2__30_,data_li_1__2__29_,data_li_1__2__28_,data_li_1__2__27_,
  data_li_1__2__26_,data_li_1__2__25_,data_li_1__2__24_,data_li_1__2__23_,
  data_li_1__2__22_,data_li_1__2__21_,data_li_1__2__20_,data_li_1__2__19_,data_li_1__2__18_,
  data_li_1__2__17_,data_li_1__2__16_,data_li_1__2__15_,data_li_1__2__14_,
  data_li_1__2__13_,data_li_1__2__12_,data_li_1__2__11_,data_li_1__2__10_,data_li_1__2__9_,
  data_li_1__2__8_,data_li_1__2__7_,data_li_1__2__6_,data_li_1__2__5_,
  data_li_1__2__4_,data_li_1__2__3_,data_li_1__2__2_,data_li_1__2__1_,data_li_1__2__0_,
  lce_packet_out_1__3_,lce_packet_out_1__2_,lce_packet_out_1__1_,lce_packet_out_1__0_,
  lce_packet_out_0__3_,lce_packet_out_0__2_,lce_packet_out_0__1_,lce_packet_out_0__0_;
  wire [9:0] ready_lo,valid_lo;
  wire [1309:0] data_lo;
  wire [1043:0] lce_packet_in;
  wire [521:0] cce_packet_in;

  bsg_wormhole_router_131_1_1_2_1_1_1_00000003_0000001a
  router_0__router
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .local_x_cord_i(1'b0),
    .local_y_cord_i(1'b1),
    .valid_i({ valid_li_0__4_, valid_li_0__3_, valid_lo[6:6], valid_li_0__1_, valid_li_0__0_ }),
    .data_i({ data_li_0__4__130_, data_li_0__4__129_, data_li_0__4__128_, data_li_0__4__127_, data_li_0__4__126_, data_li_0__4__125_, data_li_0__4__124_, data_li_0__4__123_, data_li_0__4__122_, data_li_0__4__121_, data_li_0__4__120_, data_li_0__4__119_, data_li_0__4__118_, data_li_0__4__117_, data_li_0__4__116_, data_li_0__4__115_, data_li_0__4__114_, data_li_0__4__113_, data_li_0__4__112_, data_li_0__4__111_, data_li_0__4__110_, data_li_0__4__109_, data_li_0__4__108_, data_li_0__4__107_, data_li_0__4__106_, data_li_0__4__105_, data_li_0__4__104_, data_li_0__4__103_, data_li_0__4__102_, data_li_0__4__101_, data_li_0__4__100_, data_li_0__4__99_, data_li_0__4__98_, data_li_0__4__97_, data_li_0__4__96_, data_li_0__4__95_, data_li_0__4__94_, data_li_0__4__93_, data_li_0__4__92_, data_li_0__4__91_, data_li_0__4__90_, data_li_0__4__89_, data_li_0__4__88_, data_li_0__4__87_, data_li_0__4__86_, data_li_0__4__85_, data_li_0__4__84_, data_li_0__4__83_, data_li_0__4__82_, data_li_0__4__81_, data_li_0__4__80_, data_li_0__4__79_, data_li_0__4__78_, data_li_0__4__77_, data_li_0__4__76_, data_li_0__4__75_, data_li_0__4__74_, data_li_0__4__73_, data_li_0__4__72_, data_li_0__4__71_, data_li_0__4__70_, data_li_0__4__69_, data_li_0__4__68_, data_li_0__4__67_, data_li_0__4__66_, data_li_0__4__65_, data_li_0__4__64_, data_li_0__4__63_, data_li_0__4__62_, data_li_0__4__61_, data_li_0__4__60_, data_li_0__4__59_, data_li_0__4__58_, data_li_0__4__57_, data_li_0__4__56_, data_li_0__4__55_, data_li_0__4__54_, data_li_0__4__53_, data_li_0__4__52_, data_li_0__4__51_, data_li_0__4__50_, data_li_0__4__49_, data_li_0__4__48_, data_li_0__4__47_, data_li_0__4__46_, data_li_0__4__45_, data_li_0__4__44_, data_li_0__4__43_, data_li_0__4__42_, data_li_0__4__41_, data_li_0__4__40_, data_li_0__4__39_, data_li_0__4__38_, data_li_0__4__37_, data_li_0__4__36_, data_li_0__4__35_, data_li_0__4__34_, data_li_0__4__33_, data_li_0__4__32_, data_li_0__4__31_, data_li_0__4__30_, data_li_0__4__29_, data_li_0__4__28_, data_li_0__4__27_, data_li_0__4__26_, data_li_0__4__25_, data_li_0__4__24_, data_li_0__4__23_, data_li_0__4__22_, data_li_0__4__21_, data_li_0__4__20_, data_li_0__4__19_, data_li_0__4__18_, data_li_0__4__17_, data_li_0__4__16_, data_li_0__4__15_, data_li_0__4__14_, data_li_0__4__13_, data_li_0__4__12_, data_li_0__4__11_, data_li_0__4__10_, data_li_0__4__9_, data_li_0__4__8_, data_li_0__4__7_, data_li_0__4__6_, data_li_0__4__5_, data_li_0__4__4_, data_li_0__4__3_, data_li_0__4__2_, data_li_0__4__1_, data_li_0__4__0_, data_li_0__3__130_, data_li_0__3__129_, data_li_0__3__128_, data_li_0__3__127_, data_li_0__3__126_, data_li_0__3__125_, data_li_0__3__124_, data_li_0__3__123_, data_li_0__3__122_, data_li_0__3__121_, data_li_0__3__120_, data_li_0__3__119_, data_li_0__3__118_, data_li_0__3__117_, data_li_0__3__116_, data_li_0__3__115_, data_li_0__3__114_, data_li_0__3__113_, data_li_0__3__112_, data_li_0__3__111_, data_li_0__3__110_, data_li_0__3__109_, data_li_0__3__108_, data_li_0__3__107_, data_li_0__3__106_, data_li_0__3__105_, data_li_0__3__104_, data_li_0__3__103_, data_li_0__3__102_, data_li_0__3__101_, data_li_0__3__100_, data_li_0__3__99_, data_li_0__3__98_, data_li_0__3__97_, data_li_0__3__96_, data_li_0__3__95_, data_li_0__3__94_, data_li_0__3__93_, data_li_0__3__92_, data_li_0__3__91_, data_li_0__3__90_, data_li_0__3__89_, data_li_0__3__88_, data_li_0__3__87_, data_li_0__3__86_, data_li_0__3__85_, data_li_0__3__84_, data_li_0__3__83_, data_li_0__3__82_, data_li_0__3__81_, data_li_0__3__80_, data_li_0__3__79_, data_li_0__3__78_, data_li_0__3__77_, data_li_0__3__76_, data_li_0__3__75_, data_li_0__3__74_, data_li_0__3__73_, data_li_0__3__72_, data_li_0__3__71_, data_li_0__3__70_, data_li_0__3__69_, data_li_0__3__68_, data_li_0__3__67_, data_li_0__3__66_, data_li_0__3__65_, data_li_0__3__64_, data_li_0__3__63_, data_li_0__3__62_, data_li_0__3__61_, data_li_0__3__60_, data_li_0__3__59_, data_li_0__3__58_, data_li_0__3__57_, data_li_0__3__56_, data_li_0__3__55_, data_li_0__3__54_, data_li_0__3__53_, data_li_0__3__52_, data_li_0__3__51_, data_li_0__3__50_, data_li_0__3__49_, data_li_0__3__48_, data_li_0__3__47_, data_li_0__3__46_, data_li_0__3__45_, data_li_0__3__44_, data_li_0__3__43_, data_li_0__3__42_, data_li_0__3__41_, data_li_0__3__40_, data_li_0__3__39_, data_li_0__3__38_, data_li_0__3__37_, data_li_0__3__36_, data_li_0__3__35_, data_li_0__3__34_, data_li_0__3__33_, data_li_0__3__32_, data_li_0__3__31_, data_li_0__3__30_, data_li_0__3__29_, data_li_0__3__28_, data_li_0__3__27_, data_li_0__3__26_, data_li_0__3__25_, data_li_0__3__24_, data_li_0__3__23_, data_li_0__3__22_, data_li_0__3__21_, data_li_0__3__20_, data_li_0__3__19_, data_li_0__3__18_, data_li_0__3__17_, data_li_0__3__16_, data_li_0__3__15_, data_li_0__3__14_, data_li_0__3__13_, data_li_0__3__12_, data_li_0__3__11_, data_li_0__3__10_, data_li_0__3__9_, data_li_0__3__8_, data_li_0__3__7_, data_li_0__3__6_, data_li_0__3__5_, data_li_0__3__4_, data_li_0__3__3_, data_li_0__3__2_, data_li_0__3__1_, data_li_0__3__0_, data_lo[916:786], data_li_0__1__130_, data_li_0__1__129_, data_li_0__1__128_, data_li_0__1__127_, data_li_0__1__126_, data_li_0__1__125_, data_li_0__1__124_, data_li_0__1__123_, data_li_0__1__122_, data_li_0__1__121_, data_li_0__1__120_, data_li_0__1__119_, data_li_0__1__118_, data_li_0__1__117_, data_li_0__1__116_, data_li_0__1__115_, data_li_0__1__114_, data_li_0__1__113_, data_li_0__1__112_, data_li_0__1__111_, data_li_0__1__110_, data_li_0__1__109_, data_li_0__1__108_, data_li_0__1__107_, data_li_0__1__106_, data_li_0__1__105_, data_li_0__1__104_, data_li_0__1__103_, data_li_0__1__102_, data_li_0__1__101_, data_li_0__1__100_, data_li_0__1__99_, data_li_0__1__98_, data_li_0__1__97_, data_li_0__1__96_, data_li_0__1__95_, data_li_0__1__94_, data_li_0__1__93_, data_li_0__1__92_, data_li_0__1__91_, data_li_0__1__90_, data_li_0__1__89_, data_li_0__1__88_, data_li_0__1__87_, data_li_0__1__86_, data_li_0__1__85_, data_li_0__1__84_, data_li_0__1__83_, data_li_0__1__82_, data_li_0__1__81_, data_li_0__1__80_, data_li_0__1__79_, data_li_0__1__78_, data_li_0__1__77_, data_li_0__1__76_, data_li_0__1__75_, data_li_0__1__74_, data_li_0__1__73_, data_li_0__1__72_, data_li_0__1__71_, data_li_0__1__70_, data_li_0__1__69_, data_li_0__1__68_, data_li_0__1__67_, data_li_0__1__66_, data_li_0__1__65_, data_li_0__1__64_, data_li_0__1__63_, data_li_0__1__62_, data_li_0__1__61_, data_li_0__1__60_, data_li_0__1__59_, data_li_0__1__58_, data_li_0__1__57_, data_li_0__1__56_, data_li_0__1__55_, data_li_0__1__54_, data_li_0__1__53_, data_li_0__1__52_, data_li_0__1__51_, data_li_0__1__50_, data_li_0__1__49_, data_li_0__1__48_, data_li_0__1__47_, data_li_0__1__46_, data_li_0__1__45_, data_li_0__1__44_, data_li_0__1__43_, data_li_0__1__42_, data_li_0__1__41_, data_li_0__1__40_, data_li_0__1__39_, data_li_0__1__38_, data_li_0__1__37_, data_li_0__1__36_, data_li_0__1__35_, data_li_0__1__34_, data_li_0__1__33_, data_li_0__1__32_, data_li_0__1__31_, data_li_0__1__30_, data_li_0__1__29_, data_li_0__1__28_, data_li_0__1__27_, data_li_0__1__26_, data_li_0__1__25_, data_li_0__1__24_, data_li_0__1__23_, data_li_0__1__22_, data_li_0__1__21_, data_li_0__1__20_, data_li_0__1__19_, data_li_0__1__18_, data_li_0__1__17_, data_li_0__1__16_, data_li_0__1__15_, data_li_0__1__14_, data_li_0__1__13_, data_li_0__1__12_, data_li_0__1__11_, data_li_0__1__10_, data_li_0__1__9_, data_li_0__1__8_, data_li_0__1__7_, data_li_0__1__6_, data_li_0__1__5_, data_li_0__1__4_, data_li_0__1__3_, data_li_0__1__2_, data_li_0__1__1_, data_li_0__1__0_, data_li_0__0__130_, data_li_0__0__129_, data_li_0__0__128_, data_li_0__0__127_, data_li_0__0__126_, data_li_0__0__125_, data_li_0__0__124_, data_li_0__0__123_, data_li_0__0__122_, data_li_0__0__121_, data_li_0__0__120_, data_li_0__0__119_, data_li_0__0__118_, data_li_0__0__117_, data_li_0__0__116_, data_li_0__0__115_, data_li_0__0__114_, data_li_0__0__113_, data_li_0__0__112_, data_li_0__0__111_, data_li_0__0__110_, data_li_0__0__109_, data_li_0__0__108_, data_li_0__0__107_, data_li_0__0__106_, data_li_0__0__105_, data_li_0__0__104_, data_li_0__0__103_, data_li_0__0__102_, data_li_0__0__101_, data_li_0__0__100_, data_li_0__0__99_, data_li_0__0__98_, data_li_0__0__97_, data_li_0__0__96_, data_li_0__0__95_, data_li_0__0__94_, data_li_0__0__93_, data_li_0__0__92_, data_li_0__0__91_, data_li_0__0__90_, data_li_0__0__89_, data_li_0__0__88_, data_li_0__0__87_, data_li_0__0__86_, data_li_0__0__85_, data_li_0__0__84_, data_li_0__0__83_, data_li_0__0__82_, data_li_0__0__81_, data_li_0__0__80_, data_li_0__0__79_, data_li_0__0__78_, data_li_0__0__77_, data_li_0__0__76_, data_li_0__0__75_, data_li_0__0__74_, data_li_0__0__73_, data_li_0__0__72_, data_li_0__0__71_, data_li_0__0__70_, data_li_0__0__69_, data_li_0__0__68_, data_li_0__0__67_, data_li_0__0__66_, data_li_0__0__65_, data_li_0__0__64_, data_li_0__0__63_, data_li_0__0__62_, data_li_0__0__61_, data_li_0__0__60_, data_li_0__0__59_, data_li_0__0__58_, data_li_0__0__57_, data_li_0__0__56_, data_li_0__0__55_, data_li_0__0__54_, data_li_0__0__53_, data_li_0__0__52_, data_li_0__0__51_, data_li_0__0__50_, data_li_0__0__49_, data_li_0__0__48_, data_li_0__0__47_, data_li_0__0__46_, data_li_0__0__45_, data_li_0__0__44_, data_li_0__0__43_, data_li_0__0__42_, data_li_0__0__41_, data_li_0__0__40_, data_li_0__0__39_, data_li_0__0__38_, data_li_0__0__37_, data_li_0__0__36_, data_li_0__0__35_, data_li_0__0__34_, data_li_0__0__33_, data_li_0__0__32_, data_li_0__0__31_, data_li_0__0__30_, data_li_0__0__29_, data_li_0__0__28_, data_li_0__0__27_, data_li_0__0__26_, data_li_0__0__25_, data_li_0__0__24_, data_li_0__0__23_, data_li_0__0__22_, data_li_0__0__21_, data_li_0__0__20_, data_li_0__0__19_, data_li_0__0__18_, data_li_0__0__17_, data_li_0__0__16_, data_li_0__0__15_, data_li_0__0__14_, data_li_0__0__13_, data_li_0__0__12_, data_li_0__0__11_, data_li_0__0__10_, data_li_0__0__9_, data_li_0__0__8_, data_li_0__0__7_, data_li_0__0__6_, data_li_0__0__5_, data_li_0__0__4_, data_li_0__0__3_, data_li_0__0__2_, data_li_0__0__1_, data_li_0__0__0_ }),
    .ready_o(ready_lo[4:0]),
    .valid_o(valid_lo[4:0]),
    .data_o(data_lo[654:0]),
    .ready_i({ ready_li_0__4_, ready_li_0__3_, ready_lo[6:6], ready_li_0__1_, ready_li_0__0_ })
  );


  bsg_wormhole_router_131_1_1_2_1_1_1_00000015_0000001c
  router_1__router
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .local_x_cord_i(1'b1),
    .local_y_cord_i(1'b1),
    .valid_i({ valid_li_1__4_, valid_li_1__3_, valid_li_1__2_, valid_lo[2:2], valid_li_1__0_ }),
    .data_i({ data_li_1__4__130_, data_li_1__4__129_, data_li_1__4__128_, data_li_1__4__127_, data_li_1__4__126_, data_li_1__4__125_, data_li_1__4__124_, data_li_1__4__123_, data_li_1__4__122_, data_li_1__4__121_, data_li_1__4__120_, data_li_1__4__119_, data_li_1__4__118_, data_li_1__4__117_, data_li_1__4__116_, data_li_1__4__115_, data_li_1__4__114_, data_li_1__4__113_, data_li_1__4__112_, data_li_1__4__111_, data_li_1__4__110_, data_li_1__4__109_, data_li_1__4__108_, data_li_1__4__107_, data_li_1__4__106_, data_li_1__4__105_, data_li_1__4__104_, data_li_1__4__103_, data_li_1__4__102_, data_li_1__4__101_, data_li_1__4__100_, data_li_1__4__99_, data_li_1__4__98_, data_li_1__4__97_, data_li_1__4__96_, data_li_1__4__95_, data_li_1__4__94_, data_li_1__4__93_, data_li_1__4__92_, data_li_1__4__91_, data_li_1__4__90_, data_li_1__4__89_, data_li_1__4__88_, data_li_1__4__87_, data_li_1__4__86_, data_li_1__4__85_, data_li_1__4__84_, data_li_1__4__83_, data_li_1__4__82_, data_li_1__4__81_, data_li_1__4__80_, data_li_1__4__79_, data_li_1__4__78_, data_li_1__4__77_, data_li_1__4__76_, data_li_1__4__75_, data_li_1__4__74_, data_li_1__4__73_, data_li_1__4__72_, data_li_1__4__71_, data_li_1__4__70_, data_li_1__4__69_, data_li_1__4__68_, data_li_1__4__67_, data_li_1__4__66_, data_li_1__4__65_, data_li_1__4__64_, data_li_1__4__63_, data_li_1__4__62_, data_li_1__4__61_, data_li_1__4__60_, data_li_1__4__59_, data_li_1__4__58_, data_li_1__4__57_, data_li_1__4__56_, data_li_1__4__55_, data_li_1__4__54_, data_li_1__4__53_, data_li_1__4__52_, data_li_1__4__51_, data_li_1__4__50_, data_li_1__4__49_, data_li_1__4__48_, data_li_1__4__47_, data_li_1__4__46_, data_li_1__4__45_, data_li_1__4__44_, data_li_1__4__43_, data_li_1__4__42_, data_li_1__4__41_, data_li_1__4__40_, data_li_1__4__39_, data_li_1__4__38_, data_li_1__4__37_, data_li_1__4__36_, data_li_1__4__35_, data_li_1__4__34_, data_li_1__4__33_, data_li_1__4__32_, data_li_1__4__31_, data_li_1__4__30_, data_li_1__4__29_, data_li_1__4__28_, data_li_1__4__27_, data_li_1__4__26_, data_li_1__4__25_, data_li_1__4__24_, data_li_1__4__23_, data_li_1__4__22_, data_li_1__4__21_, data_li_1__4__20_, data_li_1__4__19_, data_li_1__4__18_, data_li_1__4__17_, data_li_1__4__16_, data_li_1__4__15_, data_li_1__4__14_, data_li_1__4__13_, data_li_1__4__12_, data_li_1__4__11_, data_li_1__4__10_, data_li_1__4__9_, data_li_1__4__8_, data_li_1__4__7_, data_li_1__4__6_, data_li_1__4__5_, data_li_1__4__4_, data_li_1__4__3_, data_li_1__4__2_, data_li_1__4__1_, data_li_1__4__0_, data_li_1__3__130_, data_li_1__3__129_, data_li_1__3__128_, data_li_1__3__127_, data_li_1__3__126_, data_li_1__3__125_, data_li_1__3__124_, data_li_1__3__123_, data_li_1__3__122_, data_li_1__3__121_, data_li_1__3__120_, data_li_1__3__119_, data_li_1__3__118_, data_li_1__3__117_, data_li_1__3__116_, data_li_1__3__115_, data_li_1__3__114_, data_li_1__3__113_, data_li_1__3__112_, data_li_1__3__111_, data_li_1__3__110_, data_li_1__3__109_, data_li_1__3__108_, data_li_1__3__107_, data_li_1__3__106_, data_li_1__3__105_, data_li_1__3__104_, data_li_1__3__103_, data_li_1__3__102_, data_li_1__3__101_, data_li_1__3__100_, data_li_1__3__99_, data_li_1__3__98_, data_li_1__3__97_, data_li_1__3__96_, data_li_1__3__95_, data_li_1__3__94_, data_li_1__3__93_, data_li_1__3__92_, data_li_1__3__91_, data_li_1__3__90_, data_li_1__3__89_, data_li_1__3__88_, data_li_1__3__87_, data_li_1__3__86_, data_li_1__3__85_, data_li_1__3__84_, data_li_1__3__83_, data_li_1__3__82_, data_li_1__3__81_, data_li_1__3__80_, data_li_1__3__79_, data_li_1__3__78_, data_li_1__3__77_, data_li_1__3__76_, data_li_1__3__75_, data_li_1__3__74_, data_li_1__3__73_, data_li_1__3__72_, data_li_1__3__71_, data_li_1__3__70_, data_li_1__3__69_, data_li_1__3__68_, data_li_1__3__67_, data_li_1__3__66_, data_li_1__3__65_, data_li_1__3__64_, data_li_1__3__63_, data_li_1__3__62_, data_li_1__3__61_, data_li_1__3__60_, data_li_1__3__59_, data_li_1__3__58_, data_li_1__3__57_, data_li_1__3__56_, data_li_1__3__55_, data_li_1__3__54_, data_li_1__3__53_, data_li_1__3__52_, data_li_1__3__51_, data_li_1__3__50_, data_li_1__3__49_, data_li_1__3__48_, data_li_1__3__47_, data_li_1__3__46_, data_li_1__3__45_, data_li_1__3__44_, data_li_1__3__43_, data_li_1__3__42_, data_li_1__3__41_, data_li_1__3__40_, data_li_1__3__39_, data_li_1__3__38_, data_li_1__3__37_, data_li_1__3__36_, data_li_1__3__35_, data_li_1__3__34_, data_li_1__3__33_, data_li_1__3__32_, data_li_1__3__31_, data_li_1__3__30_, data_li_1__3__29_, data_li_1__3__28_, data_li_1__3__27_, data_li_1__3__26_, data_li_1__3__25_, data_li_1__3__24_, data_li_1__3__23_, data_li_1__3__22_, data_li_1__3__21_, data_li_1__3__20_, data_li_1__3__19_, data_li_1__3__18_, data_li_1__3__17_, data_li_1__3__16_, data_li_1__3__15_, data_li_1__3__14_, data_li_1__3__13_, data_li_1__3__12_, data_li_1__3__11_, data_li_1__3__10_, data_li_1__3__9_, data_li_1__3__8_, data_li_1__3__7_, data_li_1__3__6_, data_li_1__3__5_, data_li_1__3__4_, data_li_1__3__3_, data_li_1__3__2_, data_li_1__3__1_, data_li_1__3__0_, data_li_1__2__130_, data_li_1__2__129_, data_li_1__2__128_, data_li_1__2__127_, data_li_1__2__126_, data_li_1__2__125_, data_li_1__2__124_, data_li_1__2__123_, data_li_1__2__122_, data_li_1__2__121_, data_li_1__2__120_, data_li_1__2__119_, data_li_1__2__118_, data_li_1__2__117_, data_li_1__2__116_, data_li_1__2__115_, data_li_1__2__114_, data_li_1__2__113_, data_li_1__2__112_, data_li_1__2__111_, data_li_1__2__110_, data_li_1__2__109_, data_li_1__2__108_, data_li_1__2__107_, data_li_1__2__106_, data_li_1__2__105_, data_li_1__2__104_, data_li_1__2__103_, data_li_1__2__102_, data_li_1__2__101_, data_li_1__2__100_, data_li_1__2__99_, data_li_1__2__98_, data_li_1__2__97_, data_li_1__2__96_, data_li_1__2__95_, data_li_1__2__94_, data_li_1__2__93_, data_li_1__2__92_, data_li_1__2__91_, data_li_1__2__90_, data_li_1__2__89_, data_li_1__2__88_, data_li_1__2__87_, data_li_1__2__86_, data_li_1__2__85_, data_li_1__2__84_, data_li_1__2__83_, data_li_1__2__82_, data_li_1__2__81_, data_li_1__2__80_, data_li_1__2__79_, data_li_1__2__78_, data_li_1__2__77_, data_li_1__2__76_, data_li_1__2__75_, data_li_1__2__74_, data_li_1__2__73_, data_li_1__2__72_, data_li_1__2__71_, data_li_1__2__70_, data_li_1__2__69_, data_li_1__2__68_, data_li_1__2__67_, data_li_1__2__66_, data_li_1__2__65_, data_li_1__2__64_, data_li_1__2__63_, data_li_1__2__62_, data_li_1__2__61_, data_li_1__2__60_, data_li_1__2__59_, data_li_1__2__58_, data_li_1__2__57_, data_li_1__2__56_, data_li_1__2__55_, data_li_1__2__54_, data_li_1__2__53_, data_li_1__2__52_, data_li_1__2__51_, data_li_1__2__50_, data_li_1__2__49_, data_li_1__2__48_, data_li_1__2__47_, data_li_1__2__46_, data_li_1__2__45_, data_li_1__2__44_, data_li_1__2__43_, data_li_1__2__42_, data_li_1__2__41_, data_li_1__2__40_, data_li_1__2__39_, data_li_1__2__38_, data_li_1__2__37_, data_li_1__2__36_, data_li_1__2__35_, data_li_1__2__34_, data_li_1__2__33_, data_li_1__2__32_, data_li_1__2__31_, data_li_1__2__30_, data_li_1__2__29_, data_li_1__2__28_, data_li_1__2__27_, data_li_1__2__26_, data_li_1__2__25_, data_li_1__2__24_, data_li_1__2__23_, data_li_1__2__22_, data_li_1__2__21_, data_li_1__2__20_, data_li_1__2__19_, data_li_1__2__18_, data_li_1__2__17_, data_li_1__2__16_, data_li_1__2__15_, data_li_1__2__14_, data_li_1__2__13_, data_li_1__2__12_, data_li_1__2__11_, data_li_1__2__10_, data_li_1__2__9_, data_li_1__2__8_, data_li_1__2__7_, data_li_1__2__6_, data_li_1__2__5_, data_li_1__2__4_, data_li_1__2__3_, data_li_1__2__2_, data_li_1__2__1_, data_li_1__2__0_, data_lo[392:262], data_li_1__0__130_, data_li_1__0__129_, data_li_1__0__128_, data_li_1__0__127_, data_li_1__0__126_, data_li_1__0__125_, data_li_1__0__124_, data_li_1__0__123_, data_li_1__0__122_, data_li_1__0__121_, data_li_1__0__120_, data_li_1__0__119_, data_li_1__0__118_, data_li_1__0__117_, data_li_1__0__116_, data_li_1__0__115_, data_li_1__0__114_, data_li_1__0__113_, data_li_1__0__112_, data_li_1__0__111_, data_li_1__0__110_, data_li_1__0__109_, data_li_1__0__108_, data_li_1__0__107_, data_li_1__0__106_, data_li_1__0__105_, data_li_1__0__104_, data_li_1__0__103_, data_li_1__0__102_, data_li_1__0__101_, data_li_1__0__100_, data_li_1__0__99_, data_li_1__0__98_, data_li_1__0__97_, data_li_1__0__96_, data_li_1__0__95_, data_li_1__0__94_, data_li_1__0__93_, data_li_1__0__92_, data_li_1__0__91_, data_li_1__0__90_, data_li_1__0__89_, data_li_1__0__88_, data_li_1__0__87_, data_li_1__0__86_, data_li_1__0__85_, data_li_1__0__84_, data_li_1__0__83_, data_li_1__0__82_, data_li_1__0__81_, data_li_1__0__80_, data_li_1__0__79_, data_li_1__0__78_, data_li_1__0__77_, data_li_1__0__76_, data_li_1__0__75_, data_li_1__0__74_, data_li_1__0__73_, data_li_1__0__72_, data_li_1__0__71_, data_li_1__0__70_, data_li_1__0__69_, data_li_1__0__68_, data_li_1__0__67_, data_li_1__0__66_, data_li_1__0__65_, data_li_1__0__64_, data_li_1__0__63_, data_li_1__0__62_, data_li_1__0__61_, data_li_1__0__60_, data_li_1__0__59_, data_li_1__0__58_, data_li_1__0__57_, data_li_1__0__56_, data_li_1__0__55_, data_li_1__0__54_, data_li_1__0__53_, data_li_1__0__52_, data_li_1__0__51_, data_li_1__0__50_, data_li_1__0__49_, data_li_1__0__48_, data_li_1__0__47_, data_li_1__0__46_, data_li_1__0__45_, data_li_1__0__44_, data_li_1__0__43_, data_li_1__0__42_, data_li_1__0__41_, data_li_1__0__40_, data_li_1__0__39_, data_li_1__0__38_, data_li_1__0__37_, data_li_1__0__36_, data_li_1__0__35_, data_li_1__0__34_, data_li_1__0__33_, data_li_1__0__32_, data_li_1__0__31_, data_li_1__0__30_, data_li_1__0__29_, data_li_1__0__28_, data_li_1__0__27_, data_li_1__0__26_, data_li_1__0__25_, data_li_1__0__24_, data_li_1__0__23_, data_li_1__0__22_, data_li_1__0__21_, data_li_1__0__20_, data_li_1__0__19_, data_li_1__0__18_, data_li_1__0__17_, data_li_1__0__16_, data_li_1__0__15_, data_li_1__0__14_, data_li_1__0__13_, data_li_1__0__12_, data_li_1__0__11_, data_li_1__0__10_, data_li_1__0__9_, data_li_1__0__8_, data_li_1__0__7_, data_li_1__0__6_, data_li_1__0__5_, data_li_1__0__4_, data_li_1__0__3_, data_li_1__0__2_, data_li_1__0__1_, data_li_1__0__0_ }),
    .ready_o(ready_lo[9:5]),
    .valid_o(valid_lo[9:5]),
    .data_o(data_lo[1309:655]),
    .ready_i({ ready_li_1__4_, ready_li_1__3_, ready_li_1__2_, ready_lo[2:2], ready_li_1__0_ })
  );


  bp_me_network_pkt_encode_data_cmd_num_lce_p2_lce_assoc_p8_block_size_in_bits_p512_max_num_flit_p4_x_cord_width_p1_y_cord_width_p1
  genblk3_0__lce_pkt_encode
  (
    .payload_i(lce_lce_data_cmd_i[517:0]),
    .packet_o(lce_packet_in[521:0])
  );


  bp_me_network_pkt_encode_data_cmd_num_lce_p2_lce_assoc_p8_block_size_in_bits_p512_max_num_flit_p4_x_cord_width_p1_y_cord_width_p1
  genblk3_1__lce_pkt_encode
  (
    .payload_i(lce_lce_data_cmd_i[1035:518]),
    .packet_o(lce_packet_in[1043:522])
  );


  bsg_wormhole_router_adapter_in_max_num_flit_p4_max_payload_width_p518_x_cord_width_p1_y_cord_width_p1
  genblk4_0__lce_adapter_in
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(lce_packet_in[521:0]),
    .v_i(lce_lce_data_cmd_v_i[0]),
    .ready_o(lce_lce_data_cmd_ready_o[0]),
    .data_o({ data_li_0__3__130_, data_li_0__3__129_, data_li_0__3__128_, data_li_0__3__127_, data_li_0__3__126_, data_li_0__3__125_, data_li_0__3__124_, data_li_0__3__123_, data_li_0__3__122_, data_li_0__3__121_, data_li_0__3__120_, data_li_0__3__119_, data_li_0__3__118_, data_li_0__3__117_, data_li_0__3__116_, data_li_0__3__115_, data_li_0__3__114_, data_li_0__3__113_, data_li_0__3__112_, data_li_0__3__111_, data_li_0__3__110_, data_li_0__3__109_, data_li_0__3__108_, data_li_0__3__107_, data_li_0__3__106_, data_li_0__3__105_, data_li_0__3__104_, data_li_0__3__103_, data_li_0__3__102_, data_li_0__3__101_, data_li_0__3__100_, data_li_0__3__99_, data_li_0__3__98_, data_li_0__3__97_, data_li_0__3__96_, data_li_0__3__95_, data_li_0__3__94_, data_li_0__3__93_, data_li_0__3__92_, data_li_0__3__91_, data_li_0__3__90_, data_li_0__3__89_, data_li_0__3__88_, data_li_0__3__87_, data_li_0__3__86_, data_li_0__3__85_, data_li_0__3__84_, data_li_0__3__83_, data_li_0__3__82_, data_li_0__3__81_, data_li_0__3__80_, data_li_0__3__79_, data_li_0__3__78_, data_li_0__3__77_, data_li_0__3__76_, data_li_0__3__75_, data_li_0__3__74_, data_li_0__3__73_, data_li_0__3__72_, data_li_0__3__71_, data_li_0__3__70_, data_li_0__3__69_, data_li_0__3__68_, data_li_0__3__67_, data_li_0__3__66_, data_li_0__3__65_, data_li_0__3__64_, data_li_0__3__63_, data_li_0__3__62_, data_li_0__3__61_, data_li_0__3__60_, data_li_0__3__59_, data_li_0__3__58_, data_li_0__3__57_, data_li_0__3__56_, data_li_0__3__55_, data_li_0__3__54_, data_li_0__3__53_, data_li_0__3__52_, data_li_0__3__51_, data_li_0__3__50_, data_li_0__3__49_, data_li_0__3__48_, data_li_0__3__47_, data_li_0__3__46_, data_li_0__3__45_, data_li_0__3__44_, data_li_0__3__43_, data_li_0__3__42_, data_li_0__3__41_, data_li_0__3__40_, data_li_0__3__39_, data_li_0__3__38_, data_li_0__3__37_, data_li_0__3__36_, data_li_0__3__35_, data_li_0__3__34_, data_li_0__3__33_, data_li_0__3__32_, data_li_0__3__31_, data_li_0__3__30_, data_li_0__3__29_, data_li_0__3__28_, data_li_0__3__27_, data_li_0__3__26_, data_li_0__3__25_, data_li_0__3__24_, data_li_0__3__23_, data_li_0__3__22_, data_li_0__3__21_, data_li_0__3__20_, data_li_0__3__19_, data_li_0__3__18_, data_li_0__3__17_, data_li_0__3__16_, data_li_0__3__15_, data_li_0__3__14_, data_li_0__3__13_, data_li_0__3__12_, data_li_0__3__11_, data_li_0__3__10_, data_li_0__3__9_, data_li_0__3__8_, data_li_0__3__7_, data_li_0__3__6_, data_li_0__3__5_, data_li_0__3__4_, data_li_0__3__3_, data_li_0__3__2_, data_li_0__3__1_, data_li_0__3__0_ }),
    .v_o(valid_li_0__3_),
    .ready_i(ready_lo[3])
  );


  bsg_wormhole_router_adapter_in_max_num_flit_p4_max_payload_width_p518_x_cord_width_p1_y_cord_width_p1
  genblk4_1__lce_adapter_in
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(lce_packet_in[1043:522]),
    .v_i(lce_lce_data_cmd_v_i[1]),
    .ready_o(lce_lce_data_cmd_ready_o[1]),
    .data_o({ data_li_1__3__130_, data_li_1__3__129_, data_li_1__3__128_, data_li_1__3__127_, data_li_1__3__126_, data_li_1__3__125_, data_li_1__3__124_, data_li_1__3__123_, data_li_1__3__122_, data_li_1__3__121_, data_li_1__3__120_, data_li_1__3__119_, data_li_1__3__118_, data_li_1__3__117_, data_li_1__3__116_, data_li_1__3__115_, data_li_1__3__114_, data_li_1__3__113_, data_li_1__3__112_, data_li_1__3__111_, data_li_1__3__110_, data_li_1__3__109_, data_li_1__3__108_, data_li_1__3__107_, data_li_1__3__106_, data_li_1__3__105_, data_li_1__3__104_, data_li_1__3__103_, data_li_1__3__102_, data_li_1__3__101_, data_li_1__3__100_, data_li_1__3__99_, data_li_1__3__98_, data_li_1__3__97_, data_li_1__3__96_, data_li_1__3__95_, data_li_1__3__94_, data_li_1__3__93_, data_li_1__3__92_, data_li_1__3__91_, data_li_1__3__90_, data_li_1__3__89_, data_li_1__3__88_, data_li_1__3__87_, data_li_1__3__86_, data_li_1__3__85_, data_li_1__3__84_, data_li_1__3__83_, data_li_1__3__82_, data_li_1__3__81_, data_li_1__3__80_, data_li_1__3__79_, data_li_1__3__78_, data_li_1__3__77_, data_li_1__3__76_, data_li_1__3__75_, data_li_1__3__74_, data_li_1__3__73_, data_li_1__3__72_, data_li_1__3__71_, data_li_1__3__70_, data_li_1__3__69_, data_li_1__3__68_, data_li_1__3__67_, data_li_1__3__66_, data_li_1__3__65_, data_li_1__3__64_, data_li_1__3__63_, data_li_1__3__62_, data_li_1__3__61_, data_li_1__3__60_, data_li_1__3__59_, data_li_1__3__58_, data_li_1__3__57_, data_li_1__3__56_, data_li_1__3__55_, data_li_1__3__54_, data_li_1__3__53_, data_li_1__3__52_, data_li_1__3__51_, data_li_1__3__50_, data_li_1__3__49_, data_li_1__3__48_, data_li_1__3__47_, data_li_1__3__46_, data_li_1__3__45_, data_li_1__3__44_, data_li_1__3__43_, data_li_1__3__42_, data_li_1__3__41_, data_li_1__3__40_, data_li_1__3__39_, data_li_1__3__38_, data_li_1__3__37_, data_li_1__3__36_, data_li_1__3__35_, data_li_1__3__34_, data_li_1__3__33_, data_li_1__3__32_, data_li_1__3__31_, data_li_1__3__30_, data_li_1__3__29_, data_li_1__3__28_, data_li_1__3__27_, data_li_1__3__26_, data_li_1__3__25_, data_li_1__3__24_, data_li_1__3__23_, data_li_1__3__22_, data_li_1__3__21_, data_li_1__3__20_, data_li_1__3__19_, data_li_1__3__18_, data_li_1__3__17_, data_li_1__3__16_, data_li_1__3__15_, data_li_1__3__14_, data_li_1__3__13_, data_li_1__3__12_, data_li_1__3__11_, data_li_1__3__10_, data_li_1__3__9_, data_li_1__3__8_, data_li_1__3__7_, data_li_1__3__6_, data_li_1__3__5_, data_li_1__3__4_, data_li_1__3__3_, data_li_1__3__2_, data_li_1__3__1_, data_li_1__3__0_ }),
    .v_o(valid_li_1__3_),
    .ready_i(ready_lo[8])
  );


  bp_me_network_pkt_encode_data_cmd_num_lce_p2_lce_assoc_p8_block_size_in_bits_p512_max_num_flit_p4_x_cord_width_p1_y_cord_width_p1
  genblk5_0__cce_pkt_encode
  (
    .payload_i(cce_lce_data_cmd_i),
    .packet_o(cce_packet_in)
  );


  bsg_wormhole_router_adapter_in_max_num_flit_p4_max_payload_width_p518_x_cord_width_p1_y_cord_width_p1
  genblk6_0__cce_adapter_in
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(cce_packet_in),
    .v_i(cce_lce_data_cmd_v_i[0]),
    .ready_o(cce_lce_data_cmd_ready_o[0]),
    .data_o({ data_li_0__4__130_, data_li_0__4__129_, data_li_0__4__128_, data_li_0__4__127_, data_li_0__4__126_, data_li_0__4__125_, data_li_0__4__124_, data_li_0__4__123_, data_li_0__4__122_, data_li_0__4__121_, data_li_0__4__120_, data_li_0__4__119_, data_li_0__4__118_, data_li_0__4__117_, data_li_0__4__116_, data_li_0__4__115_, data_li_0__4__114_, data_li_0__4__113_, data_li_0__4__112_, data_li_0__4__111_, data_li_0__4__110_, data_li_0__4__109_, data_li_0__4__108_, data_li_0__4__107_, data_li_0__4__106_, data_li_0__4__105_, data_li_0__4__104_, data_li_0__4__103_, data_li_0__4__102_, data_li_0__4__101_, data_li_0__4__100_, data_li_0__4__99_, data_li_0__4__98_, data_li_0__4__97_, data_li_0__4__96_, data_li_0__4__95_, data_li_0__4__94_, data_li_0__4__93_, data_li_0__4__92_, data_li_0__4__91_, data_li_0__4__90_, data_li_0__4__89_, data_li_0__4__88_, data_li_0__4__87_, data_li_0__4__86_, data_li_0__4__85_, data_li_0__4__84_, data_li_0__4__83_, data_li_0__4__82_, data_li_0__4__81_, data_li_0__4__80_, data_li_0__4__79_, data_li_0__4__78_, data_li_0__4__77_, data_li_0__4__76_, data_li_0__4__75_, data_li_0__4__74_, data_li_0__4__73_, data_li_0__4__72_, data_li_0__4__71_, data_li_0__4__70_, data_li_0__4__69_, data_li_0__4__68_, data_li_0__4__67_, data_li_0__4__66_, data_li_0__4__65_, data_li_0__4__64_, data_li_0__4__63_, data_li_0__4__62_, data_li_0__4__61_, data_li_0__4__60_, data_li_0__4__59_, data_li_0__4__58_, data_li_0__4__57_, data_li_0__4__56_, data_li_0__4__55_, data_li_0__4__54_, data_li_0__4__53_, data_li_0__4__52_, data_li_0__4__51_, data_li_0__4__50_, data_li_0__4__49_, data_li_0__4__48_, data_li_0__4__47_, data_li_0__4__46_, data_li_0__4__45_, data_li_0__4__44_, data_li_0__4__43_, data_li_0__4__42_, data_li_0__4__41_, data_li_0__4__40_, data_li_0__4__39_, data_li_0__4__38_, data_li_0__4__37_, data_li_0__4__36_, data_li_0__4__35_, data_li_0__4__34_, data_li_0__4__33_, data_li_0__4__32_, data_li_0__4__31_, data_li_0__4__30_, data_li_0__4__29_, data_li_0__4__28_, data_li_0__4__27_, data_li_0__4__26_, data_li_0__4__25_, data_li_0__4__24_, data_li_0__4__23_, data_li_0__4__22_, data_li_0__4__21_, data_li_0__4__20_, data_li_0__4__19_, data_li_0__4__18_, data_li_0__4__17_, data_li_0__4__16_, data_li_0__4__15_, data_li_0__4__14_, data_li_0__4__13_, data_li_0__4__12_, data_li_0__4__11_, data_li_0__4__10_, data_li_0__4__9_, data_li_0__4__8_, data_li_0__4__7_, data_li_0__4__6_, data_li_0__4__5_, data_li_0__4__4_, data_li_0__4__3_, data_li_0__4__2_, data_li_0__4__1_, data_li_0__4__0_ }),
    .v_o(valid_li_0__4_),
    .ready_i(ready_lo[4])
  );


  bsg_wormhole_router_adapter_out_max_num_flit_p4_max_payload_width_p518_x_cord_width_p1_y_cord_width_p1
  genblk7_0__adapter_out
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_lo[130:0]),
    .v_i(valid_lo[0]),
    .ready_o(ready_li_0__0_),
    .data_o({ lce_data_cmd_o[517:0], lce_packet_out_0__3_, lce_packet_out_0__2_, lce_packet_out_0__1_, lce_packet_out_0__0_ }),
    .v_o(lce_data_cmd_v_o[0]),
    .ready_i(lce_data_cmd_ready_i[0])
  );


  bsg_wormhole_router_adapter_out_max_num_flit_p4_max_payload_width_p518_x_cord_width_p1_y_cord_width_p1
  genblk7_1__adapter_out
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_lo[785:655]),
    .v_i(valid_lo[5]),
    .ready_o(ready_li_1__0_),
    .data_o({ lce_data_cmd_o[1035:518], lce_packet_out_1__3_, lce_packet_out_1__2_, lce_packet_out_1__1_, lce_packet_out_1__0_ }),
    .v_o(lce_data_cmd_v_o[1]),
    .ready_i(lce_data_cmd_ready_i[1])
  );


endmodule



module bp_me_network_num_lce_p2_num_cce_p1_paddr_width_p22_lce_assoc_p8_block_size_in_bytes_p64_data_width_p64
(
  clk_i,
  reset_i,
  lce_cmd_o,
  lce_cmd_v_o,
  lce_cmd_ready_i,
  lce_cmd_i,
  lce_cmd_v_i,
  lce_cmd_ready_o,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i,
  cce_lce_data_cmd_i,
  cce_lce_data_cmd_v_i,
  cce_lce_data_cmd_ready_o,
  lce_lce_data_cmd_i,
  lce_lce_data_cmd_v_i,
  lce_lce_data_cmd_ready_o,
  lce_req_i,
  lce_req_v_i,
  lce_req_ready_o,
  lce_req_o,
  lce_req_v_o,
  lce_req_ready_i,
  lce_resp_i,
  lce_resp_v_i,
  lce_resp_ready_o,
  lce_resp_o,
  lce_resp_v_o,
  lce_resp_ready_i,
  lce_data_resp_i,
  lce_data_resp_v_i,
  lce_data_resp_ready_o,
  lce_data_resp_o,
  lce_data_resp_v_o,
  lce_data_resp_ready_i
);

  output [71:0] lce_cmd_o;
  output [1:0] lce_cmd_v_o;
  input [1:0] lce_cmd_ready_i;
  input [35:0] lce_cmd_i;
  input [0:0] lce_cmd_v_i;
  output [0:0] lce_cmd_ready_o;
  output [1035:0] lce_data_cmd_o;
  output [1:0] lce_data_cmd_v_o;
  input [1:0] lce_data_cmd_ready_i;
  input [517:0] cce_lce_data_cmd_i;
  input [0:0] cce_lce_data_cmd_v_i;
  output [0:0] cce_lce_data_cmd_ready_o;
  input [1035:0] lce_lce_data_cmd_i;
  input [1:0] lce_lce_data_cmd_v_i;
  output [1:0] lce_lce_data_cmd_ready_o;
  input [193:0] lce_req_i;
  input [1:0] lce_req_v_i;
  output [1:0] lce_req_ready_o;
  output [96:0] lce_req_o;
  output [0:0] lce_req_v_o;
  input [0:0] lce_req_ready_i;
  input [51:0] lce_resp_i;
  input [1:0] lce_resp_v_i;
  output [1:0] lce_resp_ready_o;
  output [25:0] lce_resp_o;
  output [0:0] lce_resp_v_o;
  input [0:0] lce_resp_ready_i;
  input [1073:0] lce_data_resp_i;
  input [1:0] lce_data_resp_v_i;
  output [1:0] lce_data_resp_ready_o;
  output [536:0] lce_data_resp_o;
  output [0:0] lce_data_resp_v_o;
  input [0:0] lce_data_resp_ready_i;
  input clk_i;
  input reset_i;
  wire [71:0] lce_cmd_o;
  wire [1:0] lce_cmd_v_o,lce_data_cmd_v_o,lce_lce_data_cmd_ready_o,lce_req_ready_o,
  lce_resp_ready_o,lce_data_resp_ready_o;
  wire [0:0] lce_cmd_ready_o,cce_lce_data_cmd_ready_o,lce_req_v_o,lce_resp_v_o,
  lce_data_resp_v_o;
  wire [1035:0] lce_data_cmd_o;
  wire [96:0] lce_req_o;
  wire [25:0] lce_resp_o;
  wire [536:0] lce_data_resp_o;

  bp_me_network_channel_mesh_packet_width_p36_num_src_p1_num_dst_p2_debug_p0
  cce_lce_cmd_network
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .src_data_i(lce_cmd_i),
    .src_v_i(lce_cmd_v_i[0]),
    .src_ready_o(lce_cmd_ready_o[0]),
    .dst_data_o(lce_cmd_o),
    .dst_v_o(lce_cmd_v_o),
    .dst_ready_i(lce_cmd_ready_i)
  );


  bp_me_network_channel_mesh_packet_width_p97_num_src_p2_num_dst_p1_debug_p0
  lce_cce_req_network
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .src_data_i(lce_req_i),
    .src_v_i(lce_req_v_i),
    .src_ready_o(lce_req_ready_o),
    .dst_data_o(lce_req_o),
    .dst_v_o(lce_req_v_o[0]),
    .dst_ready_i(lce_req_ready_i[0])
  );


  bp_me_network_channel_mesh_packet_width_p26_num_src_p2_num_dst_p1_debug_p0
  lce_cce_resp_network
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .src_data_i(lce_resp_i),
    .src_v_i(lce_resp_v_i),
    .src_ready_o(lce_resp_ready_o),
    .dst_data_o(lce_resp_o),
    .dst_v_o(lce_resp_v_o[0]),
    .dst_ready_i(lce_resp_ready_i[0])
  );


  bp_me_network_channel_data_resp_num_lce_p2_num_cce_p1_paddr_width_p22_block_size_in_bits_p512_max_num_flit_p4
  data_resp_channel
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .lce_data_resp_i(lce_data_resp_i),
    .lce_data_resp_v_i(lce_data_resp_v_i),
    .lce_data_resp_ready_o(lce_data_resp_ready_o),
    .lce_data_resp_o(lce_data_resp_o),
    .lce_data_resp_v_o(lce_data_resp_v_o[0]),
    .lce_data_resp_ready_i(lce_data_resp_ready_i[0])
  );


  bp_me_network_channel_data_cmd_num_lce_p2_num_cce_p1_lce_assoc_p8_block_size_in_bits_p512_max_num_flit_p4
  data_cmd_channel
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .lce_data_cmd_o(lce_data_cmd_o),
    .lce_data_cmd_v_o(lce_data_cmd_v_o),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_i),
    .cce_lce_data_cmd_i(cce_lce_data_cmd_i),
    .cce_lce_data_cmd_v_i(cce_lce_data_cmd_v_i[0]),
    .cce_lce_data_cmd_ready_o(cce_lce_data_cmd_ready_o[0]),
    .lce_lce_data_cmd_i(lce_lce_data_cmd_i),
    .lce_lce_data_cmd_v_i(lce_lce_data_cmd_v_i),
    .lce_lce_data_cmd_ready_o(lce_lce_data_cmd_ready_o)
  );


endmodule



module bsg_mem_p97
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [96:0] w_data_i;
  input [0:0] r_addr_i;
  output [96:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [96:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  reg [193:0] mem;
  assign r_data_o[96] = (N3)? mem[96] :
                        (N0)? mem[193] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[95] = (N3)? mem[95] :
                        (N0)? mem[192] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] :
                        (N0)? mem[191] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] :
                        (N0)? mem[190] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] :
                        (N0)? mem[189] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] :
                        (N0)? mem[188] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] :
                        (N0)? mem[187] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] :
                        (N0)? mem[186] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] :
                        (N0)? mem[185] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] :
                        (N0)? mem[184] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] :
                        (N0)? mem[183] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] :
                        (N0)? mem[182] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] :
                        (N0)? mem[181] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] :
                        (N0)? mem[180] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] :
                        (N0)? mem[179] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] :
                        (N0)? mem[178] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] :
                        (N0)? mem[177] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] :
                        (N0)? mem[176] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] :
                        (N0)? mem[175] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] :
                        (N0)? mem[174] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] :
                        (N0)? mem[173] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] :
                        (N0)? mem[172] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] :
                        (N0)? mem[171] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] :
                        (N0)? mem[170] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] :
                        (N0)? mem[169] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] :
                        (N0)? mem[168] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] :
                        (N0)? mem[167] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] :
                        (N0)? mem[166] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] :
                        (N0)? mem[165] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] :
                        (N0)? mem[164] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] :
                        (N0)? mem[163] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] :
                        (N0)? mem[162] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] :
                        (N0)? mem[161] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] :
                        (N0)? mem[160] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] :
                        (N0)? mem[159] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] :
                        (N0)? mem[158] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] :
                        (N0)? mem[157] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] :
                        (N0)? mem[156] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] :
                        (N0)? mem[155] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] :
                        (N0)? mem[154] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] :
                        (N0)? mem[153] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] :
                        (N0)? mem[152] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] :
                        (N0)? mem[151] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] :
                        (N0)? mem[150] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] :
                        (N0)? mem[149] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] :
                        (N0)? mem[148] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] :
                        (N0)? mem[147] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] :
                        (N0)? mem[146] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] :
                        (N0)? mem[145] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] :
                        (N0)? mem[144] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] :
                        (N0)? mem[143] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] :
                        (N0)? mem[142] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] :
                        (N0)? mem[141] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] :
                        (N0)? mem[140] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] :
                        (N0)? mem[139] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] :
                        (N0)? mem[138] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] :
                        (N0)? mem[137] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] :
                        (N0)? mem[136] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] :
                        (N0)? mem[135] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] :
                        (N0)? mem[134] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] :
                        (N0)? mem[133] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] :
                        (N0)? mem[132] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] :
                        (N0)? mem[131] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] :
                        (N0)? mem[130] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] :
                        (N0)? mem[129] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] :
                        (N0)? mem[128] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] :
                        (N0)? mem[127] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] :
                        (N0)? mem[126] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] :
                        (N0)? mem[125] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] :
                        (N0)? mem[124] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] :
                        (N0)? mem[123] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] :
                        (N0)? mem[122] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] :
                        (N0)? mem[121] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] :
                        (N0)? mem[120] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] :
                        (N0)? mem[119] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] :
                        (N0)? mem[118] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] :
                        (N0)? mem[117] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] :
                        (N0)? mem[116] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] :
                        (N0)? mem[115] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] :
                        (N0)? mem[114] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] :
                        (N0)? mem[113] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] :
                        (N0)? mem[112] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] :
                        (N0)? mem[111] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] :
                        (N0)? mem[110] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] :
                        (N0)? mem[109] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] :
                        (N0)? mem[108] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] :
                        (N0)? mem[107] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] :
                       (N0)? mem[106] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] :
                       (N0)? mem[105] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] :
                       (N0)? mem[104] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] :
                       (N0)? mem[103] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] :
                       (N0)? mem[102] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] :
                       (N0)? mem[101] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] :
                       (N0)? mem[100] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] :
                       (N0)? mem[99] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] :
                       (N0)? mem[98] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] :
                       (N0)? mem[97] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } :
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      { mem[193:97] } <= { w_data_i[96:0] };
    end
    if(N7) begin
      { mem[96:0] } <= { w_data_i[96:0] };
    end
  end


endmodule



module bsg_mem_1r1w_width_p97_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [96:0] w_data_i;
  input [0:0] r_addr_i;
  output [96:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [96:0] r_data_o;

  bsg_mem_p97
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p97
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [96:0] data_i;
  output [96:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [96:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p97_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 :
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 :
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 :
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 :
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 :
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 :
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end
    if(N9) begin
      tail_r <= N10;
    end
    if(N11) begin
      head_r <= N12;
    end
  end


endmodule



module bsg_mem_p26
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [25:0] w_data_i;
  input [0:0] r_addr_i;
  output [25:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [25:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  reg [51:0] mem;
  assign r_data_o[25] = (N3)? mem[25] :
                        (N0)? mem[51] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[24] = (N3)? mem[24] :
                        (N0)? mem[50] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] :
                        (N0)? mem[49] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] :
                        (N0)? mem[48] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] :
                        (N0)? mem[47] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] :
                        (N0)? mem[46] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] :
                        (N0)? mem[45] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] :
                        (N0)? mem[44] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] :
                        (N0)? mem[43] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] :
                        (N0)? mem[42] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] :
                        (N0)? mem[41] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] :
                        (N0)? mem[40] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] :
                        (N0)? mem[39] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] :
                        (N0)? mem[38] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] :
                        (N0)? mem[37] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] :
                        (N0)? mem[36] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] :
                       (N0)? mem[35] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] :
                       (N0)? mem[34] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] :
                       (N0)? mem[33] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] :
                       (N0)? mem[32] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] :
                       (N0)? mem[31] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] :
                       (N0)? mem[30] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] :
                       (N0)? mem[29] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] :
                       (N0)? mem[28] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] :
                       (N0)? mem[27] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] :
                       (N0)? mem[26] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } :
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      { mem[51:26] } <= { w_data_i[25:0] };
    end
    if(N7) begin
      { mem[25:0] } <= { w_data_i[25:0] };
    end
  end


endmodule



module bsg_mem_1r1w_width_p26_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [25:0] w_data_i;
  input [0:0] r_addr_i;
  output [25:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [25:0] r_data_o;

  bsg_mem_p26
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p26
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [25:0] data_i;
  output [25:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [25:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p26_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 :
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 :
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 :
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 :
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 :
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 :
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end
    if(N9) begin
      tail_r <= N10;
    end
    if(N11) begin
      head_r <= N12;
    end
  end


endmodule



module bsg_mem_p537
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [536:0] w_data_i;
  input [0:0] r_addr_i;
  output [536:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [536:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;
  reg [1073:0] mem;
  assign r_data_o[536] = (N3)? mem[536] :
                         (N0)? mem[1073] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[535] = (N3)? mem[535] :
                         (N0)? mem[1072] : 1'b0;
  assign r_data_o[534] = (N3)? mem[534] :
                         (N0)? mem[1071] : 1'b0;
  assign r_data_o[533] = (N3)? mem[533] :
                         (N0)? mem[1070] : 1'b0;
  assign r_data_o[532] = (N3)? mem[532] :
                         (N0)? mem[1069] : 1'b0;
  assign r_data_o[531] = (N3)? mem[531] :
                         (N0)? mem[1068] : 1'b0;
  assign r_data_o[530] = (N3)? mem[530] :
                         (N0)? mem[1067] : 1'b0;
  assign r_data_o[529] = (N3)? mem[529] :
                         (N0)? mem[1066] : 1'b0;
  assign r_data_o[528] = (N3)? mem[528] :
                         (N0)? mem[1065] : 1'b0;
  assign r_data_o[527] = (N3)? mem[527] :
                         (N0)? mem[1064] : 1'b0;
  assign r_data_o[526] = (N3)? mem[526] :
                         (N0)? mem[1063] : 1'b0;
  assign r_data_o[525] = (N3)? mem[525] :
                         (N0)? mem[1062] : 1'b0;
  assign r_data_o[524] = (N3)? mem[524] :
                         (N0)? mem[1061] : 1'b0;
  assign r_data_o[523] = (N3)? mem[523] :
                         (N0)? mem[1060] : 1'b0;
  assign r_data_o[522] = (N3)? mem[522] :
                         (N0)? mem[1059] : 1'b0;
  assign r_data_o[521] = (N3)? mem[521] :
                         (N0)? mem[1058] : 1'b0;
  assign r_data_o[520] = (N3)? mem[520] :
                         (N0)? mem[1057] : 1'b0;
  assign r_data_o[519] = (N3)? mem[519] :
                         (N0)? mem[1056] : 1'b0;
  assign r_data_o[518] = (N3)? mem[518] :
                         (N0)? mem[1055] : 1'b0;
  assign r_data_o[517] = (N3)? mem[517] :
                         (N0)? mem[1054] : 1'b0;
  assign r_data_o[516] = (N3)? mem[516] :
                         (N0)? mem[1053] : 1'b0;
  assign r_data_o[515] = (N3)? mem[515] :
                         (N0)? mem[1052] : 1'b0;
  assign r_data_o[514] = (N3)? mem[514] :
                         (N0)? mem[1051] : 1'b0;
  assign r_data_o[513] = (N3)? mem[513] :
                         (N0)? mem[1050] : 1'b0;
  assign r_data_o[512] = (N3)? mem[512] :
                         (N0)? mem[1049] : 1'b0;
  assign r_data_o[511] = (N3)? mem[511] :
                         (N0)? mem[1048] : 1'b0;
  assign r_data_o[510] = (N3)? mem[510] :
                         (N0)? mem[1047] : 1'b0;
  assign r_data_o[509] = (N3)? mem[509] :
                         (N0)? mem[1046] : 1'b0;
  assign r_data_o[508] = (N3)? mem[508] :
                         (N0)? mem[1045] : 1'b0;
  assign r_data_o[507] = (N3)? mem[507] :
                         (N0)? mem[1044] : 1'b0;
  assign r_data_o[506] = (N3)? mem[506] :
                         (N0)? mem[1043] : 1'b0;
  assign r_data_o[505] = (N3)? mem[505] :
                         (N0)? mem[1042] : 1'b0;
  assign r_data_o[504] = (N3)? mem[504] :
                         (N0)? mem[1041] : 1'b0;
  assign r_data_o[503] = (N3)? mem[503] :
                         (N0)? mem[1040] : 1'b0;
  assign r_data_o[502] = (N3)? mem[502] :
                         (N0)? mem[1039] : 1'b0;
  assign r_data_o[501] = (N3)? mem[501] :
                         (N0)? mem[1038] : 1'b0;
  assign r_data_o[500] = (N3)? mem[500] :
                         (N0)? mem[1037] : 1'b0;
  assign r_data_o[499] = (N3)? mem[499] :
                         (N0)? mem[1036] : 1'b0;
  assign r_data_o[498] = (N3)? mem[498] :
                         (N0)? mem[1035] : 1'b0;
  assign r_data_o[497] = (N3)? mem[497] :
                         (N0)? mem[1034] : 1'b0;
  assign r_data_o[496] = (N3)? mem[496] :
                         (N0)? mem[1033] : 1'b0;
  assign r_data_o[495] = (N3)? mem[495] :
                         (N0)? mem[1032] : 1'b0;
  assign r_data_o[494] = (N3)? mem[494] :
                         (N0)? mem[1031] : 1'b0;
  assign r_data_o[493] = (N3)? mem[493] :
                         (N0)? mem[1030] : 1'b0;
  assign r_data_o[492] = (N3)? mem[492] :
                         (N0)? mem[1029] : 1'b0;
  assign r_data_o[491] = (N3)? mem[491] :
                         (N0)? mem[1028] : 1'b0;
  assign r_data_o[490] = (N3)? mem[490] :
                         (N0)? mem[1027] : 1'b0;
  assign r_data_o[489] = (N3)? mem[489] :
                         (N0)? mem[1026] : 1'b0;
  assign r_data_o[488] = (N3)? mem[488] :
                         (N0)? mem[1025] : 1'b0;
  assign r_data_o[487] = (N3)? mem[487] :
                         (N0)? mem[1024] : 1'b0;
  assign r_data_o[486] = (N3)? mem[486] :
                         (N0)? mem[1023] : 1'b0;
  assign r_data_o[485] = (N3)? mem[485] :
                         (N0)? mem[1022] : 1'b0;
  assign r_data_o[484] = (N3)? mem[484] :
                         (N0)? mem[1021] : 1'b0;
  assign r_data_o[483] = (N3)? mem[483] :
                         (N0)? mem[1020] : 1'b0;
  assign r_data_o[482] = (N3)? mem[482] :
                         (N0)? mem[1019] : 1'b0;
  assign r_data_o[481] = (N3)? mem[481] :
                         (N0)? mem[1018] : 1'b0;
  assign r_data_o[480] = (N3)? mem[480] :
                         (N0)? mem[1017] : 1'b0;
  assign r_data_o[479] = (N3)? mem[479] :
                         (N0)? mem[1016] : 1'b0;
  assign r_data_o[478] = (N3)? mem[478] :
                         (N0)? mem[1015] : 1'b0;
  assign r_data_o[477] = (N3)? mem[477] :
                         (N0)? mem[1014] : 1'b0;
  assign r_data_o[476] = (N3)? mem[476] :
                         (N0)? mem[1013] : 1'b0;
  assign r_data_o[475] = (N3)? mem[475] :
                         (N0)? mem[1012] : 1'b0;
  assign r_data_o[474] = (N3)? mem[474] :
                         (N0)? mem[1011] : 1'b0;
  assign r_data_o[473] = (N3)? mem[473] :
                         (N0)? mem[1010] : 1'b0;
  assign r_data_o[472] = (N3)? mem[472] :
                         (N0)? mem[1009] : 1'b0;
  assign r_data_o[471] = (N3)? mem[471] :
                         (N0)? mem[1008] : 1'b0;
  assign r_data_o[470] = (N3)? mem[470] :
                         (N0)? mem[1007] : 1'b0;
  assign r_data_o[469] = (N3)? mem[469] :
                         (N0)? mem[1006] : 1'b0;
  assign r_data_o[468] = (N3)? mem[468] :
                         (N0)? mem[1005] : 1'b0;
  assign r_data_o[467] = (N3)? mem[467] :
                         (N0)? mem[1004] : 1'b0;
  assign r_data_o[466] = (N3)? mem[466] :
                         (N0)? mem[1003] : 1'b0;
  assign r_data_o[465] = (N3)? mem[465] :
                         (N0)? mem[1002] : 1'b0;
  assign r_data_o[464] = (N3)? mem[464] :
                         (N0)? mem[1001] : 1'b0;
  assign r_data_o[463] = (N3)? mem[463] :
                         (N0)? mem[1000] : 1'b0;
  assign r_data_o[462] = (N3)? mem[462] :
                         (N0)? mem[999] : 1'b0;
  assign r_data_o[461] = (N3)? mem[461] :
                         (N0)? mem[998] : 1'b0;
  assign r_data_o[460] = (N3)? mem[460] :
                         (N0)? mem[997] : 1'b0;
  assign r_data_o[459] = (N3)? mem[459] :
                         (N0)? mem[996] : 1'b0;
  assign r_data_o[458] = (N3)? mem[458] :
                         (N0)? mem[995] : 1'b0;
  assign r_data_o[457] = (N3)? mem[457] :
                         (N0)? mem[994] : 1'b0;
  assign r_data_o[456] = (N3)? mem[456] :
                         (N0)? mem[993] : 1'b0;
  assign r_data_o[455] = (N3)? mem[455] :
                         (N0)? mem[992] : 1'b0;
  assign r_data_o[454] = (N3)? mem[454] :
                         (N0)? mem[991] : 1'b0;
  assign r_data_o[453] = (N3)? mem[453] :
                         (N0)? mem[990] : 1'b0;
  assign r_data_o[452] = (N3)? mem[452] :
                         (N0)? mem[989] : 1'b0;
  assign r_data_o[451] = (N3)? mem[451] :
                         (N0)? mem[988] : 1'b0;
  assign r_data_o[450] = (N3)? mem[450] :
                         (N0)? mem[987] : 1'b0;
  assign r_data_o[449] = (N3)? mem[449] :
                         (N0)? mem[986] : 1'b0;
  assign r_data_o[448] = (N3)? mem[448] :
                         (N0)? mem[985] : 1'b0;
  assign r_data_o[447] = (N3)? mem[447] :
                         (N0)? mem[984] : 1'b0;
  assign r_data_o[446] = (N3)? mem[446] :
                         (N0)? mem[983] : 1'b0;
  assign r_data_o[445] = (N3)? mem[445] :
                         (N0)? mem[982] : 1'b0;
  assign r_data_o[444] = (N3)? mem[444] :
                         (N0)? mem[981] : 1'b0;
  assign r_data_o[443] = (N3)? mem[443] :
                         (N0)? mem[980] : 1'b0;
  assign r_data_o[442] = (N3)? mem[442] :
                         (N0)? mem[979] : 1'b0;
  assign r_data_o[441] = (N3)? mem[441] :
                         (N0)? mem[978] : 1'b0;
  assign r_data_o[440] = (N3)? mem[440] :
                         (N0)? mem[977] : 1'b0;
  assign r_data_o[439] = (N3)? mem[439] :
                         (N0)? mem[976] : 1'b0;
  assign r_data_o[438] = (N3)? mem[438] :
                         (N0)? mem[975] : 1'b0;
  assign r_data_o[437] = (N3)? mem[437] :
                         (N0)? mem[974] : 1'b0;
  assign r_data_o[436] = (N3)? mem[436] :
                         (N0)? mem[973] : 1'b0;
  assign r_data_o[435] = (N3)? mem[435] :
                         (N0)? mem[972] : 1'b0;
  assign r_data_o[434] = (N3)? mem[434] :
                         (N0)? mem[971] : 1'b0;
  assign r_data_o[433] = (N3)? mem[433] :
                         (N0)? mem[970] : 1'b0;
  assign r_data_o[432] = (N3)? mem[432] :
                         (N0)? mem[969] : 1'b0;
  assign r_data_o[431] = (N3)? mem[431] :
                         (N0)? mem[968] : 1'b0;
  assign r_data_o[430] = (N3)? mem[430] :
                         (N0)? mem[967] : 1'b0;
  assign r_data_o[429] = (N3)? mem[429] :
                         (N0)? mem[966] : 1'b0;
  assign r_data_o[428] = (N3)? mem[428] :
                         (N0)? mem[965] : 1'b0;
  assign r_data_o[427] = (N3)? mem[427] :
                         (N0)? mem[964] : 1'b0;
  assign r_data_o[426] = (N3)? mem[426] :
                         (N0)? mem[963] : 1'b0;
  assign r_data_o[425] = (N3)? mem[425] :
                         (N0)? mem[962] : 1'b0;
  assign r_data_o[424] = (N3)? mem[424] :
                         (N0)? mem[961] : 1'b0;
  assign r_data_o[423] = (N3)? mem[423] :
                         (N0)? mem[960] : 1'b0;
  assign r_data_o[422] = (N3)? mem[422] :
                         (N0)? mem[959] : 1'b0;
  assign r_data_o[421] = (N3)? mem[421] :
                         (N0)? mem[958] : 1'b0;
  assign r_data_o[420] = (N3)? mem[420] :
                         (N0)? mem[957] : 1'b0;
  assign r_data_o[419] = (N3)? mem[419] :
                         (N0)? mem[956] : 1'b0;
  assign r_data_o[418] = (N3)? mem[418] :
                         (N0)? mem[955] : 1'b0;
  assign r_data_o[417] = (N3)? mem[417] :
                         (N0)? mem[954] : 1'b0;
  assign r_data_o[416] = (N3)? mem[416] :
                         (N0)? mem[953] : 1'b0;
  assign r_data_o[415] = (N3)? mem[415] :
                         (N0)? mem[952] : 1'b0;
  assign r_data_o[414] = (N3)? mem[414] :
                         (N0)? mem[951] : 1'b0;
  assign r_data_o[413] = (N3)? mem[413] :
                         (N0)? mem[950] : 1'b0;
  assign r_data_o[412] = (N3)? mem[412] :
                         (N0)? mem[949] : 1'b0;
  assign r_data_o[411] = (N3)? mem[411] :
                         (N0)? mem[948] : 1'b0;
  assign r_data_o[410] = (N3)? mem[410] :
                         (N0)? mem[947] : 1'b0;
  assign r_data_o[409] = (N3)? mem[409] :
                         (N0)? mem[946] : 1'b0;
  assign r_data_o[408] = (N3)? mem[408] :
                         (N0)? mem[945] : 1'b0;
  assign r_data_o[407] = (N3)? mem[407] :
                         (N0)? mem[944] : 1'b0;
  assign r_data_o[406] = (N3)? mem[406] :
                         (N0)? mem[943] : 1'b0;
  assign r_data_o[405] = (N3)? mem[405] :
                         (N0)? mem[942] : 1'b0;
  assign r_data_o[404] = (N3)? mem[404] :
                         (N0)? mem[941] : 1'b0;
  assign r_data_o[403] = (N3)? mem[403] :
                         (N0)? mem[940] : 1'b0;
  assign r_data_o[402] = (N3)? mem[402] :
                         (N0)? mem[939] : 1'b0;
  assign r_data_o[401] = (N3)? mem[401] :
                         (N0)? mem[938] : 1'b0;
  assign r_data_o[400] = (N3)? mem[400] :
                         (N0)? mem[937] : 1'b0;
  assign r_data_o[399] = (N3)? mem[399] :
                         (N0)? mem[936] : 1'b0;
  assign r_data_o[398] = (N3)? mem[398] :
                         (N0)? mem[935] : 1'b0;
  assign r_data_o[397] = (N3)? mem[397] :
                         (N0)? mem[934] : 1'b0;
  assign r_data_o[396] = (N3)? mem[396] :
                         (N0)? mem[933] : 1'b0;
  assign r_data_o[395] = (N3)? mem[395] :
                         (N0)? mem[932] : 1'b0;
  assign r_data_o[394] = (N3)? mem[394] :
                         (N0)? mem[931] : 1'b0;
  assign r_data_o[393] = (N3)? mem[393] :
                         (N0)? mem[930] : 1'b0;
  assign r_data_o[392] = (N3)? mem[392] :
                         (N0)? mem[929] : 1'b0;
  assign r_data_o[391] = (N3)? mem[391] :
                         (N0)? mem[928] : 1'b0;
  assign r_data_o[390] = (N3)? mem[390] :
                         (N0)? mem[927] : 1'b0;
  assign r_data_o[389] = (N3)? mem[389] :
                         (N0)? mem[926] : 1'b0;
  assign r_data_o[388] = (N3)? mem[388] :
                         (N0)? mem[925] : 1'b0;
  assign r_data_o[387] = (N3)? mem[387] :
                         (N0)? mem[924] : 1'b0;
  assign r_data_o[386] = (N3)? mem[386] :
                         (N0)? mem[923] : 1'b0;
  assign r_data_o[385] = (N3)? mem[385] :
                         (N0)? mem[922] : 1'b0;
  assign r_data_o[384] = (N3)? mem[384] :
                         (N0)? mem[921] : 1'b0;
  assign r_data_o[383] = (N3)? mem[383] :
                         (N0)? mem[920] : 1'b0;
  assign r_data_o[382] = (N3)? mem[382] :
                         (N0)? mem[919] : 1'b0;
  assign r_data_o[381] = (N3)? mem[381] :
                         (N0)? mem[918] : 1'b0;
  assign r_data_o[380] = (N3)? mem[380] :
                         (N0)? mem[917] : 1'b0;
  assign r_data_o[379] = (N3)? mem[379] :
                         (N0)? mem[916] : 1'b0;
  assign r_data_o[378] = (N3)? mem[378] :
                         (N0)? mem[915] : 1'b0;
  assign r_data_o[377] = (N3)? mem[377] :
                         (N0)? mem[914] : 1'b0;
  assign r_data_o[376] = (N3)? mem[376] :
                         (N0)? mem[913] : 1'b0;
  assign r_data_o[375] = (N3)? mem[375] :
                         (N0)? mem[912] : 1'b0;
  assign r_data_o[374] = (N3)? mem[374] :
                         (N0)? mem[911] : 1'b0;
  assign r_data_o[373] = (N3)? mem[373] :
                         (N0)? mem[910] : 1'b0;
  assign r_data_o[372] = (N3)? mem[372] :
                         (N0)? mem[909] : 1'b0;
  assign r_data_o[371] = (N3)? mem[371] :
                         (N0)? mem[908] : 1'b0;
  assign r_data_o[370] = (N3)? mem[370] :
                         (N0)? mem[907] : 1'b0;
  assign r_data_o[369] = (N3)? mem[369] :
                         (N0)? mem[906] : 1'b0;
  assign r_data_o[368] = (N3)? mem[368] :
                         (N0)? mem[905] : 1'b0;
  assign r_data_o[367] = (N3)? mem[367] :
                         (N0)? mem[904] : 1'b0;
  assign r_data_o[366] = (N3)? mem[366] :
                         (N0)? mem[903] : 1'b0;
  assign r_data_o[365] = (N3)? mem[365] :
                         (N0)? mem[902] : 1'b0;
  assign r_data_o[364] = (N3)? mem[364] :
                         (N0)? mem[901] : 1'b0;
  assign r_data_o[363] = (N3)? mem[363] :
                         (N0)? mem[900] : 1'b0;
  assign r_data_o[362] = (N3)? mem[362] :
                         (N0)? mem[899] : 1'b0;
  assign r_data_o[361] = (N3)? mem[361] :
                         (N0)? mem[898] : 1'b0;
  assign r_data_o[360] = (N3)? mem[360] :
                         (N0)? mem[897] : 1'b0;
  assign r_data_o[359] = (N3)? mem[359] :
                         (N0)? mem[896] : 1'b0;
  assign r_data_o[358] = (N3)? mem[358] :
                         (N0)? mem[895] : 1'b0;
  assign r_data_o[357] = (N3)? mem[357] :
                         (N0)? mem[894] : 1'b0;
  assign r_data_o[356] = (N3)? mem[356] :
                         (N0)? mem[893] : 1'b0;
  assign r_data_o[355] = (N3)? mem[355] :
                         (N0)? mem[892] : 1'b0;
  assign r_data_o[354] = (N3)? mem[354] :
                         (N0)? mem[891] : 1'b0;
  assign r_data_o[353] = (N3)? mem[353] :
                         (N0)? mem[890] : 1'b0;
  assign r_data_o[352] = (N3)? mem[352] :
                         (N0)? mem[889] : 1'b0;
  assign r_data_o[351] = (N3)? mem[351] :
                         (N0)? mem[888] : 1'b0;
  assign r_data_o[350] = (N3)? mem[350] :
                         (N0)? mem[887] : 1'b0;
  assign r_data_o[349] = (N3)? mem[349] :
                         (N0)? mem[886] : 1'b0;
  assign r_data_o[348] = (N3)? mem[348] :
                         (N0)? mem[885] : 1'b0;
  assign r_data_o[347] = (N3)? mem[347] :
                         (N0)? mem[884] : 1'b0;
  assign r_data_o[346] = (N3)? mem[346] :
                         (N0)? mem[883] : 1'b0;
  assign r_data_o[345] = (N3)? mem[345] :
                         (N0)? mem[882] : 1'b0;
  assign r_data_o[344] = (N3)? mem[344] :
                         (N0)? mem[881] : 1'b0;
  assign r_data_o[343] = (N3)? mem[343] :
                         (N0)? mem[880] : 1'b0;
  assign r_data_o[342] = (N3)? mem[342] :
                         (N0)? mem[879] : 1'b0;
  assign r_data_o[341] = (N3)? mem[341] :
                         (N0)? mem[878] : 1'b0;
  assign r_data_o[340] = (N3)? mem[340] :
                         (N0)? mem[877] : 1'b0;
  assign r_data_o[339] = (N3)? mem[339] :
                         (N0)? mem[876] : 1'b0;
  assign r_data_o[338] = (N3)? mem[338] :
                         (N0)? mem[875] : 1'b0;
  assign r_data_o[337] = (N3)? mem[337] :
                         (N0)? mem[874] : 1'b0;
  assign r_data_o[336] = (N3)? mem[336] :
                         (N0)? mem[873] : 1'b0;
  assign r_data_o[335] = (N3)? mem[335] :
                         (N0)? mem[872] : 1'b0;
  assign r_data_o[334] = (N3)? mem[334] :
                         (N0)? mem[871] : 1'b0;
  assign r_data_o[333] = (N3)? mem[333] :
                         (N0)? mem[870] : 1'b0;
  assign r_data_o[332] = (N3)? mem[332] :
                         (N0)? mem[869] : 1'b0;
  assign r_data_o[331] = (N3)? mem[331] :
                         (N0)? mem[868] : 1'b0;
  assign r_data_o[330] = (N3)? mem[330] :
                         (N0)? mem[867] : 1'b0;
  assign r_data_o[329] = (N3)? mem[329] :
                         (N0)? mem[866] : 1'b0;
  assign r_data_o[328] = (N3)? mem[328] :
                         (N0)? mem[865] : 1'b0;
  assign r_data_o[327] = (N3)? mem[327] :
                         (N0)? mem[864] : 1'b0;
  assign r_data_o[326] = (N3)? mem[326] :
                         (N0)? mem[863] : 1'b0;
  assign r_data_o[325] = (N3)? mem[325] :
                         (N0)? mem[862] : 1'b0;
  assign r_data_o[324] = (N3)? mem[324] :
                         (N0)? mem[861] : 1'b0;
  assign r_data_o[323] = (N3)? mem[323] :
                         (N0)? mem[860] : 1'b0;
  assign r_data_o[322] = (N3)? mem[322] :
                         (N0)? mem[859] : 1'b0;
  assign r_data_o[321] = (N3)? mem[321] :
                         (N0)? mem[858] : 1'b0;
  assign r_data_o[320] = (N3)? mem[320] :
                         (N0)? mem[857] : 1'b0;
  assign r_data_o[319] = (N3)? mem[319] :
                         (N0)? mem[856] : 1'b0;
  assign r_data_o[318] = (N3)? mem[318] :
                         (N0)? mem[855] : 1'b0;
  assign r_data_o[317] = (N3)? mem[317] :
                         (N0)? mem[854] : 1'b0;
  assign r_data_o[316] = (N3)? mem[316] :
                         (N0)? mem[853] : 1'b0;
  assign r_data_o[315] = (N3)? mem[315] :
                         (N0)? mem[852] : 1'b0;
  assign r_data_o[314] = (N3)? mem[314] :
                         (N0)? mem[851] : 1'b0;
  assign r_data_o[313] = (N3)? mem[313] :
                         (N0)? mem[850] : 1'b0;
  assign r_data_o[312] = (N3)? mem[312] :
                         (N0)? mem[849] : 1'b0;
  assign r_data_o[311] = (N3)? mem[311] :
                         (N0)? mem[848] : 1'b0;
  assign r_data_o[310] = (N3)? mem[310] :
                         (N0)? mem[847] : 1'b0;
  assign r_data_o[309] = (N3)? mem[309] :
                         (N0)? mem[846] : 1'b0;
  assign r_data_o[308] = (N3)? mem[308] :
                         (N0)? mem[845] : 1'b0;
  assign r_data_o[307] = (N3)? mem[307] :
                         (N0)? mem[844] : 1'b0;
  assign r_data_o[306] = (N3)? mem[306] :
                         (N0)? mem[843] : 1'b0;
  assign r_data_o[305] = (N3)? mem[305] :
                         (N0)? mem[842] : 1'b0;
  assign r_data_o[304] = (N3)? mem[304] :
                         (N0)? mem[841] : 1'b0;
  assign r_data_o[303] = (N3)? mem[303] :
                         (N0)? mem[840] : 1'b0;
  assign r_data_o[302] = (N3)? mem[302] :
                         (N0)? mem[839] : 1'b0;
  assign r_data_o[301] = (N3)? mem[301] :
                         (N0)? mem[838] : 1'b0;
  assign r_data_o[300] = (N3)? mem[300] :
                         (N0)? mem[837] : 1'b0;
  assign r_data_o[299] = (N3)? mem[299] :
                         (N0)? mem[836] : 1'b0;
  assign r_data_o[298] = (N3)? mem[298] :
                         (N0)? mem[835] : 1'b0;
  assign r_data_o[297] = (N3)? mem[297] :
                         (N0)? mem[834] : 1'b0;
  assign r_data_o[296] = (N3)? mem[296] :
                         (N0)? mem[833] : 1'b0;
  assign r_data_o[295] = (N3)? mem[295] :
                         (N0)? mem[832] : 1'b0;
  assign r_data_o[294] = (N3)? mem[294] :
                         (N0)? mem[831] : 1'b0;
  assign r_data_o[293] = (N3)? mem[293] :
                         (N0)? mem[830] : 1'b0;
  assign r_data_o[292] = (N3)? mem[292] :
                         (N0)? mem[829] : 1'b0;
  assign r_data_o[291] = (N3)? mem[291] :
                         (N0)? mem[828] : 1'b0;
  assign r_data_o[290] = (N3)? mem[290] :
                         (N0)? mem[827] : 1'b0;
  assign r_data_o[289] = (N3)? mem[289] :
                         (N0)? mem[826] : 1'b0;
  assign r_data_o[288] = (N3)? mem[288] :
                         (N0)? mem[825] : 1'b0;
  assign r_data_o[287] = (N3)? mem[287] :
                         (N0)? mem[824] : 1'b0;
  assign r_data_o[286] = (N3)? mem[286] :
                         (N0)? mem[823] : 1'b0;
  assign r_data_o[285] = (N3)? mem[285] :
                         (N0)? mem[822] : 1'b0;
  assign r_data_o[284] = (N3)? mem[284] :
                         (N0)? mem[821] : 1'b0;
  assign r_data_o[283] = (N3)? mem[283] :
                         (N0)? mem[820] : 1'b0;
  assign r_data_o[282] = (N3)? mem[282] :
                         (N0)? mem[819] : 1'b0;
  assign r_data_o[281] = (N3)? mem[281] :
                         (N0)? mem[818] : 1'b0;
  assign r_data_o[280] = (N3)? mem[280] :
                         (N0)? mem[817] : 1'b0;
  assign r_data_o[279] = (N3)? mem[279] :
                         (N0)? mem[816] : 1'b0;
  assign r_data_o[278] = (N3)? mem[278] :
                         (N0)? mem[815] : 1'b0;
  assign r_data_o[277] = (N3)? mem[277] :
                         (N0)? mem[814] : 1'b0;
  assign r_data_o[276] = (N3)? mem[276] :
                         (N0)? mem[813] : 1'b0;
  assign r_data_o[275] = (N3)? mem[275] :
                         (N0)? mem[812] : 1'b0;
  assign r_data_o[274] = (N3)? mem[274] :
                         (N0)? mem[811] : 1'b0;
  assign r_data_o[273] = (N3)? mem[273] :
                         (N0)? mem[810] : 1'b0;
  assign r_data_o[272] = (N3)? mem[272] :
                         (N0)? mem[809] : 1'b0;
  assign r_data_o[271] = (N3)? mem[271] :
                         (N0)? mem[808] : 1'b0;
  assign r_data_o[270] = (N3)? mem[270] :
                         (N0)? mem[807] : 1'b0;
  assign r_data_o[269] = (N3)? mem[269] :
                         (N0)? mem[806] : 1'b0;
  assign r_data_o[268] = (N3)? mem[268] :
                         (N0)? mem[805] : 1'b0;
  assign r_data_o[267] = (N3)? mem[267] :
                         (N0)? mem[804] : 1'b0;
  assign r_data_o[266] = (N3)? mem[266] :
                         (N0)? mem[803] : 1'b0;
  assign r_data_o[265] = (N3)? mem[265] :
                         (N0)? mem[802] : 1'b0;
  assign r_data_o[264] = (N3)? mem[264] :
                         (N0)? mem[801] : 1'b0;
  assign r_data_o[263] = (N3)? mem[263] :
                         (N0)? mem[800] : 1'b0;
  assign r_data_o[262] = (N3)? mem[262] :
                         (N0)? mem[799] : 1'b0;
  assign r_data_o[261] = (N3)? mem[261] :
                         (N0)? mem[798] : 1'b0;
  assign r_data_o[260] = (N3)? mem[260] :
                         (N0)? mem[797] : 1'b0;
  assign r_data_o[259] = (N3)? mem[259] :
                         (N0)? mem[796] : 1'b0;
  assign r_data_o[258] = (N3)? mem[258] :
                         (N0)? mem[795] : 1'b0;
  assign r_data_o[257] = (N3)? mem[257] :
                         (N0)? mem[794] : 1'b0;
  assign r_data_o[256] = (N3)? mem[256] :
                         (N0)? mem[793] : 1'b0;
  assign r_data_o[255] = (N3)? mem[255] :
                         (N0)? mem[792] : 1'b0;
  assign r_data_o[254] = (N3)? mem[254] :
                         (N0)? mem[791] : 1'b0;
  assign r_data_o[253] = (N3)? mem[253] :
                         (N0)? mem[790] : 1'b0;
  assign r_data_o[252] = (N3)? mem[252] :
                         (N0)? mem[789] : 1'b0;
  assign r_data_o[251] = (N3)? mem[251] :
                         (N0)? mem[788] : 1'b0;
  assign r_data_o[250] = (N3)? mem[250] :
                         (N0)? mem[787] : 1'b0;
  assign r_data_o[249] = (N3)? mem[249] :
                         (N0)? mem[786] : 1'b0;
  assign r_data_o[248] = (N3)? mem[248] :
                         (N0)? mem[785] : 1'b0;
  assign r_data_o[247] = (N3)? mem[247] :
                         (N0)? mem[784] : 1'b0;
  assign r_data_o[246] = (N3)? mem[246] :
                         (N0)? mem[783] : 1'b0;
  assign r_data_o[245] = (N3)? mem[245] :
                         (N0)? mem[782] : 1'b0;
  assign r_data_o[244] = (N3)? mem[244] :
                         (N0)? mem[781] : 1'b0;
  assign r_data_o[243] = (N3)? mem[243] :
                         (N0)? mem[780] : 1'b0;
  assign r_data_o[242] = (N3)? mem[242] :
                         (N0)? mem[779] : 1'b0;
  assign r_data_o[241] = (N3)? mem[241] :
                         (N0)? mem[778] : 1'b0;
  assign r_data_o[240] = (N3)? mem[240] :
                         (N0)? mem[777] : 1'b0;
  assign r_data_o[239] = (N3)? mem[239] :
                         (N0)? mem[776] : 1'b0;
  assign r_data_o[238] = (N3)? mem[238] :
                         (N0)? mem[775] : 1'b0;
  assign r_data_o[237] = (N3)? mem[237] :
                         (N0)? mem[774] : 1'b0;
  assign r_data_o[236] = (N3)? mem[236] :
                         (N0)? mem[773] : 1'b0;
  assign r_data_o[235] = (N3)? mem[235] :
                         (N0)? mem[772] : 1'b0;
  assign r_data_o[234] = (N3)? mem[234] :
                         (N0)? mem[771] : 1'b0;
  assign r_data_o[233] = (N3)? mem[233] :
                         (N0)? mem[770] : 1'b0;
  assign r_data_o[232] = (N3)? mem[232] :
                         (N0)? mem[769] : 1'b0;
  assign r_data_o[231] = (N3)? mem[231] :
                         (N0)? mem[768] : 1'b0;
  assign r_data_o[230] = (N3)? mem[230] :
                         (N0)? mem[767] : 1'b0;
  assign r_data_o[229] = (N3)? mem[229] :
                         (N0)? mem[766] : 1'b0;
  assign r_data_o[228] = (N3)? mem[228] :
                         (N0)? mem[765] : 1'b0;
  assign r_data_o[227] = (N3)? mem[227] :
                         (N0)? mem[764] : 1'b0;
  assign r_data_o[226] = (N3)? mem[226] :
                         (N0)? mem[763] : 1'b0;
  assign r_data_o[225] = (N3)? mem[225] :
                         (N0)? mem[762] : 1'b0;
  assign r_data_o[224] = (N3)? mem[224] :
                         (N0)? mem[761] : 1'b0;
  assign r_data_o[223] = (N3)? mem[223] :
                         (N0)? mem[760] : 1'b0;
  assign r_data_o[222] = (N3)? mem[222] :
                         (N0)? mem[759] : 1'b0;
  assign r_data_o[221] = (N3)? mem[221] :
                         (N0)? mem[758] : 1'b0;
  assign r_data_o[220] = (N3)? mem[220] :
                         (N0)? mem[757] : 1'b0;
  assign r_data_o[219] = (N3)? mem[219] :
                         (N0)? mem[756] : 1'b0;
  assign r_data_o[218] = (N3)? mem[218] :
                         (N0)? mem[755] : 1'b0;
  assign r_data_o[217] = (N3)? mem[217] :
                         (N0)? mem[754] : 1'b0;
  assign r_data_o[216] = (N3)? mem[216] :
                         (N0)? mem[753] : 1'b0;
  assign r_data_o[215] = (N3)? mem[215] :
                         (N0)? mem[752] : 1'b0;
  assign r_data_o[214] = (N3)? mem[214] :
                         (N0)? mem[751] : 1'b0;
  assign r_data_o[213] = (N3)? mem[213] :
                         (N0)? mem[750] : 1'b0;
  assign r_data_o[212] = (N3)? mem[212] :
                         (N0)? mem[749] : 1'b0;
  assign r_data_o[211] = (N3)? mem[211] :
                         (N0)? mem[748] : 1'b0;
  assign r_data_o[210] = (N3)? mem[210] :
                         (N0)? mem[747] : 1'b0;
  assign r_data_o[209] = (N3)? mem[209] :
                         (N0)? mem[746] : 1'b0;
  assign r_data_o[208] = (N3)? mem[208] :
                         (N0)? mem[745] : 1'b0;
  assign r_data_o[207] = (N3)? mem[207] :
                         (N0)? mem[744] : 1'b0;
  assign r_data_o[206] = (N3)? mem[206] :
                         (N0)? mem[743] : 1'b0;
  assign r_data_o[205] = (N3)? mem[205] :
                         (N0)? mem[742] : 1'b0;
  assign r_data_o[204] = (N3)? mem[204] :
                         (N0)? mem[741] : 1'b0;
  assign r_data_o[203] = (N3)? mem[203] :
                         (N0)? mem[740] : 1'b0;
  assign r_data_o[202] = (N3)? mem[202] :
                         (N0)? mem[739] : 1'b0;
  assign r_data_o[201] = (N3)? mem[201] :
                         (N0)? mem[738] : 1'b0;
  assign r_data_o[200] = (N3)? mem[200] :
                         (N0)? mem[737] : 1'b0;
  assign r_data_o[199] = (N3)? mem[199] :
                         (N0)? mem[736] : 1'b0;
  assign r_data_o[198] = (N3)? mem[198] :
                         (N0)? mem[735] : 1'b0;
  assign r_data_o[197] = (N3)? mem[197] :
                         (N0)? mem[734] : 1'b0;
  assign r_data_o[196] = (N3)? mem[196] :
                         (N0)? mem[733] : 1'b0;
  assign r_data_o[195] = (N3)? mem[195] :
                         (N0)? mem[732] : 1'b0;
  assign r_data_o[194] = (N3)? mem[194] :
                         (N0)? mem[731] : 1'b0;
  assign r_data_o[193] = (N3)? mem[193] :
                         (N0)? mem[730] : 1'b0;
  assign r_data_o[192] = (N3)? mem[192] :
                         (N0)? mem[729] : 1'b0;
  assign r_data_o[191] = (N3)? mem[191] :
                         (N0)? mem[728] : 1'b0;
  assign r_data_o[190] = (N3)? mem[190] :
                         (N0)? mem[727] : 1'b0;
  assign r_data_o[189] = (N3)? mem[189] :
                         (N0)? mem[726] : 1'b0;
  assign r_data_o[188] = (N3)? mem[188] :
                         (N0)? mem[725] : 1'b0;
  assign r_data_o[187] = (N3)? mem[187] :
                         (N0)? mem[724] : 1'b0;
  assign r_data_o[186] = (N3)? mem[186] :
                         (N0)? mem[723] : 1'b0;
  assign r_data_o[185] = (N3)? mem[185] :
                         (N0)? mem[722] : 1'b0;
  assign r_data_o[184] = (N3)? mem[184] :
                         (N0)? mem[721] : 1'b0;
  assign r_data_o[183] = (N3)? mem[183] :
                         (N0)? mem[720] : 1'b0;
  assign r_data_o[182] = (N3)? mem[182] :
                         (N0)? mem[719] : 1'b0;
  assign r_data_o[181] = (N3)? mem[181] :
                         (N0)? mem[718] : 1'b0;
  assign r_data_o[180] = (N3)? mem[180] :
                         (N0)? mem[717] : 1'b0;
  assign r_data_o[179] = (N3)? mem[179] :
                         (N0)? mem[716] : 1'b0;
  assign r_data_o[178] = (N3)? mem[178] :
                         (N0)? mem[715] : 1'b0;
  assign r_data_o[177] = (N3)? mem[177] :
                         (N0)? mem[714] : 1'b0;
  assign r_data_o[176] = (N3)? mem[176] :
                         (N0)? mem[713] : 1'b0;
  assign r_data_o[175] = (N3)? mem[175] :
                         (N0)? mem[712] : 1'b0;
  assign r_data_o[174] = (N3)? mem[174] :
                         (N0)? mem[711] : 1'b0;
  assign r_data_o[173] = (N3)? mem[173] :
                         (N0)? mem[710] : 1'b0;
  assign r_data_o[172] = (N3)? mem[172] :
                         (N0)? mem[709] : 1'b0;
  assign r_data_o[171] = (N3)? mem[171] :
                         (N0)? mem[708] : 1'b0;
  assign r_data_o[170] = (N3)? mem[170] :
                         (N0)? mem[707] : 1'b0;
  assign r_data_o[169] = (N3)? mem[169] :
                         (N0)? mem[706] : 1'b0;
  assign r_data_o[168] = (N3)? mem[168] :
                         (N0)? mem[705] : 1'b0;
  assign r_data_o[167] = (N3)? mem[167] :
                         (N0)? mem[704] : 1'b0;
  assign r_data_o[166] = (N3)? mem[166] :
                         (N0)? mem[703] : 1'b0;
  assign r_data_o[165] = (N3)? mem[165] :
                         (N0)? mem[702] : 1'b0;
  assign r_data_o[164] = (N3)? mem[164] :
                         (N0)? mem[701] : 1'b0;
  assign r_data_o[163] = (N3)? mem[163] :
                         (N0)? mem[700] : 1'b0;
  assign r_data_o[162] = (N3)? mem[162] :
                         (N0)? mem[699] : 1'b0;
  assign r_data_o[161] = (N3)? mem[161] :
                         (N0)? mem[698] : 1'b0;
  assign r_data_o[160] = (N3)? mem[160] :
                         (N0)? mem[697] : 1'b0;
  assign r_data_o[159] = (N3)? mem[159] :
                         (N0)? mem[696] : 1'b0;
  assign r_data_o[158] = (N3)? mem[158] :
                         (N0)? mem[695] : 1'b0;
  assign r_data_o[157] = (N3)? mem[157] :
                         (N0)? mem[694] : 1'b0;
  assign r_data_o[156] = (N3)? mem[156] :
                         (N0)? mem[693] : 1'b0;
  assign r_data_o[155] = (N3)? mem[155] :
                         (N0)? mem[692] : 1'b0;
  assign r_data_o[154] = (N3)? mem[154] :
                         (N0)? mem[691] : 1'b0;
  assign r_data_o[153] = (N3)? mem[153] :
                         (N0)? mem[690] : 1'b0;
  assign r_data_o[152] = (N3)? mem[152] :
                         (N0)? mem[689] : 1'b0;
  assign r_data_o[151] = (N3)? mem[151] :
                         (N0)? mem[688] : 1'b0;
  assign r_data_o[150] = (N3)? mem[150] :
                         (N0)? mem[687] : 1'b0;
  assign r_data_o[149] = (N3)? mem[149] :
                         (N0)? mem[686] : 1'b0;
  assign r_data_o[148] = (N3)? mem[148] :
                         (N0)? mem[685] : 1'b0;
  assign r_data_o[147] = (N3)? mem[147] :
                         (N0)? mem[684] : 1'b0;
  assign r_data_o[146] = (N3)? mem[146] :
                         (N0)? mem[683] : 1'b0;
  assign r_data_o[145] = (N3)? mem[145] :
                         (N0)? mem[682] : 1'b0;
  assign r_data_o[144] = (N3)? mem[144] :
                         (N0)? mem[681] : 1'b0;
  assign r_data_o[143] = (N3)? mem[143] :
                         (N0)? mem[680] : 1'b0;
  assign r_data_o[142] = (N3)? mem[142] :
                         (N0)? mem[679] : 1'b0;
  assign r_data_o[141] = (N3)? mem[141] :
                         (N0)? mem[678] : 1'b0;
  assign r_data_o[140] = (N3)? mem[140] :
                         (N0)? mem[677] : 1'b0;
  assign r_data_o[139] = (N3)? mem[139] :
                         (N0)? mem[676] : 1'b0;
  assign r_data_o[138] = (N3)? mem[138] :
                         (N0)? mem[675] : 1'b0;
  assign r_data_o[137] = (N3)? mem[137] :
                         (N0)? mem[674] : 1'b0;
  assign r_data_o[136] = (N3)? mem[136] :
                         (N0)? mem[673] : 1'b0;
  assign r_data_o[135] = (N3)? mem[135] :
                         (N0)? mem[672] : 1'b0;
  assign r_data_o[134] = (N3)? mem[134] :
                         (N0)? mem[671] : 1'b0;
  assign r_data_o[133] = (N3)? mem[133] :
                         (N0)? mem[670] : 1'b0;
  assign r_data_o[132] = (N3)? mem[132] :
                         (N0)? mem[669] : 1'b0;
  assign r_data_o[131] = (N3)? mem[131] :
                         (N0)? mem[668] : 1'b0;
  assign r_data_o[130] = (N3)? mem[130] :
                         (N0)? mem[667] : 1'b0;
  assign r_data_o[129] = (N3)? mem[129] :
                         (N0)? mem[666] : 1'b0;
  assign r_data_o[128] = (N3)? mem[128] :
                         (N0)? mem[665] : 1'b0;
  assign r_data_o[127] = (N3)? mem[127] :
                         (N0)? mem[664] : 1'b0;
  assign r_data_o[126] = (N3)? mem[126] :
                         (N0)? mem[663] : 1'b0;
  assign r_data_o[125] = (N3)? mem[125] :
                         (N0)? mem[662] : 1'b0;
  assign r_data_o[124] = (N3)? mem[124] :
                         (N0)? mem[661] : 1'b0;
  assign r_data_o[123] = (N3)? mem[123] :
                         (N0)? mem[660] : 1'b0;
  assign r_data_o[122] = (N3)? mem[122] :
                         (N0)? mem[659] : 1'b0;
  assign r_data_o[121] = (N3)? mem[121] :
                         (N0)? mem[658] : 1'b0;
  assign r_data_o[120] = (N3)? mem[120] :
                         (N0)? mem[657] : 1'b0;
  assign r_data_o[119] = (N3)? mem[119] :
                         (N0)? mem[656] : 1'b0;
  assign r_data_o[118] = (N3)? mem[118] :
                         (N0)? mem[655] : 1'b0;
  assign r_data_o[117] = (N3)? mem[117] :
                         (N0)? mem[654] : 1'b0;
  assign r_data_o[116] = (N3)? mem[116] :
                         (N0)? mem[653] : 1'b0;
  assign r_data_o[115] = (N3)? mem[115] :
                         (N0)? mem[652] : 1'b0;
  assign r_data_o[114] = (N3)? mem[114] :
                         (N0)? mem[651] : 1'b0;
  assign r_data_o[113] = (N3)? mem[113] :
                         (N0)? mem[650] : 1'b0;
  assign r_data_o[112] = (N3)? mem[112] :
                         (N0)? mem[649] : 1'b0;
  assign r_data_o[111] = (N3)? mem[111] :
                         (N0)? mem[648] : 1'b0;
  assign r_data_o[110] = (N3)? mem[110] :
                         (N0)? mem[647] : 1'b0;
  assign r_data_o[109] = (N3)? mem[109] :
                         (N0)? mem[646] : 1'b0;
  assign r_data_o[108] = (N3)? mem[108] :
                         (N0)? mem[645] : 1'b0;
  assign r_data_o[107] = (N3)? mem[107] :
                         (N0)? mem[644] : 1'b0;
  assign r_data_o[106] = (N3)? mem[106] :
                         (N0)? mem[643] : 1'b0;
  assign r_data_o[105] = (N3)? mem[105] :
                         (N0)? mem[642] : 1'b0;
  assign r_data_o[104] = (N3)? mem[104] :
                         (N0)? mem[641] : 1'b0;
  assign r_data_o[103] = (N3)? mem[103] :
                         (N0)? mem[640] : 1'b0;
  assign r_data_o[102] = (N3)? mem[102] :
                         (N0)? mem[639] : 1'b0;
  assign r_data_o[101] = (N3)? mem[101] :
                         (N0)? mem[638] : 1'b0;
  assign r_data_o[100] = (N3)? mem[100] :
                         (N0)? mem[637] : 1'b0;
  assign r_data_o[99] = (N3)? mem[99] :
                        (N0)? mem[636] : 1'b0;
  assign r_data_o[98] = (N3)? mem[98] :
                        (N0)? mem[635] : 1'b0;
  assign r_data_o[97] = (N3)? mem[97] :
                        (N0)? mem[634] : 1'b0;
  assign r_data_o[96] = (N3)? mem[96] :
                        (N0)? mem[633] : 1'b0;
  assign r_data_o[95] = (N3)? mem[95] :
                        (N0)? mem[632] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] :
                        (N0)? mem[631] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] :
                        (N0)? mem[630] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] :
                        (N0)? mem[629] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] :
                        (N0)? mem[628] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] :
                        (N0)? mem[627] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] :
                        (N0)? mem[626] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] :
                        (N0)? mem[625] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] :
                        (N0)? mem[624] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] :
                        (N0)? mem[623] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] :
                        (N0)? mem[622] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] :
                        (N0)? mem[621] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] :
                        (N0)? mem[620] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] :
                        (N0)? mem[619] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] :
                        (N0)? mem[618] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] :
                        (N0)? mem[617] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] :
                        (N0)? mem[616] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] :
                        (N0)? mem[615] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] :
                        (N0)? mem[614] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] :
                        (N0)? mem[613] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] :
                        (N0)? mem[612] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] :
                        (N0)? mem[611] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] :
                        (N0)? mem[610] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] :
                        (N0)? mem[609] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] :
                        (N0)? mem[608] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] :
                        (N0)? mem[607] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] :
                        (N0)? mem[606] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] :
                        (N0)? mem[605] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] :
                        (N0)? mem[604] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] :
                        (N0)? mem[603] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] :
                        (N0)? mem[602] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] :
                        (N0)? mem[601] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] :
                        (N0)? mem[600] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] :
                        (N0)? mem[599] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] :
                        (N0)? mem[598] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] :
                        (N0)? mem[597] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] :
                        (N0)? mem[596] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] :
                        (N0)? mem[595] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] :
                        (N0)? mem[594] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] :
                        (N0)? mem[593] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] :
                        (N0)? mem[592] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] :
                        (N0)? mem[591] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] :
                        (N0)? mem[590] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] :
                        (N0)? mem[589] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] :
                        (N0)? mem[588] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] :
                        (N0)? mem[587] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] :
                        (N0)? mem[586] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] :
                        (N0)? mem[585] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] :
                        (N0)? mem[584] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] :
                        (N0)? mem[583] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] :
                        (N0)? mem[582] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] :
                        (N0)? mem[581] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] :
                        (N0)? mem[580] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] :
                        (N0)? mem[579] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] :
                        (N0)? mem[578] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] :
                        (N0)? mem[577] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] :
                        (N0)? mem[576] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] :
                        (N0)? mem[575] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] :
                        (N0)? mem[574] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] :
                        (N0)? mem[573] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] :
                        (N0)? mem[572] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] :
                        (N0)? mem[571] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] :
                        (N0)? mem[570] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] :
                        (N0)? mem[569] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] :
                        (N0)? mem[568] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] :
                        (N0)? mem[567] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] :
                        (N0)? mem[566] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] :
                        (N0)? mem[565] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] :
                        (N0)? mem[564] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] :
                        (N0)? mem[563] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] :
                        (N0)? mem[562] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] :
                        (N0)? mem[561] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] :
                        (N0)? mem[560] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] :
                        (N0)? mem[559] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] :
                        (N0)? mem[558] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] :
                        (N0)? mem[557] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] :
                        (N0)? mem[556] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] :
                        (N0)? mem[555] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] :
                        (N0)? mem[554] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] :
                        (N0)? mem[553] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] :
                        (N0)? mem[552] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] :
                        (N0)? mem[551] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] :
                        (N0)? mem[550] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] :
                        (N0)? mem[549] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] :
                        (N0)? mem[548] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] :
                        (N0)? mem[547] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] :
                       (N0)? mem[546] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] :
                       (N0)? mem[545] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] :
                       (N0)? mem[544] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] :
                       (N0)? mem[543] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] :
                       (N0)? mem[542] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] :
                       (N0)? mem[541] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] :
                       (N0)? mem[540] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] :
                       (N0)? mem[539] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] :
                       (N0)? mem[538] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] :
                       (N0)? mem[537] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], N5, N5, N5, N5, N5, N5 } :
                                                                       (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N13) begin
      { mem[1073:975], mem[537:537] } <= { w_data_i[536:438], w_data_i[0:0] };
    end
    if(N14) begin
      { mem[974:876], mem[538:538] } <= { w_data_i[437:339], w_data_i[1:1] };
    end
    if(N15) begin
      { mem[875:777], mem[539:539] } <= { w_data_i[338:240], w_data_i[2:2] };
    end
    if(N16) begin
      { mem[776:678], mem[540:540] } <= { w_data_i[239:141], w_data_i[3:3] };
    end
    if(N17) begin
      { mem[677:579], mem[541:541] } <= { w_data_i[140:42], w_data_i[4:4] };
    end
    if(N18) begin
      { mem[578:542] } <= { w_data_i[41:5] };
    end
    if(N7) begin
      { mem[536:438], mem[0:0] } <= { w_data_i[536:438], w_data_i[0:0] };
    end
    if(N8) begin
      { mem[437:339], mem[1:1] } <= { w_data_i[437:339], w_data_i[1:1] };
    end
    if(N9) begin
      { mem[338:240], mem[2:2] } <= { w_data_i[338:240], w_data_i[2:2] };
    end
    if(N10) begin
      { mem[239:141], mem[3:3] } <= { w_data_i[239:141], w_data_i[3:3] };
    end
    if(N11) begin
      { mem[140:42], mem[4:4] } <= { w_data_i[140:42], w_data_i[4:4] };
    end
    if(N12) begin
      { mem[41:5] } <= { w_data_i[41:5] };
    end
  end


endmodule



module bsg_mem_1r1w_width_p537_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [536:0] w_data_i;
  input [0:0] r_addr_i;
  output [536:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [536:0] r_data_o;

  bsg_mem_p537
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p537
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [536:0] data_i;
  output [536:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [536:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p537_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 :
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 :
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 :
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 :
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 :
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 :
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end
    if(N9) begin
      tail_r <= N10;
    end
    if(N11) begin
      head_r <= N12;
    end
  end


endmodule



module bsg_mem_p58
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [57:0] w_data_i;
  input [0:0] r_addr_i;
  output [57:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [57:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  reg [115:0] mem;
  assign r_data_o[57] = (N3)? mem[57] :
                        (N0)? mem[115] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[56] = (N3)? mem[56] :
                        (N0)? mem[114] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] :
                        (N0)? mem[113] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] :
                        (N0)? mem[112] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] :
                        (N0)? mem[111] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] :
                        (N0)? mem[110] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] :
                        (N0)? mem[109] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] :
                        (N0)? mem[108] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] :
                        (N0)? mem[107] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] :
                        (N0)? mem[106] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] :
                        (N0)? mem[105] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] :
                        (N0)? mem[104] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] :
                        (N0)? mem[103] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] :
                        (N0)? mem[102] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] :
                        (N0)? mem[101] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] :
                        (N0)? mem[100] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] :
                        (N0)? mem[99] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] :
                        (N0)? mem[98] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] :
                        (N0)? mem[97] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] :
                        (N0)? mem[96] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] :
                        (N0)? mem[95] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] :
                        (N0)? mem[94] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] :
                        (N0)? mem[93] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] :
                        (N0)? mem[92] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] :
                        (N0)? mem[91] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] :
                        (N0)? mem[90] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] :
                        (N0)? mem[89] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] :
                        (N0)? mem[88] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] :
                        (N0)? mem[87] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] :
                        (N0)? mem[86] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] :
                        (N0)? mem[85] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] :
                        (N0)? mem[84] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] :
                        (N0)? mem[83] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] :
                        (N0)? mem[82] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] :
                        (N0)? mem[81] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] :
                        (N0)? mem[80] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] :
                        (N0)? mem[79] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] :
                        (N0)? mem[78] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] :
                        (N0)? mem[77] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] :
                        (N0)? mem[76] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] :
                        (N0)? mem[75] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] :
                        (N0)? mem[74] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] :
                        (N0)? mem[73] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] :
                        (N0)? mem[72] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] :
                        (N0)? mem[71] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] :
                        (N0)? mem[70] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] :
                        (N0)? mem[69] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] :
                        (N0)? mem[68] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] :
                       (N0)? mem[67] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] :
                       (N0)? mem[66] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] :
                       (N0)? mem[65] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] :
                       (N0)? mem[64] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] :
                       (N0)? mem[63] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] :
                       (N0)? mem[62] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] :
                       (N0)? mem[61] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] :
                       (N0)? mem[60] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] :
                       (N0)? mem[59] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] :
                       (N0)? mem[58] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } :
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      { mem[115:58] } <= { w_data_i[57:0] };
    end
    if(N7) begin
      { mem[57:0] } <= { w_data_i[57:0] };
    end
  end


endmodule



module bsg_mem_1r1w_width_p58_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [57:0] w_data_i;
  input [0:0] r_addr_i;
  output [57:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [57:0] r_data_o;

  bsg_mem_p58
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p58
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [57:0] data_i;
  output [57:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [57:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p58_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 :
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 :
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 :
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 :
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 :
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 :
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end
    if(N9) begin
      tail_r <= N10;
    end
    if(N11) begin
      head_r <= N12;
    end
  end


endmodule



module bsg_mem_p542
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [541:0] w_data_i;
  input [0:0] r_addr_i;
  output [541:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [541:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;
  reg [1083:0] mem;
  assign r_data_o[541] = (N3)? mem[541] :
                         (N0)? mem[1083] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[540] = (N3)? mem[540] :
                         (N0)? mem[1082] : 1'b0;
  assign r_data_o[539] = (N3)? mem[539] :
                         (N0)? mem[1081] : 1'b0;
  assign r_data_o[538] = (N3)? mem[538] :
                         (N0)? mem[1080] : 1'b0;
  assign r_data_o[537] = (N3)? mem[537] :
                         (N0)? mem[1079] : 1'b0;
  assign r_data_o[536] = (N3)? mem[536] :
                         (N0)? mem[1078] : 1'b0;
  assign r_data_o[535] = (N3)? mem[535] :
                         (N0)? mem[1077] : 1'b0;
  assign r_data_o[534] = (N3)? mem[534] :
                         (N0)? mem[1076] : 1'b0;
  assign r_data_o[533] = (N3)? mem[533] :
                         (N0)? mem[1075] : 1'b0;
  assign r_data_o[532] = (N3)? mem[532] :
                         (N0)? mem[1074] : 1'b0;
  assign r_data_o[531] = (N3)? mem[531] :
                         (N0)? mem[1073] : 1'b0;
  assign r_data_o[530] = (N3)? mem[530] :
                         (N0)? mem[1072] : 1'b0;
  assign r_data_o[529] = (N3)? mem[529] :
                         (N0)? mem[1071] : 1'b0;
  assign r_data_o[528] = (N3)? mem[528] :
                         (N0)? mem[1070] : 1'b0;
  assign r_data_o[527] = (N3)? mem[527] :
                         (N0)? mem[1069] : 1'b0;
  assign r_data_o[526] = (N3)? mem[526] :
                         (N0)? mem[1068] : 1'b0;
  assign r_data_o[525] = (N3)? mem[525] :
                         (N0)? mem[1067] : 1'b0;
  assign r_data_o[524] = (N3)? mem[524] :
                         (N0)? mem[1066] : 1'b0;
  assign r_data_o[523] = (N3)? mem[523] :
                         (N0)? mem[1065] : 1'b0;
  assign r_data_o[522] = (N3)? mem[522] :
                         (N0)? mem[1064] : 1'b0;
  assign r_data_o[521] = (N3)? mem[521] :
                         (N0)? mem[1063] : 1'b0;
  assign r_data_o[520] = (N3)? mem[520] :
                         (N0)? mem[1062] : 1'b0;
  assign r_data_o[519] = (N3)? mem[519] :
                         (N0)? mem[1061] : 1'b0;
  assign r_data_o[518] = (N3)? mem[518] :
                         (N0)? mem[1060] : 1'b0;
  assign r_data_o[517] = (N3)? mem[517] :
                         (N0)? mem[1059] : 1'b0;
  assign r_data_o[516] = (N3)? mem[516] :
                         (N0)? mem[1058] : 1'b0;
  assign r_data_o[515] = (N3)? mem[515] :
                         (N0)? mem[1057] : 1'b0;
  assign r_data_o[514] = (N3)? mem[514] :
                         (N0)? mem[1056] : 1'b0;
  assign r_data_o[513] = (N3)? mem[513] :
                         (N0)? mem[1055] : 1'b0;
  assign r_data_o[512] = (N3)? mem[512] :
                         (N0)? mem[1054] : 1'b0;
  assign r_data_o[511] = (N3)? mem[511] :
                         (N0)? mem[1053] : 1'b0;
  assign r_data_o[510] = (N3)? mem[510] :
                         (N0)? mem[1052] : 1'b0;
  assign r_data_o[509] = (N3)? mem[509] :
                         (N0)? mem[1051] : 1'b0;
  assign r_data_o[508] = (N3)? mem[508] :
                         (N0)? mem[1050] : 1'b0;
  assign r_data_o[507] = (N3)? mem[507] :
                         (N0)? mem[1049] : 1'b0;
  assign r_data_o[506] = (N3)? mem[506] :
                         (N0)? mem[1048] : 1'b0;
  assign r_data_o[505] = (N3)? mem[505] :
                         (N0)? mem[1047] : 1'b0;
  assign r_data_o[504] = (N3)? mem[504] :
                         (N0)? mem[1046] : 1'b0;
  assign r_data_o[503] = (N3)? mem[503] :
                         (N0)? mem[1045] : 1'b0;
  assign r_data_o[502] = (N3)? mem[502] :
                         (N0)? mem[1044] : 1'b0;
  assign r_data_o[501] = (N3)? mem[501] :
                         (N0)? mem[1043] : 1'b0;
  assign r_data_o[500] = (N3)? mem[500] :
                         (N0)? mem[1042] : 1'b0;
  assign r_data_o[499] = (N3)? mem[499] :
                         (N0)? mem[1041] : 1'b0;
  assign r_data_o[498] = (N3)? mem[498] :
                         (N0)? mem[1040] : 1'b0;
  assign r_data_o[497] = (N3)? mem[497] :
                         (N0)? mem[1039] : 1'b0;
  assign r_data_o[496] = (N3)? mem[496] :
                         (N0)? mem[1038] : 1'b0;
  assign r_data_o[495] = (N3)? mem[495] :
                         (N0)? mem[1037] : 1'b0;
  assign r_data_o[494] = (N3)? mem[494] :
                         (N0)? mem[1036] : 1'b0;
  assign r_data_o[493] = (N3)? mem[493] :
                         (N0)? mem[1035] : 1'b0;
  assign r_data_o[492] = (N3)? mem[492] :
                         (N0)? mem[1034] : 1'b0;
  assign r_data_o[491] = (N3)? mem[491] :
                         (N0)? mem[1033] : 1'b0;
  assign r_data_o[490] = (N3)? mem[490] :
                         (N0)? mem[1032] : 1'b0;
  assign r_data_o[489] = (N3)? mem[489] :
                         (N0)? mem[1031] : 1'b0;
  assign r_data_o[488] = (N3)? mem[488] :
                         (N0)? mem[1030] : 1'b0;
  assign r_data_o[487] = (N3)? mem[487] :
                         (N0)? mem[1029] : 1'b0;
  assign r_data_o[486] = (N3)? mem[486] :
                         (N0)? mem[1028] : 1'b0;
  assign r_data_o[485] = (N3)? mem[485] :
                         (N0)? mem[1027] : 1'b0;
  assign r_data_o[484] = (N3)? mem[484] :
                         (N0)? mem[1026] : 1'b0;
  assign r_data_o[483] = (N3)? mem[483] :
                         (N0)? mem[1025] : 1'b0;
  assign r_data_o[482] = (N3)? mem[482] :
                         (N0)? mem[1024] : 1'b0;
  assign r_data_o[481] = (N3)? mem[481] :
                         (N0)? mem[1023] : 1'b0;
  assign r_data_o[480] = (N3)? mem[480] :
                         (N0)? mem[1022] : 1'b0;
  assign r_data_o[479] = (N3)? mem[479] :
                         (N0)? mem[1021] : 1'b0;
  assign r_data_o[478] = (N3)? mem[478] :
                         (N0)? mem[1020] : 1'b0;
  assign r_data_o[477] = (N3)? mem[477] :
                         (N0)? mem[1019] : 1'b0;
  assign r_data_o[476] = (N3)? mem[476] :
                         (N0)? mem[1018] : 1'b0;
  assign r_data_o[475] = (N3)? mem[475] :
                         (N0)? mem[1017] : 1'b0;
  assign r_data_o[474] = (N3)? mem[474] :
                         (N0)? mem[1016] : 1'b0;
  assign r_data_o[473] = (N3)? mem[473] :
                         (N0)? mem[1015] : 1'b0;
  assign r_data_o[472] = (N3)? mem[472] :
                         (N0)? mem[1014] : 1'b0;
  assign r_data_o[471] = (N3)? mem[471] :
                         (N0)? mem[1013] : 1'b0;
  assign r_data_o[470] = (N3)? mem[470] :
                         (N0)? mem[1012] : 1'b0;
  assign r_data_o[469] = (N3)? mem[469] :
                         (N0)? mem[1011] : 1'b0;
  assign r_data_o[468] = (N3)? mem[468] :
                         (N0)? mem[1010] : 1'b0;
  assign r_data_o[467] = (N3)? mem[467] :
                         (N0)? mem[1009] : 1'b0;
  assign r_data_o[466] = (N3)? mem[466] :
                         (N0)? mem[1008] : 1'b0;
  assign r_data_o[465] = (N3)? mem[465] :
                         (N0)? mem[1007] : 1'b0;
  assign r_data_o[464] = (N3)? mem[464] :
                         (N0)? mem[1006] : 1'b0;
  assign r_data_o[463] = (N3)? mem[463] :
                         (N0)? mem[1005] : 1'b0;
  assign r_data_o[462] = (N3)? mem[462] :
                         (N0)? mem[1004] : 1'b0;
  assign r_data_o[461] = (N3)? mem[461] :
                         (N0)? mem[1003] : 1'b0;
  assign r_data_o[460] = (N3)? mem[460] :
                         (N0)? mem[1002] : 1'b0;
  assign r_data_o[459] = (N3)? mem[459] :
                         (N0)? mem[1001] : 1'b0;
  assign r_data_o[458] = (N3)? mem[458] :
                         (N0)? mem[1000] : 1'b0;
  assign r_data_o[457] = (N3)? mem[457] :
                         (N0)? mem[999] : 1'b0;
  assign r_data_o[456] = (N3)? mem[456] :
                         (N0)? mem[998] : 1'b0;
  assign r_data_o[455] = (N3)? mem[455] :
                         (N0)? mem[997] : 1'b0;
  assign r_data_o[454] = (N3)? mem[454] :
                         (N0)? mem[996] : 1'b0;
  assign r_data_o[453] = (N3)? mem[453] :
                         (N0)? mem[995] : 1'b0;
  assign r_data_o[452] = (N3)? mem[452] :
                         (N0)? mem[994] : 1'b0;
  assign r_data_o[451] = (N3)? mem[451] :
                         (N0)? mem[993] : 1'b0;
  assign r_data_o[450] = (N3)? mem[450] :
                         (N0)? mem[992] : 1'b0;
  assign r_data_o[449] = (N3)? mem[449] :
                         (N0)? mem[991] : 1'b0;
  assign r_data_o[448] = (N3)? mem[448] :
                         (N0)? mem[990] : 1'b0;
  assign r_data_o[447] = (N3)? mem[447] :
                         (N0)? mem[989] : 1'b0;
  assign r_data_o[446] = (N3)? mem[446] :
                         (N0)? mem[988] : 1'b0;
  assign r_data_o[445] = (N3)? mem[445] :
                         (N0)? mem[987] : 1'b0;
  assign r_data_o[444] = (N3)? mem[444] :
                         (N0)? mem[986] : 1'b0;
  assign r_data_o[443] = (N3)? mem[443] :
                         (N0)? mem[985] : 1'b0;
  assign r_data_o[442] = (N3)? mem[442] :
                         (N0)? mem[984] : 1'b0;
  assign r_data_o[441] = (N3)? mem[441] :
                         (N0)? mem[983] : 1'b0;
  assign r_data_o[440] = (N3)? mem[440] :
                         (N0)? mem[982] : 1'b0;
  assign r_data_o[439] = (N3)? mem[439] :
                         (N0)? mem[981] : 1'b0;
  assign r_data_o[438] = (N3)? mem[438] :
                         (N0)? mem[980] : 1'b0;
  assign r_data_o[437] = (N3)? mem[437] :
                         (N0)? mem[979] : 1'b0;
  assign r_data_o[436] = (N3)? mem[436] :
                         (N0)? mem[978] : 1'b0;
  assign r_data_o[435] = (N3)? mem[435] :
                         (N0)? mem[977] : 1'b0;
  assign r_data_o[434] = (N3)? mem[434] :
                         (N0)? mem[976] : 1'b0;
  assign r_data_o[433] = (N3)? mem[433] :
                         (N0)? mem[975] : 1'b0;
  assign r_data_o[432] = (N3)? mem[432] :
                         (N0)? mem[974] : 1'b0;
  assign r_data_o[431] = (N3)? mem[431] :
                         (N0)? mem[973] : 1'b0;
  assign r_data_o[430] = (N3)? mem[430] :
                         (N0)? mem[972] : 1'b0;
  assign r_data_o[429] = (N3)? mem[429] :
                         (N0)? mem[971] : 1'b0;
  assign r_data_o[428] = (N3)? mem[428] :
                         (N0)? mem[970] : 1'b0;
  assign r_data_o[427] = (N3)? mem[427] :
                         (N0)? mem[969] : 1'b0;
  assign r_data_o[426] = (N3)? mem[426] :
                         (N0)? mem[968] : 1'b0;
  assign r_data_o[425] = (N3)? mem[425] :
                         (N0)? mem[967] : 1'b0;
  assign r_data_o[424] = (N3)? mem[424] :
                         (N0)? mem[966] : 1'b0;
  assign r_data_o[423] = (N3)? mem[423] :
                         (N0)? mem[965] : 1'b0;
  assign r_data_o[422] = (N3)? mem[422] :
                         (N0)? mem[964] : 1'b0;
  assign r_data_o[421] = (N3)? mem[421] :
                         (N0)? mem[963] : 1'b0;
  assign r_data_o[420] = (N3)? mem[420] :
                         (N0)? mem[962] : 1'b0;
  assign r_data_o[419] = (N3)? mem[419] :
                         (N0)? mem[961] : 1'b0;
  assign r_data_o[418] = (N3)? mem[418] :
                         (N0)? mem[960] : 1'b0;
  assign r_data_o[417] = (N3)? mem[417] :
                         (N0)? mem[959] : 1'b0;
  assign r_data_o[416] = (N3)? mem[416] :
                         (N0)? mem[958] : 1'b0;
  assign r_data_o[415] = (N3)? mem[415] :
                         (N0)? mem[957] : 1'b0;
  assign r_data_o[414] = (N3)? mem[414] :
                         (N0)? mem[956] : 1'b0;
  assign r_data_o[413] = (N3)? mem[413] :
                         (N0)? mem[955] : 1'b0;
  assign r_data_o[412] = (N3)? mem[412] :
                         (N0)? mem[954] : 1'b0;
  assign r_data_o[411] = (N3)? mem[411] :
                         (N0)? mem[953] : 1'b0;
  assign r_data_o[410] = (N3)? mem[410] :
                         (N0)? mem[952] : 1'b0;
  assign r_data_o[409] = (N3)? mem[409] :
                         (N0)? mem[951] : 1'b0;
  assign r_data_o[408] = (N3)? mem[408] :
                         (N0)? mem[950] : 1'b0;
  assign r_data_o[407] = (N3)? mem[407] :
                         (N0)? mem[949] : 1'b0;
  assign r_data_o[406] = (N3)? mem[406] :
                         (N0)? mem[948] : 1'b0;
  assign r_data_o[405] = (N3)? mem[405] :
                         (N0)? mem[947] : 1'b0;
  assign r_data_o[404] = (N3)? mem[404] :
                         (N0)? mem[946] : 1'b0;
  assign r_data_o[403] = (N3)? mem[403] :
                         (N0)? mem[945] : 1'b0;
  assign r_data_o[402] = (N3)? mem[402] :
                         (N0)? mem[944] : 1'b0;
  assign r_data_o[401] = (N3)? mem[401] :
                         (N0)? mem[943] : 1'b0;
  assign r_data_o[400] = (N3)? mem[400] :
                         (N0)? mem[942] : 1'b0;
  assign r_data_o[399] = (N3)? mem[399] :
                         (N0)? mem[941] : 1'b0;
  assign r_data_o[398] = (N3)? mem[398] :
                         (N0)? mem[940] : 1'b0;
  assign r_data_o[397] = (N3)? mem[397] :
                         (N0)? mem[939] : 1'b0;
  assign r_data_o[396] = (N3)? mem[396] :
                         (N0)? mem[938] : 1'b0;
  assign r_data_o[395] = (N3)? mem[395] :
                         (N0)? mem[937] : 1'b0;
  assign r_data_o[394] = (N3)? mem[394] :
                         (N0)? mem[936] : 1'b0;
  assign r_data_o[393] = (N3)? mem[393] :
                         (N0)? mem[935] : 1'b0;
  assign r_data_o[392] = (N3)? mem[392] :
                         (N0)? mem[934] : 1'b0;
  assign r_data_o[391] = (N3)? mem[391] :
                         (N0)? mem[933] : 1'b0;
  assign r_data_o[390] = (N3)? mem[390] :
                         (N0)? mem[932] : 1'b0;
  assign r_data_o[389] = (N3)? mem[389] :
                         (N0)? mem[931] : 1'b0;
  assign r_data_o[388] = (N3)? mem[388] :
                         (N0)? mem[930] : 1'b0;
  assign r_data_o[387] = (N3)? mem[387] :
                         (N0)? mem[929] : 1'b0;
  assign r_data_o[386] = (N3)? mem[386] :
                         (N0)? mem[928] : 1'b0;
  assign r_data_o[385] = (N3)? mem[385] :
                         (N0)? mem[927] : 1'b0;
  assign r_data_o[384] = (N3)? mem[384] :
                         (N0)? mem[926] : 1'b0;
  assign r_data_o[383] = (N3)? mem[383] :
                         (N0)? mem[925] : 1'b0;
  assign r_data_o[382] = (N3)? mem[382] :
                         (N0)? mem[924] : 1'b0;
  assign r_data_o[381] = (N3)? mem[381] :
                         (N0)? mem[923] : 1'b0;
  assign r_data_o[380] = (N3)? mem[380] :
                         (N0)? mem[922] : 1'b0;
  assign r_data_o[379] = (N3)? mem[379] :
                         (N0)? mem[921] : 1'b0;
  assign r_data_o[378] = (N3)? mem[378] :
                         (N0)? mem[920] : 1'b0;
  assign r_data_o[377] = (N3)? mem[377] :
                         (N0)? mem[919] : 1'b0;
  assign r_data_o[376] = (N3)? mem[376] :
                         (N0)? mem[918] : 1'b0;
  assign r_data_o[375] = (N3)? mem[375] :
                         (N0)? mem[917] : 1'b0;
  assign r_data_o[374] = (N3)? mem[374] :
                         (N0)? mem[916] : 1'b0;
  assign r_data_o[373] = (N3)? mem[373] :
                         (N0)? mem[915] : 1'b0;
  assign r_data_o[372] = (N3)? mem[372] :
                         (N0)? mem[914] : 1'b0;
  assign r_data_o[371] = (N3)? mem[371] :
                         (N0)? mem[913] : 1'b0;
  assign r_data_o[370] = (N3)? mem[370] :
                         (N0)? mem[912] : 1'b0;
  assign r_data_o[369] = (N3)? mem[369] :
                         (N0)? mem[911] : 1'b0;
  assign r_data_o[368] = (N3)? mem[368] :
                         (N0)? mem[910] : 1'b0;
  assign r_data_o[367] = (N3)? mem[367] :
                         (N0)? mem[909] : 1'b0;
  assign r_data_o[366] = (N3)? mem[366] :
                         (N0)? mem[908] : 1'b0;
  assign r_data_o[365] = (N3)? mem[365] :
                         (N0)? mem[907] : 1'b0;
  assign r_data_o[364] = (N3)? mem[364] :
                         (N0)? mem[906] : 1'b0;
  assign r_data_o[363] = (N3)? mem[363] :
                         (N0)? mem[905] : 1'b0;
  assign r_data_o[362] = (N3)? mem[362] :
                         (N0)? mem[904] : 1'b0;
  assign r_data_o[361] = (N3)? mem[361] :
                         (N0)? mem[903] : 1'b0;
  assign r_data_o[360] = (N3)? mem[360] :
                         (N0)? mem[902] : 1'b0;
  assign r_data_o[359] = (N3)? mem[359] :
                         (N0)? mem[901] : 1'b0;
  assign r_data_o[358] = (N3)? mem[358] :
                         (N0)? mem[900] : 1'b0;
  assign r_data_o[357] = (N3)? mem[357] :
                         (N0)? mem[899] : 1'b0;
  assign r_data_o[356] = (N3)? mem[356] :
                         (N0)? mem[898] : 1'b0;
  assign r_data_o[355] = (N3)? mem[355] :
                         (N0)? mem[897] : 1'b0;
  assign r_data_o[354] = (N3)? mem[354] :
                         (N0)? mem[896] : 1'b0;
  assign r_data_o[353] = (N3)? mem[353] :
                         (N0)? mem[895] : 1'b0;
  assign r_data_o[352] = (N3)? mem[352] :
                         (N0)? mem[894] : 1'b0;
  assign r_data_o[351] = (N3)? mem[351] :
                         (N0)? mem[893] : 1'b0;
  assign r_data_o[350] = (N3)? mem[350] :
                         (N0)? mem[892] : 1'b0;
  assign r_data_o[349] = (N3)? mem[349] :
                         (N0)? mem[891] : 1'b0;
  assign r_data_o[348] = (N3)? mem[348] :
                         (N0)? mem[890] : 1'b0;
  assign r_data_o[347] = (N3)? mem[347] :
                         (N0)? mem[889] : 1'b0;
  assign r_data_o[346] = (N3)? mem[346] :
                         (N0)? mem[888] : 1'b0;
  assign r_data_o[345] = (N3)? mem[345] :
                         (N0)? mem[887] : 1'b0;
  assign r_data_o[344] = (N3)? mem[344] :
                         (N0)? mem[886] : 1'b0;
  assign r_data_o[343] = (N3)? mem[343] :
                         (N0)? mem[885] : 1'b0;
  assign r_data_o[342] = (N3)? mem[342] :
                         (N0)? mem[884] : 1'b0;
  assign r_data_o[341] = (N3)? mem[341] :
                         (N0)? mem[883] : 1'b0;
  assign r_data_o[340] = (N3)? mem[340] :
                         (N0)? mem[882] : 1'b0;
  assign r_data_o[339] = (N3)? mem[339] :
                         (N0)? mem[881] : 1'b0;
  assign r_data_o[338] = (N3)? mem[338] :
                         (N0)? mem[880] : 1'b0;
  assign r_data_o[337] = (N3)? mem[337] :
                         (N0)? mem[879] : 1'b0;
  assign r_data_o[336] = (N3)? mem[336] :
                         (N0)? mem[878] : 1'b0;
  assign r_data_o[335] = (N3)? mem[335] :
                         (N0)? mem[877] : 1'b0;
  assign r_data_o[334] = (N3)? mem[334] :
                         (N0)? mem[876] : 1'b0;
  assign r_data_o[333] = (N3)? mem[333] :
                         (N0)? mem[875] : 1'b0;
  assign r_data_o[332] = (N3)? mem[332] :
                         (N0)? mem[874] : 1'b0;
  assign r_data_o[331] = (N3)? mem[331] :
                         (N0)? mem[873] : 1'b0;
  assign r_data_o[330] = (N3)? mem[330] :
                         (N0)? mem[872] : 1'b0;
  assign r_data_o[329] = (N3)? mem[329] :
                         (N0)? mem[871] : 1'b0;
  assign r_data_o[328] = (N3)? mem[328] :
                         (N0)? mem[870] : 1'b0;
  assign r_data_o[327] = (N3)? mem[327] :
                         (N0)? mem[869] : 1'b0;
  assign r_data_o[326] = (N3)? mem[326] :
                         (N0)? mem[868] : 1'b0;
  assign r_data_o[325] = (N3)? mem[325] :
                         (N0)? mem[867] : 1'b0;
  assign r_data_o[324] = (N3)? mem[324] :
                         (N0)? mem[866] : 1'b0;
  assign r_data_o[323] = (N3)? mem[323] :
                         (N0)? mem[865] : 1'b0;
  assign r_data_o[322] = (N3)? mem[322] :
                         (N0)? mem[864] : 1'b0;
  assign r_data_o[321] = (N3)? mem[321] :
                         (N0)? mem[863] : 1'b0;
  assign r_data_o[320] = (N3)? mem[320] :
                         (N0)? mem[862] : 1'b0;
  assign r_data_o[319] = (N3)? mem[319] :
                         (N0)? mem[861] : 1'b0;
  assign r_data_o[318] = (N3)? mem[318] :
                         (N0)? mem[860] : 1'b0;
  assign r_data_o[317] = (N3)? mem[317] :
                         (N0)? mem[859] : 1'b0;
  assign r_data_o[316] = (N3)? mem[316] :
                         (N0)? mem[858] : 1'b0;
  assign r_data_o[315] = (N3)? mem[315] :
                         (N0)? mem[857] : 1'b0;
  assign r_data_o[314] = (N3)? mem[314] :
                         (N0)? mem[856] : 1'b0;
  assign r_data_o[313] = (N3)? mem[313] :
                         (N0)? mem[855] : 1'b0;
  assign r_data_o[312] = (N3)? mem[312] :
                         (N0)? mem[854] : 1'b0;
  assign r_data_o[311] = (N3)? mem[311] :
                         (N0)? mem[853] : 1'b0;
  assign r_data_o[310] = (N3)? mem[310] :
                         (N0)? mem[852] : 1'b0;
  assign r_data_o[309] = (N3)? mem[309] :
                         (N0)? mem[851] : 1'b0;
  assign r_data_o[308] = (N3)? mem[308] :
                         (N0)? mem[850] : 1'b0;
  assign r_data_o[307] = (N3)? mem[307] :
                         (N0)? mem[849] : 1'b0;
  assign r_data_o[306] = (N3)? mem[306] :
                         (N0)? mem[848] : 1'b0;
  assign r_data_o[305] = (N3)? mem[305] :
                         (N0)? mem[847] : 1'b0;
  assign r_data_o[304] = (N3)? mem[304] :
                         (N0)? mem[846] : 1'b0;
  assign r_data_o[303] = (N3)? mem[303] :
                         (N0)? mem[845] : 1'b0;
  assign r_data_o[302] = (N3)? mem[302] :
                         (N0)? mem[844] : 1'b0;
  assign r_data_o[301] = (N3)? mem[301] :
                         (N0)? mem[843] : 1'b0;
  assign r_data_o[300] = (N3)? mem[300] :
                         (N0)? mem[842] : 1'b0;
  assign r_data_o[299] = (N3)? mem[299] :
                         (N0)? mem[841] : 1'b0;
  assign r_data_o[298] = (N3)? mem[298] :
                         (N0)? mem[840] : 1'b0;
  assign r_data_o[297] = (N3)? mem[297] :
                         (N0)? mem[839] : 1'b0;
  assign r_data_o[296] = (N3)? mem[296] :
                         (N0)? mem[838] : 1'b0;
  assign r_data_o[295] = (N3)? mem[295] :
                         (N0)? mem[837] : 1'b0;
  assign r_data_o[294] = (N3)? mem[294] :
                         (N0)? mem[836] : 1'b0;
  assign r_data_o[293] = (N3)? mem[293] :
                         (N0)? mem[835] : 1'b0;
  assign r_data_o[292] = (N3)? mem[292] :
                         (N0)? mem[834] : 1'b0;
  assign r_data_o[291] = (N3)? mem[291] :
                         (N0)? mem[833] : 1'b0;
  assign r_data_o[290] = (N3)? mem[290] :
                         (N0)? mem[832] : 1'b0;
  assign r_data_o[289] = (N3)? mem[289] :
                         (N0)? mem[831] : 1'b0;
  assign r_data_o[288] = (N3)? mem[288] :
                         (N0)? mem[830] : 1'b0;
  assign r_data_o[287] = (N3)? mem[287] :
                         (N0)? mem[829] : 1'b0;
  assign r_data_o[286] = (N3)? mem[286] :
                         (N0)? mem[828] : 1'b0;
  assign r_data_o[285] = (N3)? mem[285] :
                         (N0)? mem[827] : 1'b0;
  assign r_data_o[284] = (N3)? mem[284] :
                         (N0)? mem[826] : 1'b0;
  assign r_data_o[283] = (N3)? mem[283] :
                         (N0)? mem[825] : 1'b0;
  assign r_data_o[282] = (N3)? mem[282] :
                         (N0)? mem[824] : 1'b0;
  assign r_data_o[281] = (N3)? mem[281] :
                         (N0)? mem[823] : 1'b0;
  assign r_data_o[280] = (N3)? mem[280] :
                         (N0)? mem[822] : 1'b0;
  assign r_data_o[279] = (N3)? mem[279] :
                         (N0)? mem[821] : 1'b0;
  assign r_data_o[278] = (N3)? mem[278] :
                         (N0)? mem[820] : 1'b0;
  assign r_data_o[277] = (N3)? mem[277] :
                         (N0)? mem[819] : 1'b0;
  assign r_data_o[276] = (N3)? mem[276] :
                         (N0)? mem[818] : 1'b0;
  assign r_data_o[275] = (N3)? mem[275] :
                         (N0)? mem[817] : 1'b0;
  assign r_data_o[274] = (N3)? mem[274] :
                         (N0)? mem[816] : 1'b0;
  assign r_data_o[273] = (N3)? mem[273] :
                         (N0)? mem[815] : 1'b0;
  assign r_data_o[272] = (N3)? mem[272] :
                         (N0)? mem[814] : 1'b0;
  assign r_data_o[271] = (N3)? mem[271] :
                         (N0)? mem[813] : 1'b0;
  assign r_data_o[270] = (N3)? mem[270] :
                         (N0)? mem[812] : 1'b0;
  assign r_data_o[269] = (N3)? mem[269] :
                         (N0)? mem[811] : 1'b0;
  assign r_data_o[268] = (N3)? mem[268] :
                         (N0)? mem[810] : 1'b0;
  assign r_data_o[267] = (N3)? mem[267] :
                         (N0)? mem[809] : 1'b0;
  assign r_data_o[266] = (N3)? mem[266] :
                         (N0)? mem[808] : 1'b0;
  assign r_data_o[265] = (N3)? mem[265] :
                         (N0)? mem[807] : 1'b0;
  assign r_data_o[264] = (N3)? mem[264] :
                         (N0)? mem[806] : 1'b0;
  assign r_data_o[263] = (N3)? mem[263] :
                         (N0)? mem[805] : 1'b0;
  assign r_data_o[262] = (N3)? mem[262] :
                         (N0)? mem[804] : 1'b0;
  assign r_data_o[261] = (N3)? mem[261] :
                         (N0)? mem[803] : 1'b0;
  assign r_data_o[260] = (N3)? mem[260] :
                         (N0)? mem[802] : 1'b0;
  assign r_data_o[259] = (N3)? mem[259] :
                         (N0)? mem[801] : 1'b0;
  assign r_data_o[258] = (N3)? mem[258] :
                         (N0)? mem[800] : 1'b0;
  assign r_data_o[257] = (N3)? mem[257] :
                         (N0)? mem[799] : 1'b0;
  assign r_data_o[256] = (N3)? mem[256] :
                         (N0)? mem[798] : 1'b0;
  assign r_data_o[255] = (N3)? mem[255] :
                         (N0)? mem[797] : 1'b0;
  assign r_data_o[254] = (N3)? mem[254] :
                         (N0)? mem[796] : 1'b0;
  assign r_data_o[253] = (N3)? mem[253] :
                         (N0)? mem[795] : 1'b0;
  assign r_data_o[252] = (N3)? mem[252] :
                         (N0)? mem[794] : 1'b0;
  assign r_data_o[251] = (N3)? mem[251] :
                         (N0)? mem[793] : 1'b0;
  assign r_data_o[250] = (N3)? mem[250] :
                         (N0)? mem[792] : 1'b0;
  assign r_data_o[249] = (N3)? mem[249] :
                         (N0)? mem[791] : 1'b0;
  assign r_data_o[248] = (N3)? mem[248] :
                         (N0)? mem[790] : 1'b0;
  assign r_data_o[247] = (N3)? mem[247] :
                         (N0)? mem[789] : 1'b0;
  assign r_data_o[246] = (N3)? mem[246] :
                         (N0)? mem[788] : 1'b0;
  assign r_data_o[245] = (N3)? mem[245] :
                         (N0)? mem[787] : 1'b0;
  assign r_data_o[244] = (N3)? mem[244] :
                         (N0)? mem[786] : 1'b0;
  assign r_data_o[243] = (N3)? mem[243] :
                         (N0)? mem[785] : 1'b0;
  assign r_data_o[242] = (N3)? mem[242] :
                         (N0)? mem[784] : 1'b0;
  assign r_data_o[241] = (N3)? mem[241] :
                         (N0)? mem[783] : 1'b0;
  assign r_data_o[240] = (N3)? mem[240] :
                         (N0)? mem[782] : 1'b0;
  assign r_data_o[239] = (N3)? mem[239] :
                         (N0)? mem[781] : 1'b0;
  assign r_data_o[238] = (N3)? mem[238] :
                         (N0)? mem[780] : 1'b0;
  assign r_data_o[237] = (N3)? mem[237] :
                         (N0)? mem[779] : 1'b0;
  assign r_data_o[236] = (N3)? mem[236] :
                         (N0)? mem[778] : 1'b0;
  assign r_data_o[235] = (N3)? mem[235] :
                         (N0)? mem[777] : 1'b0;
  assign r_data_o[234] = (N3)? mem[234] :
                         (N0)? mem[776] : 1'b0;
  assign r_data_o[233] = (N3)? mem[233] :
                         (N0)? mem[775] : 1'b0;
  assign r_data_o[232] = (N3)? mem[232] :
                         (N0)? mem[774] : 1'b0;
  assign r_data_o[231] = (N3)? mem[231] :
                         (N0)? mem[773] : 1'b0;
  assign r_data_o[230] = (N3)? mem[230] :
                         (N0)? mem[772] : 1'b0;
  assign r_data_o[229] = (N3)? mem[229] :
                         (N0)? mem[771] : 1'b0;
  assign r_data_o[228] = (N3)? mem[228] :
                         (N0)? mem[770] : 1'b0;
  assign r_data_o[227] = (N3)? mem[227] :
                         (N0)? mem[769] : 1'b0;
  assign r_data_o[226] = (N3)? mem[226] :
                         (N0)? mem[768] : 1'b0;
  assign r_data_o[225] = (N3)? mem[225] :
                         (N0)? mem[767] : 1'b0;
  assign r_data_o[224] = (N3)? mem[224] :
                         (N0)? mem[766] : 1'b0;
  assign r_data_o[223] = (N3)? mem[223] :
                         (N0)? mem[765] : 1'b0;
  assign r_data_o[222] = (N3)? mem[222] :
                         (N0)? mem[764] : 1'b0;
  assign r_data_o[221] = (N3)? mem[221] :
                         (N0)? mem[763] : 1'b0;
  assign r_data_o[220] = (N3)? mem[220] :
                         (N0)? mem[762] : 1'b0;
  assign r_data_o[219] = (N3)? mem[219] :
                         (N0)? mem[761] : 1'b0;
  assign r_data_o[218] = (N3)? mem[218] :
                         (N0)? mem[760] : 1'b0;
  assign r_data_o[217] = (N3)? mem[217] :
                         (N0)? mem[759] : 1'b0;
  assign r_data_o[216] = (N3)? mem[216] :
                         (N0)? mem[758] : 1'b0;
  assign r_data_o[215] = (N3)? mem[215] :
                         (N0)? mem[757] : 1'b0;
  assign r_data_o[214] = (N3)? mem[214] :
                         (N0)? mem[756] : 1'b0;
  assign r_data_o[213] = (N3)? mem[213] :
                         (N0)? mem[755] : 1'b0;
  assign r_data_o[212] = (N3)? mem[212] :
                         (N0)? mem[754] : 1'b0;
  assign r_data_o[211] = (N3)? mem[211] :
                         (N0)? mem[753] : 1'b0;
  assign r_data_o[210] = (N3)? mem[210] :
                         (N0)? mem[752] : 1'b0;
  assign r_data_o[209] = (N3)? mem[209] :
                         (N0)? mem[751] : 1'b0;
  assign r_data_o[208] = (N3)? mem[208] :
                         (N0)? mem[750] : 1'b0;
  assign r_data_o[207] = (N3)? mem[207] :
                         (N0)? mem[749] : 1'b0;
  assign r_data_o[206] = (N3)? mem[206] :
                         (N0)? mem[748] : 1'b0;
  assign r_data_o[205] = (N3)? mem[205] :
                         (N0)? mem[747] : 1'b0;
  assign r_data_o[204] = (N3)? mem[204] :
                         (N0)? mem[746] : 1'b0;
  assign r_data_o[203] = (N3)? mem[203] :
                         (N0)? mem[745] : 1'b0;
  assign r_data_o[202] = (N3)? mem[202] :
                         (N0)? mem[744] : 1'b0;
  assign r_data_o[201] = (N3)? mem[201] :
                         (N0)? mem[743] : 1'b0;
  assign r_data_o[200] = (N3)? mem[200] :
                         (N0)? mem[742] : 1'b0;
  assign r_data_o[199] = (N3)? mem[199] :
                         (N0)? mem[741] : 1'b0;
  assign r_data_o[198] = (N3)? mem[198] :
                         (N0)? mem[740] : 1'b0;
  assign r_data_o[197] = (N3)? mem[197] :
                         (N0)? mem[739] : 1'b0;
  assign r_data_o[196] = (N3)? mem[196] :
                         (N0)? mem[738] : 1'b0;
  assign r_data_o[195] = (N3)? mem[195] :
                         (N0)? mem[737] : 1'b0;
  assign r_data_o[194] = (N3)? mem[194] :
                         (N0)? mem[736] : 1'b0;
  assign r_data_o[193] = (N3)? mem[193] :
                         (N0)? mem[735] : 1'b0;
  assign r_data_o[192] = (N3)? mem[192] :
                         (N0)? mem[734] : 1'b0;
  assign r_data_o[191] = (N3)? mem[191] :
                         (N0)? mem[733] : 1'b0;
  assign r_data_o[190] = (N3)? mem[190] :
                         (N0)? mem[732] : 1'b0;
  assign r_data_o[189] = (N3)? mem[189] :
                         (N0)? mem[731] : 1'b0;
  assign r_data_o[188] = (N3)? mem[188] :
                         (N0)? mem[730] : 1'b0;
  assign r_data_o[187] = (N3)? mem[187] :
                         (N0)? mem[729] : 1'b0;
  assign r_data_o[186] = (N3)? mem[186] :
                         (N0)? mem[728] : 1'b0;
  assign r_data_o[185] = (N3)? mem[185] :
                         (N0)? mem[727] : 1'b0;
  assign r_data_o[184] = (N3)? mem[184] :
                         (N0)? mem[726] : 1'b0;
  assign r_data_o[183] = (N3)? mem[183] :
                         (N0)? mem[725] : 1'b0;
  assign r_data_o[182] = (N3)? mem[182] :
                         (N0)? mem[724] : 1'b0;
  assign r_data_o[181] = (N3)? mem[181] :
                         (N0)? mem[723] : 1'b0;
  assign r_data_o[180] = (N3)? mem[180] :
                         (N0)? mem[722] : 1'b0;
  assign r_data_o[179] = (N3)? mem[179] :
                         (N0)? mem[721] : 1'b0;
  assign r_data_o[178] = (N3)? mem[178] :
                         (N0)? mem[720] : 1'b0;
  assign r_data_o[177] = (N3)? mem[177] :
                         (N0)? mem[719] : 1'b0;
  assign r_data_o[176] = (N3)? mem[176] :
                         (N0)? mem[718] : 1'b0;
  assign r_data_o[175] = (N3)? mem[175] :
                         (N0)? mem[717] : 1'b0;
  assign r_data_o[174] = (N3)? mem[174] :
                         (N0)? mem[716] : 1'b0;
  assign r_data_o[173] = (N3)? mem[173] :
                         (N0)? mem[715] : 1'b0;
  assign r_data_o[172] = (N3)? mem[172] :
                         (N0)? mem[714] : 1'b0;
  assign r_data_o[171] = (N3)? mem[171] :
                         (N0)? mem[713] : 1'b0;
  assign r_data_o[170] = (N3)? mem[170] :
                         (N0)? mem[712] : 1'b0;
  assign r_data_o[169] = (N3)? mem[169] :
                         (N0)? mem[711] : 1'b0;
  assign r_data_o[168] = (N3)? mem[168] :
                         (N0)? mem[710] : 1'b0;
  assign r_data_o[167] = (N3)? mem[167] :
                         (N0)? mem[709] : 1'b0;
  assign r_data_o[166] = (N3)? mem[166] :
                         (N0)? mem[708] : 1'b0;
  assign r_data_o[165] = (N3)? mem[165] :
                         (N0)? mem[707] : 1'b0;
  assign r_data_o[164] = (N3)? mem[164] :
                         (N0)? mem[706] : 1'b0;
  assign r_data_o[163] = (N3)? mem[163] :
                         (N0)? mem[705] : 1'b0;
  assign r_data_o[162] = (N3)? mem[162] :
                         (N0)? mem[704] : 1'b0;
  assign r_data_o[161] = (N3)? mem[161] :
                         (N0)? mem[703] : 1'b0;
  assign r_data_o[160] = (N3)? mem[160] :
                         (N0)? mem[702] : 1'b0;
  assign r_data_o[159] = (N3)? mem[159] :
                         (N0)? mem[701] : 1'b0;
  assign r_data_o[158] = (N3)? mem[158] :
                         (N0)? mem[700] : 1'b0;
  assign r_data_o[157] = (N3)? mem[157] :
                         (N0)? mem[699] : 1'b0;
  assign r_data_o[156] = (N3)? mem[156] :
                         (N0)? mem[698] : 1'b0;
  assign r_data_o[155] = (N3)? mem[155] :
                         (N0)? mem[697] : 1'b0;
  assign r_data_o[154] = (N3)? mem[154] :
                         (N0)? mem[696] : 1'b0;
  assign r_data_o[153] = (N3)? mem[153] :
                         (N0)? mem[695] : 1'b0;
  assign r_data_o[152] = (N3)? mem[152] :
                         (N0)? mem[694] : 1'b0;
  assign r_data_o[151] = (N3)? mem[151] :
                         (N0)? mem[693] : 1'b0;
  assign r_data_o[150] = (N3)? mem[150] :
                         (N0)? mem[692] : 1'b0;
  assign r_data_o[149] = (N3)? mem[149] :
                         (N0)? mem[691] : 1'b0;
  assign r_data_o[148] = (N3)? mem[148] :
                         (N0)? mem[690] : 1'b0;
  assign r_data_o[147] = (N3)? mem[147] :
                         (N0)? mem[689] : 1'b0;
  assign r_data_o[146] = (N3)? mem[146] :
                         (N0)? mem[688] : 1'b0;
  assign r_data_o[145] = (N3)? mem[145] :
                         (N0)? mem[687] : 1'b0;
  assign r_data_o[144] = (N3)? mem[144] :
                         (N0)? mem[686] : 1'b0;
  assign r_data_o[143] = (N3)? mem[143] :
                         (N0)? mem[685] : 1'b0;
  assign r_data_o[142] = (N3)? mem[142] :
                         (N0)? mem[684] : 1'b0;
  assign r_data_o[141] = (N3)? mem[141] :
                         (N0)? mem[683] : 1'b0;
  assign r_data_o[140] = (N3)? mem[140] :
                         (N0)? mem[682] : 1'b0;
  assign r_data_o[139] = (N3)? mem[139] :
                         (N0)? mem[681] : 1'b0;
  assign r_data_o[138] = (N3)? mem[138] :
                         (N0)? mem[680] : 1'b0;
  assign r_data_o[137] = (N3)? mem[137] :
                         (N0)? mem[679] : 1'b0;
  assign r_data_o[136] = (N3)? mem[136] :
                         (N0)? mem[678] : 1'b0;
  assign r_data_o[135] = (N3)? mem[135] :
                         (N0)? mem[677] : 1'b0;
  assign r_data_o[134] = (N3)? mem[134] :
                         (N0)? mem[676] : 1'b0;
  assign r_data_o[133] = (N3)? mem[133] :
                         (N0)? mem[675] : 1'b0;
  assign r_data_o[132] = (N3)? mem[132] :
                         (N0)? mem[674] : 1'b0;
  assign r_data_o[131] = (N3)? mem[131] :
                         (N0)? mem[673] : 1'b0;
  assign r_data_o[130] = (N3)? mem[130] :
                         (N0)? mem[672] : 1'b0;
  assign r_data_o[129] = (N3)? mem[129] :
                         (N0)? mem[671] : 1'b0;
  assign r_data_o[128] = (N3)? mem[128] :
                         (N0)? mem[670] : 1'b0;
  assign r_data_o[127] = (N3)? mem[127] :
                         (N0)? mem[669] : 1'b0;
  assign r_data_o[126] = (N3)? mem[126] :
                         (N0)? mem[668] : 1'b0;
  assign r_data_o[125] = (N3)? mem[125] :
                         (N0)? mem[667] : 1'b0;
  assign r_data_o[124] = (N3)? mem[124] :
                         (N0)? mem[666] : 1'b0;
  assign r_data_o[123] = (N3)? mem[123] :
                         (N0)? mem[665] : 1'b0;
  assign r_data_o[122] = (N3)? mem[122] :
                         (N0)? mem[664] : 1'b0;
  assign r_data_o[121] = (N3)? mem[121] :
                         (N0)? mem[663] : 1'b0;
  assign r_data_o[120] = (N3)? mem[120] :
                         (N0)? mem[662] : 1'b0;
  assign r_data_o[119] = (N3)? mem[119] :
                         (N0)? mem[661] : 1'b0;
  assign r_data_o[118] = (N3)? mem[118] :
                         (N0)? mem[660] : 1'b0;
  assign r_data_o[117] = (N3)? mem[117] :
                         (N0)? mem[659] : 1'b0;
  assign r_data_o[116] = (N3)? mem[116] :
                         (N0)? mem[658] : 1'b0;
  assign r_data_o[115] = (N3)? mem[115] :
                         (N0)? mem[657] : 1'b0;
  assign r_data_o[114] = (N3)? mem[114] :
                         (N0)? mem[656] : 1'b0;
  assign r_data_o[113] = (N3)? mem[113] :
                         (N0)? mem[655] : 1'b0;
  assign r_data_o[112] = (N3)? mem[112] :
                         (N0)? mem[654] : 1'b0;
  assign r_data_o[111] = (N3)? mem[111] :
                         (N0)? mem[653] : 1'b0;
  assign r_data_o[110] = (N3)? mem[110] :
                         (N0)? mem[652] : 1'b0;
  assign r_data_o[109] = (N3)? mem[109] :
                         (N0)? mem[651] : 1'b0;
  assign r_data_o[108] = (N3)? mem[108] :
                         (N0)? mem[650] : 1'b0;
  assign r_data_o[107] = (N3)? mem[107] :
                         (N0)? mem[649] : 1'b0;
  assign r_data_o[106] = (N3)? mem[106] :
                         (N0)? mem[648] : 1'b0;
  assign r_data_o[105] = (N3)? mem[105] :
                         (N0)? mem[647] : 1'b0;
  assign r_data_o[104] = (N3)? mem[104] :
                         (N0)? mem[646] : 1'b0;
  assign r_data_o[103] = (N3)? mem[103] :
                         (N0)? mem[645] : 1'b0;
  assign r_data_o[102] = (N3)? mem[102] :
                         (N0)? mem[644] : 1'b0;
  assign r_data_o[101] = (N3)? mem[101] :
                         (N0)? mem[643] : 1'b0;
  assign r_data_o[100] = (N3)? mem[100] :
                         (N0)? mem[642] : 1'b0;
  assign r_data_o[99] = (N3)? mem[99] :
                        (N0)? mem[641] : 1'b0;
  assign r_data_o[98] = (N3)? mem[98] :
                        (N0)? mem[640] : 1'b0;
  assign r_data_o[97] = (N3)? mem[97] :
                        (N0)? mem[639] : 1'b0;
  assign r_data_o[96] = (N3)? mem[96] :
                        (N0)? mem[638] : 1'b0;
  assign r_data_o[95] = (N3)? mem[95] :
                        (N0)? mem[637] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] :
                        (N0)? mem[636] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] :
                        (N0)? mem[635] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] :
                        (N0)? mem[634] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] :
                        (N0)? mem[633] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] :
                        (N0)? mem[632] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] :
                        (N0)? mem[631] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] :
                        (N0)? mem[630] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] :
                        (N0)? mem[629] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] :
                        (N0)? mem[628] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] :
                        (N0)? mem[627] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] :
                        (N0)? mem[626] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] :
                        (N0)? mem[625] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] :
                        (N0)? mem[624] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] :
                        (N0)? mem[623] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] :
                        (N0)? mem[622] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] :
                        (N0)? mem[621] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] :
                        (N0)? mem[620] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] :
                        (N0)? mem[619] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] :
                        (N0)? mem[618] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] :
                        (N0)? mem[617] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] :
                        (N0)? mem[616] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] :
                        (N0)? mem[615] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] :
                        (N0)? mem[614] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] :
                        (N0)? mem[613] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] :
                        (N0)? mem[612] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] :
                        (N0)? mem[611] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] :
                        (N0)? mem[610] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] :
                        (N0)? mem[609] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] :
                        (N0)? mem[608] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] :
                        (N0)? mem[607] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] :
                        (N0)? mem[606] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] :
                        (N0)? mem[605] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] :
                        (N0)? mem[604] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] :
                        (N0)? mem[603] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] :
                        (N0)? mem[602] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] :
                        (N0)? mem[601] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] :
                        (N0)? mem[600] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] :
                        (N0)? mem[599] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] :
                        (N0)? mem[598] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] :
                        (N0)? mem[597] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] :
                        (N0)? mem[596] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] :
                        (N0)? mem[595] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] :
                        (N0)? mem[594] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] :
                        (N0)? mem[593] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] :
                        (N0)? mem[592] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] :
                        (N0)? mem[591] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] :
                        (N0)? mem[590] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] :
                        (N0)? mem[589] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] :
                        (N0)? mem[588] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] :
                        (N0)? mem[587] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] :
                        (N0)? mem[586] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] :
                        (N0)? mem[585] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] :
                        (N0)? mem[584] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] :
                        (N0)? mem[583] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] :
                        (N0)? mem[582] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] :
                        (N0)? mem[581] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] :
                        (N0)? mem[580] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] :
                        (N0)? mem[579] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] :
                        (N0)? mem[578] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] :
                        (N0)? mem[577] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] :
                        (N0)? mem[576] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] :
                        (N0)? mem[575] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] :
                        (N0)? mem[574] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] :
                        (N0)? mem[573] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] :
                        (N0)? mem[572] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] :
                        (N0)? mem[571] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] :
                        (N0)? mem[570] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] :
                        (N0)? mem[569] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] :
                        (N0)? mem[568] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] :
                        (N0)? mem[567] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] :
                        (N0)? mem[566] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] :
                        (N0)? mem[565] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] :
                        (N0)? mem[564] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] :
                        (N0)? mem[563] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] :
                        (N0)? mem[562] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] :
                        (N0)? mem[561] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] :
                        (N0)? mem[560] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] :
                        (N0)? mem[559] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] :
                        (N0)? mem[558] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] :
                        (N0)? mem[557] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] :
                        (N0)? mem[556] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] :
                        (N0)? mem[555] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] :
                        (N0)? mem[554] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] :
                        (N0)? mem[553] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] :
                        (N0)? mem[552] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] :
                       (N0)? mem[551] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] :
                       (N0)? mem[550] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] :
                       (N0)? mem[549] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] :
                       (N0)? mem[548] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] :
                       (N0)? mem[547] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] :
                       (N0)? mem[546] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] :
                       (N0)? mem[545] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] :
                       (N0)? mem[544] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] :
                       (N0)? mem[543] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] :
                       (N0)? mem[542] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], N5, N5, N5, N5, N5, N5 } :
                                                                       (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N13) begin
      { mem[1083:985], mem[542:542] } <= { w_data_i[541:443], w_data_i[0:0] };
    end
    if(N14) begin
      { mem[984:886], mem[543:543] } <= { w_data_i[442:344], w_data_i[1:1] };
    end
    if(N15) begin
      { mem[885:787], mem[544:544] } <= { w_data_i[343:245], w_data_i[2:2] };
    end
    if(N16) begin
      { mem[786:688], mem[545:545] } <= { w_data_i[244:146], w_data_i[3:3] };
    end
    if(N17) begin
      { mem[687:589], mem[546:546] } <= { w_data_i[145:47], w_data_i[4:4] };
    end
    if(N18) begin
      { mem[588:547] } <= { w_data_i[46:5] };
    end
    if(N7) begin
      { mem[541:443], mem[0:0] } <= { w_data_i[541:443], w_data_i[0:0] };
    end
    if(N8) begin
      { mem[442:344], mem[1:1] } <= { w_data_i[442:344], w_data_i[1:1] };
    end
    if(N9) begin
      { mem[343:245], mem[2:2] } <= { w_data_i[343:245], w_data_i[2:2] };
    end
    if(N10) begin
      { mem[244:146], mem[3:3] } <= { w_data_i[244:146], w_data_i[3:3] };
    end
    if(N11) begin
      { mem[145:47], mem[4:4] } <= { w_data_i[145:47], w_data_i[4:4] };
    end
    if(N12) begin
      { mem[46:5] } <= { w_data_i[46:5] };
    end
  end


endmodule



module bsg_mem_1r1w_width_p542_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [541:0] w_data_i;
  input [0:0] r_addr_i;
  output [541:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [541:0] r_data_o;

  bsg_mem_p542
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p542
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [541:0] data_i;
  output [541:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [541:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p542_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 :
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 :
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 :
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 :
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 :
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 :
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end
    if(N9) begin
      tail_r <= N10;
    end
    if(N11) begin
      head_r <= N12;
    end
  end


endmodule



module bsg_mem_p30
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [29:0] w_data_i;
  input [0:0] r_addr_i;
  output [29:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [29:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  reg [59:0] mem;
  assign r_data_o[29] = (N3)? mem[29] :
                        (N0)? mem[59] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[28] = (N3)? mem[28] :
                        (N0)? mem[58] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] :
                        (N0)? mem[57] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] :
                        (N0)? mem[56] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] :
                        (N0)? mem[55] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] :
                        (N0)? mem[54] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] :
                        (N0)? mem[53] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] :
                        (N0)? mem[52] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] :
                        (N0)? mem[51] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] :
                        (N0)? mem[50] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] :
                        (N0)? mem[49] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] :
                        (N0)? mem[48] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] :
                        (N0)? mem[47] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] :
                        (N0)? mem[46] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] :
                        (N0)? mem[45] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] :
                        (N0)? mem[44] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] :
                        (N0)? mem[43] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] :
                        (N0)? mem[42] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] :
                        (N0)? mem[41] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] :
                        (N0)? mem[40] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] :
                       (N0)? mem[39] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] :
                       (N0)? mem[38] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] :
                       (N0)? mem[37] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] :
                       (N0)? mem[36] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] :
                       (N0)? mem[35] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] :
                       (N0)? mem[34] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] :
                       (N0)? mem[33] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] :
                       (N0)? mem[32] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] :
                       (N0)? mem[31] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] :
                       (N0)? mem[30] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } :
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      { mem[59:30] } <= { w_data_i[29:0] };
    end
    if(N7) begin
      { mem[29:0] } <= { w_data_i[29:0] };
    end
  end


endmodule



module bsg_mem_1r1w_width_p30_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [29:0] w_data_i;
  input [0:0] r_addr_i;
  output [29:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [29:0] r_data_o;

  bsg_mem_p30
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p30
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [29:0] data_i;
  output [29:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [29:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p30_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 :
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 :
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 :
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 :
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 :
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 :
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end
    if(N9) begin
      tail_r <= N10;
    end
    if(N11) begin
      head_r <= N12;
    end
  end


endmodule



module bsg_mem_p570
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [569:0] w_data_i;
  input [0:0] r_addr_i;
  output [569:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [569:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;
  reg [1139:0] mem;
  assign r_data_o[569] = (N3)? mem[569] :
                         (N0)? mem[1139] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[568] = (N3)? mem[568] :
                         (N0)? mem[1138] : 1'b0;
  assign r_data_o[567] = (N3)? mem[567] :
                         (N0)? mem[1137] : 1'b0;
  assign r_data_o[566] = (N3)? mem[566] :
                         (N0)? mem[1136] : 1'b0;
  assign r_data_o[565] = (N3)? mem[565] :
                         (N0)? mem[1135] : 1'b0;
  assign r_data_o[564] = (N3)? mem[564] :
                         (N0)? mem[1134] : 1'b0;
  assign r_data_o[563] = (N3)? mem[563] :
                         (N0)? mem[1133] : 1'b0;
  assign r_data_o[562] = (N3)? mem[562] :
                         (N0)? mem[1132] : 1'b0;
  assign r_data_o[561] = (N3)? mem[561] :
                         (N0)? mem[1131] : 1'b0;
  assign r_data_o[560] = (N3)? mem[560] :
                         (N0)? mem[1130] : 1'b0;
  assign r_data_o[559] = (N3)? mem[559] :
                         (N0)? mem[1129] : 1'b0;
  assign r_data_o[558] = (N3)? mem[558] :
                         (N0)? mem[1128] : 1'b0;
  assign r_data_o[557] = (N3)? mem[557] :
                         (N0)? mem[1127] : 1'b0;
  assign r_data_o[556] = (N3)? mem[556] :
                         (N0)? mem[1126] : 1'b0;
  assign r_data_o[555] = (N3)? mem[555] :
                         (N0)? mem[1125] : 1'b0;
  assign r_data_o[554] = (N3)? mem[554] :
                         (N0)? mem[1124] : 1'b0;
  assign r_data_o[553] = (N3)? mem[553] :
                         (N0)? mem[1123] : 1'b0;
  assign r_data_o[552] = (N3)? mem[552] :
                         (N0)? mem[1122] : 1'b0;
  assign r_data_o[551] = (N3)? mem[551] :
                         (N0)? mem[1121] : 1'b0;
  assign r_data_o[550] = (N3)? mem[550] :
                         (N0)? mem[1120] : 1'b0;
  assign r_data_o[549] = (N3)? mem[549] :
                         (N0)? mem[1119] : 1'b0;
  assign r_data_o[548] = (N3)? mem[548] :
                         (N0)? mem[1118] : 1'b0;
  assign r_data_o[547] = (N3)? mem[547] :
                         (N0)? mem[1117] : 1'b0;
  assign r_data_o[546] = (N3)? mem[546] :
                         (N0)? mem[1116] : 1'b0;
  assign r_data_o[545] = (N3)? mem[545] :
                         (N0)? mem[1115] : 1'b0;
  assign r_data_o[544] = (N3)? mem[544] :
                         (N0)? mem[1114] : 1'b0;
  assign r_data_o[543] = (N3)? mem[543] :
                         (N0)? mem[1113] : 1'b0;
  assign r_data_o[542] = (N3)? mem[542] :
                         (N0)? mem[1112] : 1'b0;
  assign r_data_o[541] = (N3)? mem[541] :
                         (N0)? mem[1111] : 1'b0;
  assign r_data_o[540] = (N3)? mem[540] :
                         (N0)? mem[1110] : 1'b0;
  assign r_data_o[539] = (N3)? mem[539] :
                         (N0)? mem[1109] : 1'b0;
  assign r_data_o[538] = (N3)? mem[538] :
                         (N0)? mem[1108] : 1'b0;
  assign r_data_o[537] = (N3)? mem[537] :
                         (N0)? mem[1107] : 1'b0;
  assign r_data_o[536] = (N3)? mem[536] :
                         (N0)? mem[1106] : 1'b0;
  assign r_data_o[535] = (N3)? mem[535] :
                         (N0)? mem[1105] : 1'b0;
  assign r_data_o[534] = (N3)? mem[534] :
                         (N0)? mem[1104] : 1'b0;
  assign r_data_o[533] = (N3)? mem[533] :
                         (N0)? mem[1103] : 1'b0;
  assign r_data_o[532] = (N3)? mem[532] :
                         (N0)? mem[1102] : 1'b0;
  assign r_data_o[531] = (N3)? mem[531] :
                         (N0)? mem[1101] : 1'b0;
  assign r_data_o[530] = (N3)? mem[530] :
                         (N0)? mem[1100] : 1'b0;
  assign r_data_o[529] = (N3)? mem[529] :
                         (N0)? mem[1099] : 1'b0;
  assign r_data_o[528] = (N3)? mem[528] :
                         (N0)? mem[1098] : 1'b0;
  assign r_data_o[527] = (N3)? mem[527] :
                         (N0)? mem[1097] : 1'b0;
  assign r_data_o[526] = (N3)? mem[526] :
                         (N0)? mem[1096] : 1'b0;
  assign r_data_o[525] = (N3)? mem[525] :
                         (N0)? mem[1095] : 1'b0;
  assign r_data_o[524] = (N3)? mem[524] :
                         (N0)? mem[1094] : 1'b0;
  assign r_data_o[523] = (N3)? mem[523] :
                         (N0)? mem[1093] : 1'b0;
  assign r_data_o[522] = (N3)? mem[522] :
                         (N0)? mem[1092] : 1'b0;
  assign r_data_o[521] = (N3)? mem[521] :
                         (N0)? mem[1091] : 1'b0;
  assign r_data_o[520] = (N3)? mem[520] :
                         (N0)? mem[1090] : 1'b0;
  assign r_data_o[519] = (N3)? mem[519] :
                         (N0)? mem[1089] : 1'b0;
  assign r_data_o[518] = (N3)? mem[518] :
                         (N0)? mem[1088] : 1'b0;
  assign r_data_o[517] = (N3)? mem[517] :
                         (N0)? mem[1087] : 1'b0;
  assign r_data_o[516] = (N3)? mem[516] :
                         (N0)? mem[1086] : 1'b0;
  assign r_data_o[515] = (N3)? mem[515] :
                         (N0)? mem[1085] : 1'b0;
  assign r_data_o[514] = (N3)? mem[514] :
                         (N0)? mem[1084] : 1'b0;
  assign r_data_o[513] = (N3)? mem[513] :
                         (N0)? mem[1083] : 1'b0;
  assign r_data_o[512] = (N3)? mem[512] :
                         (N0)? mem[1082] : 1'b0;
  assign r_data_o[511] = (N3)? mem[511] :
                         (N0)? mem[1081] : 1'b0;
  assign r_data_o[510] = (N3)? mem[510] :
                         (N0)? mem[1080] : 1'b0;
  assign r_data_o[509] = (N3)? mem[509] :
                         (N0)? mem[1079] : 1'b0;
  assign r_data_o[508] = (N3)? mem[508] :
                         (N0)? mem[1078] : 1'b0;
  assign r_data_o[507] = (N3)? mem[507] :
                         (N0)? mem[1077] : 1'b0;
  assign r_data_o[506] = (N3)? mem[506] :
                         (N0)? mem[1076] : 1'b0;
  assign r_data_o[505] = (N3)? mem[505] :
                         (N0)? mem[1075] : 1'b0;
  assign r_data_o[504] = (N3)? mem[504] :
                         (N0)? mem[1074] : 1'b0;
  assign r_data_o[503] = (N3)? mem[503] :
                         (N0)? mem[1073] : 1'b0;
  assign r_data_o[502] = (N3)? mem[502] :
                         (N0)? mem[1072] : 1'b0;
  assign r_data_o[501] = (N3)? mem[501] :
                         (N0)? mem[1071] : 1'b0;
  assign r_data_o[500] = (N3)? mem[500] :
                         (N0)? mem[1070] : 1'b0;
  assign r_data_o[499] = (N3)? mem[499] :
                         (N0)? mem[1069] : 1'b0;
  assign r_data_o[498] = (N3)? mem[498] :
                         (N0)? mem[1068] : 1'b0;
  assign r_data_o[497] = (N3)? mem[497] :
                         (N0)? mem[1067] : 1'b0;
  assign r_data_o[496] = (N3)? mem[496] :
                         (N0)? mem[1066] : 1'b0;
  assign r_data_o[495] = (N3)? mem[495] :
                         (N0)? mem[1065] : 1'b0;
  assign r_data_o[494] = (N3)? mem[494] :
                         (N0)? mem[1064] : 1'b0;
  assign r_data_o[493] = (N3)? mem[493] :
                         (N0)? mem[1063] : 1'b0;
  assign r_data_o[492] = (N3)? mem[492] :
                         (N0)? mem[1062] : 1'b0;
  assign r_data_o[491] = (N3)? mem[491] :
                         (N0)? mem[1061] : 1'b0;
  assign r_data_o[490] = (N3)? mem[490] :
                         (N0)? mem[1060] : 1'b0;
  assign r_data_o[489] = (N3)? mem[489] :
                         (N0)? mem[1059] : 1'b0;
  assign r_data_o[488] = (N3)? mem[488] :
                         (N0)? mem[1058] : 1'b0;
  assign r_data_o[487] = (N3)? mem[487] :
                         (N0)? mem[1057] : 1'b0;
  assign r_data_o[486] = (N3)? mem[486] :
                         (N0)? mem[1056] : 1'b0;
  assign r_data_o[485] = (N3)? mem[485] :
                         (N0)? mem[1055] : 1'b0;
  assign r_data_o[484] = (N3)? mem[484] :
                         (N0)? mem[1054] : 1'b0;
  assign r_data_o[483] = (N3)? mem[483] :
                         (N0)? mem[1053] : 1'b0;
  assign r_data_o[482] = (N3)? mem[482] :
                         (N0)? mem[1052] : 1'b0;
  assign r_data_o[481] = (N3)? mem[481] :
                         (N0)? mem[1051] : 1'b0;
  assign r_data_o[480] = (N3)? mem[480] :
                         (N0)? mem[1050] : 1'b0;
  assign r_data_o[479] = (N3)? mem[479] :
                         (N0)? mem[1049] : 1'b0;
  assign r_data_o[478] = (N3)? mem[478] :
                         (N0)? mem[1048] : 1'b0;
  assign r_data_o[477] = (N3)? mem[477] :
                         (N0)? mem[1047] : 1'b0;
  assign r_data_o[476] = (N3)? mem[476] :
                         (N0)? mem[1046] : 1'b0;
  assign r_data_o[475] = (N3)? mem[475] :
                         (N0)? mem[1045] : 1'b0;
  assign r_data_o[474] = (N3)? mem[474] :
                         (N0)? mem[1044] : 1'b0;
  assign r_data_o[473] = (N3)? mem[473] :
                         (N0)? mem[1043] : 1'b0;
  assign r_data_o[472] = (N3)? mem[472] :
                         (N0)? mem[1042] : 1'b0;
  assign r_data_o[471] = (N3)? mem[471] :
                         (N0)? mem[1041] : 1'b0;
  assign r_data_o[470] = (N3)? mem[470] :
                         (N0)? mem[1040] : 1'b0;
  assign r_data_o[469] = (N3)? mem[469] :
                         (N0)? mem[1039] : 1'b0;
  assign r_data_o[468] = (N3)? mem[468] :
                         (N0)? mem[1038] : 1'b0;
  assign r_data_o[467] = (N3)? mem[467] :
                         (N0)? mem[1037] : 1'b0;
  assign r_data_o[466] = (N3)? mem[466] :
                         (N0)? mem[1036] : 1'b0;
  assign r_data_o[465] = (N3)? mem[465] :
                         (N0)? mem[1035] : 1'b0;
  assign r_data_o[464] = (N3)? mem[464] :
                         (N0)? mem[1034] : 1'b0;
  assign r_data_o[463] = (N3)? mem[463] :
                         (N0)? mem[1033] : 1'b0;
  assign r_data_o[462] = (N3)? mem[462] :
                         (N0)? mem[1032] : 1'b0;
  assign r_data_o[461] = (N3)? mem[461] :
                         (N0)? mem[1031] : 1'b0;
  assign r_data_o[460] = (N3)? mem[460] :
                         (N0)? mem[1030] : 1'b0;
  assign r_data_o[459] = (N3)? mem[459] :
                         (N0)? mem[1029] : 1'b0;
  assign r_data_o[458] = (N3)? mem[458] :
                         (N0)? mem[1028] : 1'b0;
  assign r_data_o[457] = (N3)? mem[457] :
                         (N0)? mem[1027] : 1'b0;
  assign r_data_o[456] = (N3)? mem[456] :
                         (N0)? mem[1026] : 1'b0;
  assign r_data_o[455] = (N3)? mem[455] :
                         (N0)? mem[1025] : 1'b0;
  assign r_data_o[454] = (N3)? mem[454] :
                         (N0)? mem[1024] : 1'b0;
  assign r_data_o[453] = (N3)? mem[453] :
                         (N0)? mem[1023] : 1'b0;
  assign r_data_o[452] = (N3)? mem[452] :
                         (N0)? mem[1022] : 1'b0;
  assign r_data_o[451] = (N3)? mem[451] :
                         (N0)? mem[1021] : 1'b0;
  assign r_data_o[450] = (N3)? mem[450] :
                         (N0)? mem[1020] : 1'b0;
  assign r_data_o[449] = (N3)? mem[449] :
                         (N0)? mem[1019] : 1'b0;
  assign r_data_o[448] = (N3)? mem[448] :
                         (N0)? mem[1018] : 1'b0;
  assign r_data_o[447] = (N3)? mem[447] :
                         (N0)? mem[1017] : 1'b0;
  assign r_data_o[446] = (N3)? mem[446] :
                         (N0)? mem[1016] : 1'b0;
  assign r_data_o[445] = (N3)? mem[445] :
                         (N0)? mem[1015] : 1'b0;
  assign r_data_o[444] = (N3)? mem[444] :
                         (N0)? mem[1014] : 1'b0;
  assign r_data_o[443] = (N3)? mem[443] :
                         (N0)? mem[1013] : 1'b0;
  assign r_data_o[442] = (N3)? mem[442] :
                         (N0)? mem[1012] : 1'b0;
  assign r_data_o[441] = (N3)? mem[441] :
                         (N0)? mem[1011] : 1'b0;
  assign r_data_o[440] = (N3)? mem[440] :
                         (N0)? mem[1010] : 1'b0;
  assign r_data_o[439] = (N3)? mem[439] :
                         (N0)? mem[1009] : 1'b0;
  assign r_data_o[438] = (N3)? mem[438] :
                         (N0)? mem[1008] : 1'b0;
  assign r_data_o[437] = (N3)? mem[437] :
                         (N0)? mem[1007] : 1'b0;
  assign r_data_o[436] = (N3)? mem[436] :
                         (N0)? mem[1006] : 1'b0;
  assign r_data_o[435] = (N3)? mem[435] :
                         (N0)? mem[1005] : 1'b0;
  assign r_data_o[434] = (N3)? mem[434] :
                         (N0)? mem[1004] : 1'b0;
  assign r_data_o[433] = (N3)? mem[433] :
                         (N0)? mem[1003] : 1'b0;
  assign r_data_o[432] = (N3)? mem[432] :
                         (N0)? mem[1002] : 1'b0;
  assign r_data_o[431] = (N3)? mem[431] :
                         (N0)? mem[1001] : 1'b0;
  assign r_data_o[430] = (N3)? mem[430] :
                         (N0)? mem[1000] : 1'b0;
  assign r_data_o[429] = (N3)? mem[429] :
                         (N0)? mem[999] : 1'b0;
  assign r_data_o[428] = (N3)? mem[428] :
                         (N0)? mem[998] : 1'b0;
  assign r_data_o[427] = (N3)? mem[427] :
                         (N0)? mem[997] : 1'b0;
  assign r_data_o[426] = (N3)? mem[426] :
                         (N0)? mem[996] : 1'b0;
  assign r_data_o[425] = (N3)? mem[425] :
                         (N0)? mem[995] : 1'b0;
  assign r_data_o[424] = (N3)? mem[424] :
                         (N0)? mem[994] : 1'b0;
  assign r_data_o[423] = (N3)? mem[423] :
                         (N0)? mem[993] : 1'b0;
  assign r_data_o[422] = (N3)? mem[422] :
                         (N0)? mem[992] : 1'b0;
  assign r_data_o[421] = (N3)? mem[421] :
                         (N0)? mem[991] : 1'b0;
  assign r_data_o[420] = (N3)? mem[420] :
                         (N0)? mem[990] : 1'b0;
  assign r_data_o[419] = (N3)? mem[419] :
                         (N0)? mem[989] : 1'b0;
  assign r_data_o[418] = (N3)? mem[418] :
                         (N0)? mem[988] : 1'b0;
  assign r_data_o[417] = (N3)? mem[417] :
                         (N0)? mem[987] : 1'b0;
  assign r_data_o[416] = (N3)? mem[416] :
                         (N0)? mem[986] : 1'b0;
  assign r_data_o[415] = (N3)? mem[415] :
                         (N0)? mem[985] : 1'b0;
  assign r_data_o[414] = (N3)? mem[414] :
                         (N0)? mem[984] : 1'b0;
  assign r_data_o[413] = (N3)? mem[413] :
                         (N0)? mem[983] : 1'b0;
  assign r_data_o[412] = (N3)? mem[412] :
                         (N0)? mem[982] : 1'b0;
  assign r_data_o[411] = (N3)? mem[411] :
                         (N0)? mem[981] : 1'b0;
  assign r_data_o[410] = (N3)? mem[410] :
                         (N0)? mem[980] : 1'b0;
  assign r_data_o[409] = (N3)? mem[409] :
                         (N0)? mem[979] : 1'b0;
  assign r_data_o[408] = (N3)? mem[408] :
                         (N0)? mem[978] : 1'b0;
  assign r_data_o[407] = (N3)? mem[407] :
                         (N0)? mem[977] : 1'b0;
  assign r_data_o[406] = (N3)? mem[406] :
                         (N0)? mem[976] : 1'b0;
  assign r_data_o[405] = (N3)? mem[405] :
                         (N0)? mem[975] : 1'b0;
  assign r_data_o[404] = (N3)? mem[404] :
                         (N0)? mem[974] : 1'b0;
  assign r_data_o[403] = (N3)? mem[403] :
                         (N0)? mem[973] : 1'b0;
  assign r_data_o[402] = (N3)? mem[402] :
                         (N0)? mem[972] : 1'b0;
  assign r_data_o[401] = (N3)? mem[401] :
                         (N0)? mem[971] : 1'b0;
  assign r_data_o[400] = (N3)? mem[400] :
                         (N0)? mem[970] : 1'b0;
  assign r_data_o[399] = (N3)? mem[399] :
                         (N0)? mem[969] : 1'b0;
  assign r_data_o[398] = (N3)? mem[398] :
                         (N0)? mem[968] : 1'b0;
  assign r_data_o[397] = (N3)? mem[397] :
                         (N0)? mem[967] : 1'b0;
  assign r_data_o[396] = (N3)? mem[396] :
                         (N0)? mem[966] : 1'b0;
  assign r_data_o[395] = (N3)? mem[395] :
                         (N0)? mem[965] : 1'b0;
  assign r_data_o[394] = (N3)? mem[394] :
                         (N0)? mem[964] : 1'b0;
  assign r_data_o[393] = (N3)? mem[393] :
                         (N0)? mem[963] : 1'b0;
  assign r_data_o[392] = (N3)? mem[392] :
                         (N0)? mem[962] : 1'b0;
  assign r_data_o[391] = (N3)? mem[391] :
                         (N0)? mem[961] : 1'b0;
  assign r_data_o[390] = (N3)? mem[390] :
                         (N0)? mem[960] : 1'b0;
  assign r_data_o[389] = (N3)? mem[389] :
                         (N0)? mem[959] : 1'b0;
  assign r_data_o[388] = (N3)? mem[388] :
                         (N0)? mem[958] : 1'b0;
  assign r_data_o[387] = (N3)? mem[387] :
                         (N0)? mem[957] : 1'b0;
  assign r_data_o[386] = (N3)? mem[386] :
                         (N0)? mem[956] : 1'b0;
  assign r_data_o[385] = (N3)? mem[385] :
                         (N0)? mem[955] : 1'b0;
  assign r_data_o[384] = (N3)? mem[384] :
                         (N0)? mem[954] : 1'b0;
  assign r_data_o[383] = (N3)? mem[383] :
                         (N0)? mem[953] : 1'b0;
  assign r_data_o[382] = (N3)? mem[382] :
                         (N0)? mem[952] : 1'b0;
  assign r_data_o[381] = (N3)? mem[381] :
                         (N0)? mem[951] : 1'b0;
  assign r_data_o[380] = (N3)? mem[380] :
                         (N0)? mem[950] : 1'b0;
  assign r_data_o[379] = (N3)? mem[379] :
                         (N0)? mem[949] : 1'b0;
  assign r_data_o[378] = (N3)? mem[378] :
                         (N0)? mem[948] : 1'b0;
  assign r_data_o[377] = (N3)? mem[377] :
                         (N0)? mem[947] : 1'b0;
  assign r_data_o[376] = (N3)? mem[376] :
                         (N0)? mem[946] : 1'b0;
  assign r_data_o[375] = (N3)? mem[375] :
                         (N0)? mem[945] : 1'b0;
  assign r_data_o[374] = (N3)? mem[374] :
                         (N0)? mem[944] : 1'b0;
  assign r_data_o[373] = (N3)? mem[373] :
                         (N0)? mem[943] : 1'b0;
  assign r_data_o[372] = (N3)? mem[372] :
                         (N0)? mem[942] : 1'b0;
  assign r_data_o[371] = (N3)? mem[371] :
                         (N0)? mem[941] : 1'b0;
  assign r_data_o[370] = (N3)? mem[370] :
                         (N0)? mem[940] : 1'b0;
  assign r_data_o[369] = (N3)? mem[369] :
                         (N0)? mem[939] : 1'b0;
  assign r_data_o[368] = (N3)? mem[368] :
                         (N0)? mem[938] : 1'b0;
  assign r_data_o[367] = (N3)? mem[367] :
                         (N0)? mem[937] : 1'b0;
  assign r_data_o[366] = (N3)? mem[366] :
                         (N0)? mem[936] : 1'b0;
  assign r_data_o[365] = (N3)? mem[365] :
                         (N0)? mem[935] : 1'b0;
  assign r_data_o[364] = (N3)? mem[364] :
                         (N0)? mem[934] : 1'b0;
  assign r_data_o[363] = (N3)? mem[363] :
                         (N0)? mem[933] : 1'b0;
  assign r_data_o[362] = (N3)? mem[362] :
                         (N0)? mem[932] : 1'b0;
  assign r_data_o[361] = (N3)? mem[361] :
                         (N0)? mem[931] : 1'b0;
  assign r_data_o[360] = (N3)? mem[360] :
                         (N0)? mem[930] : 1'b0;
  assign r_data_o[359] = (N3)? mem[359] :
                         (N0)? mem[929] : 1'b0;
  assign r_data_o[358] = (N3)? mem[358] :
                         (N0)? mem[928] : 1'b0;
  assign r_data_o[357] = (N3)? mem[357] :
                         (N0)? mem[927] : 1'b0;
  assign r_data_o[356] = (N3)? mem[356] :
                         (N0)? mem[926] : 1'b0;
  assign r_data_o[355] = (N3)? mem[355] :
                         (N0)? mem[925] : 1'b0;
  assign r_data_o[354] = (N3)? mem[354] :
                         (N0)? mem[924] : 1'b0;
  assign r_data_o[353] = (N3)? mem[353] :
                         (N0)? mem[923] : 1'b0;
  assign r_data_o[352] = (N3)? mem[352] :
                         (N0)? mem[922] : 1'b0;
  assign r_data_o[351] = (N3)? mem[351] :
                         (N0)? mem[921] : 1'b0;
  assign r_data_o[350] = (N3)? mem[350] :
                         (N0)? mem[920] : 1'b0;
  assign r_data_o[349] = (N3)? mem[349] :
                         (N0)? mem[919] : 1'b0;
  assign r_data_o[348] = (N3)? mem[348] :
                         (N0)? mem[918] : 1'b0;
  assign r_data_o[347] = (N3)? mem[347] :
                         (N0)? mem[917] : 1'b0;
  assign r_data_o[346] = (N3)? mem[346] :
                         (N0)? mem[916] : 1'b0;
  assign r_data_o[345] = (N3)? mem[345] :
                         (N0)? mem[915] : 1'b0;
  assign r_data_o[344] = (N3)? mem[344] :
                         (N0)? mem[914] : 1'b0;
  assign r_data_o[343] = (N3)? mem[343] :
                         (N0)? mem[913] : 1'b0;
  assign r_data_o[342] = (N3)? mem[342] :
                         (N0)? mem[912] : 1'b0;
  assign r_data_o[341] = (N3)? mem[341] :
                         (N0)? mem[911] : 1'b0;
  assign r_data_o[340] = (N3)? mem[340] :
                         (N0)? mem[910] : 1'b0;
  assign r_data_o[339] = (N3)? mem[339] :
                         (N0)? mem[909] : 1'b0;
  assign r_data_o[338] = (N3)? mem[338] :
                         (N0)? mem[908] : 1'b0;
  assign r_data_o[337] = (N3)? mem[337] :
                         (N0)? mem[907] : 1'b0;
  assign r_data_o[336] = (N3)? mem[336] :
                         (N0)? mem[906] : 1'b0;
  assign r_data_o[335] = (N3)? mem[335] :
                         (N0)? mem[905] : 1'b0;
  assign r_data_o[334] = (N3)? mem[334] :
                         (N0)? mem[904] : 1'b0;
  assign r_data_o[333] = (N3)? mem[333] :
                         (N0)? mem[903] : 1'b0;
  assign r_data_o[332] = (N3)? mem[332] :
                         (N0)? mem[902] : 1'b0;
  assign r_data_o[331] = (N3)? mem[331] :
                         (N0)? mem[901] : 1'b0;
  assign r_data_o[330] = (N3)? mem[330] :
                         (N0)? mem[900] : 1'b0;
  assign r_data_o[329] = (N3)? mem[329] :
                         (N0)? mem[899] : 1'b0;
  assign r_data_o[328] = (N3)? mem[328] :
                         (N0)? mem[898] : 1'b0;
  assign r_data_o[327] = (N3)? mem[327] :
                         (N0)? mem[897] : 1'b0;
  assign r_data_o[326] = (N3)? mem[326] :
                         (N0)? mem[896] : 1'b0;
  assign r_data_o[325] = (N3)? mem[325] :
                         (N0)? mem[895] : 1'b0;
  assign r_data_o[324] = (N3)? mem[324] :
                         (N0)? mem[894] : 1'b0;
  assign r_data_o[323] = (N3)? mem[323] :
                         (N0)? mem[893] : 1'b0;
  assign r_data_o[322] = (N3)? mem[322] :
                         (N0)? mem[892] : 1'b0;
  assign r_data_o[321] = (N3)? mem[321] :
                         (N0)? mem[891] : 1'b0;
  assign r_data_o[320] = (N3)? mem[320] :
                         (N0)? mem[890] : 1'b0;
  assign r_data_o[319] = (N3)? mem[319] :
                         (N0)? mem[889] : 1'b0;
  assign r_data_o[318] = (N3)? mem[318] :
                         (N0)? mem[888] : 1'b0;
  assign r_data_o[317] = (N3)? mem[317] :
                         (N0)? mem[887] : 1'b0;
  assign r_data_o[316] = (N3)? mem[316] :
                         (N0)? mem[886] : 1'b0;
  assign r_data_o[315] = (N3)? mem[315] :
                         (N0)? mem[885] : 1'b0;
  assign r_data_o[314] = (N3)? mem[314] :
                         (N0)? mem[884] : 1'b0;
  assign r_data_o[313] = (N3)? mem[313] :
                         (N0)? mem[883] : 1'b0;
  assign r_data_o[312] = (N3)? mem[312] :
                         (N0)? mem[882] : 1'b0;
  assign r_data_o[311] = (N3)? mem[311] :
                         (N0)? mem[881] : 1'b0;
  assign r_data_o[310] = (N3)? mem[310] :
                         (N0)? mem[880] : 1'b0;
  assign r_data_o[309] = (N3)? mem[309] :
                         (N0)? mem[879] : 1'b0;
  assign r_data_o[308] = (N3)? mem[308] :
                         (N0)? mem[878] : 1'b0;
  assign r_data_o[307] = (N3)? mem[307] :
                         (N0)? mem[877] : 1'b0;
  assign r_data_o[306] = (N3)? mem[306] :
                         (N0)? mem[876] : 1'b0;
  assign r_data_o[305] = (N3)? mem[305] :
                         (N0)? mem[875] : 1'b0;
  assign r_data_o[304] = (N3)? mem[304] :
                         (N0)? mem[874] : 1'b0;
  assign r_data_o[303] = (N3)? mem[303] :
                         (N0)? mem[873] : 1'b0;
  assign r_data_o[302] = (N3)? mem[302] :
                         (N0)? mem[872] : 1'b0;
  assign r_data_o[301] = (N3)? mem[301] :
                         (N0)? mem[871] : 1'b0;
  assign r_data_o[300] = (N3)? mem[300] :
                         (N0)? mem[870] : 1'b0;
  assign r_data_o[299] = (N3)? mem[299] :
                         (N0)? mem[869] : 1'b0;
  assign r_data_o[298] = (N3)? mem[298] :
                         (N0)? mem[868] : 1'b0;
  assign r_data_o[297] = (N3)? mem[297] :
                         (N0)? mem[867] : 1'b0;
  assign r_data_o[296] = (N3)? mem[296] :
                         (N0)? mem[866] : 1'b0;
  assign r_data_o[295] = (N3)? mem[295] :
                         (N0)? mem[865] : 1'b0;
  assign r_data_o[294] = (N3)? mem[294] :
                         (N0)? mem[864] : 1'b0;
  assign r_data_o[293] = (N3)? mem[293] :
                         (N0)? mem[863] : 1'b0;
  assign r_data_o[292] = (N3)? mem[292] :
                         (N0)? mem[862] : 1'b0;
  assign r_data_o[291] = (N3)? mem[291] :
                         (N0)? mem[861] : 1'b0;
  assign r_data_o[290] = (N3)? mem[290] :
                         (N0)? mem[860] : 1'b0;
  assign r_data_o[289] = (N3)? mem[289] :
                         (N0)? mem[859] : 1'b0;
  assign r_data_o[288] = (N3)? mem[288] :
                         (N0)? mem[858] : 1'b0;
  assign r_data_o[287] = (N3)? mem[287] :
                         (N0)? mem[857] : 1'b0;
  assign r_data_o[286] = (N3)? mem[286] :
                         (N0)? mem[856] : 1'b0;
  assign r_data_o[285] = (N3)? mem[285] :
                         (N0)? mem[855] : 1'b0;
  assign r_data_o[284] = (N3)? mem[284] :
                         (N0)? mem[854] : 1'b0;
  assign r_data_o[283] = (N3)? mem[283] :
                         (N0)? mem[853] : 1'b0;
  assign r_data_o[282] = (N3)? mem[282] :
                         (N0)? mem[852] : 1'b0;
  assign r_data_o[281] = (N3)? mem[281] :
                         (N0)? mem[851] : 1'b0;
  assign r_data_o[280] = (N3)? mem[280] :
                         (N0)? mem[850] : 1'b0;
  assign r_data_o[279] = (N3)? mem[279] :
                         (N0)? mem[849] : 1'b0;
  assign r_data_o[278] = (N3)? mem[278] :
                         (N0)? mem[848] : 1'b0;
  assign r_data_o[277] = (N3)? mem[277] :
                         (N0)? mem[847] : 1'b0;
  assign r_data_o[276] = (N3)? mem[276] :
                         (N0)? mem[846] : 1'b0;
  assign r_data_o[275] = (N3)? mem[275] :
                         (N0)? mem[845] : 1'b0;
  assign r_data_o[274] = (N3)? mem[274] :
                         (N0)? mem[844] : 1'b0;
  assign r_data_o[273] = (N3)? mem[273] :
                         (N0)? mem[843] : 1'b0;
  assign r_data_o[272] = (N3)? mem[272] :
                         (N0)? mem[842] : 1'b0;
  assign r_data_o[271] = (N3)? mem[271] :
                         (N0)? mem[841] : 1'b0;
  assign r_data_o[270] = (N3)? mem[270] :
                         (N0)? mem[840] : 1'b0;
  assign r_data_o[269] = (N3)? mem[269] :
                         (N0)? mem[839] : 1'b0;
  assign r_data_o[268] = (N3)? mem[268] :
                         (N0)? mem[838] : 1'b0;
  assign r_data_o[267] = (N3)? mem[267] :
                         (N0)? mem[837] : 1'b0;
  assign r_data_o[266] = (N3)? mem[266] :
                         (N0)? mem[836] : 1'b0;
  assign r_data_o[265] = (N3)? mem[265] :
                         (N0)? mem[835] : 1'b0;
  assign r_data_o[264] = (N3)? mem[264] :
                         (N0)? mem[834] : 1'b0;
  assign r_data_o[263] = (N3)? mem[263] :
                         (N0)? mem[833] : 1'b0;
  assign r_data_o[262] = (N3)? mem[262] :
                         (N0)? mem[832] : 1'b0;
  assign r_data_o[261] = (N3)? mem[261] :
                         (N0)? mem[831] : 1'b0;
  assign r_data_o[260] = (N3)? mem[260] :
                         (N0)? mem[830] : 1'b0;
  assign r_data_o[259] = (N3)? mem[259] :
                         (N0)? mem[829] : 1'b0;
  assign r_data_o[258] = (N3)? mem[258] :
                         (N0)? mem[828] : 1'b0;
  assign r_data_o[257] = (N3)? mem[257] :
                         (N0)? mem[827] : 1'b0;
  assign r_data_o[256] = (N3)? mem[256] :
                         (N0)? mem[826] : 1'b0;
  assign r_data_o[255] = (N3)? mem[255] :
                         (N0)? mem[825] : 1'b0;
  assign r_data_o[254] = (N3)? mem[254] :
                         (N0)? mem[824] : 1'b0;
  assign r_data_o[253] = (N3)? mem[253] :
                         (N0)? mem[823] : 1'b0;
  assign r_data_o[252] = (N3)? mem[252] :
                         (N0)? mem[822] : 1'b0;
  assign r_data_o[251] = (N3)? mem[251] :
                         (N0)? mem[821] : 1'b0;
  assign r_data_o[250] = (N3)? mem[250] :
                         (N0)? mem[820] : 1'b0;
  assign r_data_o[249] = (N3)? mem[249] :
                         (N0)? mem[819] : 1'b0;
  assign r_data_o[248] = (N3)? mem[248] :
                         (N0)? mem[818] : 1'b0;
  assign r_data_o[247] = (N3)? mem[247] :
                         (N0)? mem[817] : 1'b0;
  assign r_data_o[246] = (N3)? mem[246] :
                         (N0)? mem[816] : 1'b0;
  assign r_data_o[245] = (N3)? mem[245] :
                         (N0)? mem[815] : 1'b0;
  assign r_data_o[244] = (N3)? mem[244] :
                         (N0)? mem[814] : 1'b0;
  assign r_data_o[243] = (N3)? mem[243] :
                         (N0)? mem[813] : 1'b0;
  assign r_data_o[242] = (N3)? mem[242] :
                         (N0)? mem[812] : 1'b0;
  assign r_data_o[241] = (N3)? mem[241] :
                         (N0)? mem[811] : 1'b0;
  assign r_data_o[240] = (N3)? mem[240] :
                         (N0)? mem[810] : 1'b0;
  assign r_data_o[239] = (N3)? mem[239] :
                         (N0)? mem[809] : 1'b0;
  assign r_data_o[238] = (N3)? mem[238] :
                         (N0)? mem[808] : 1'b0;
  assign r_data_o[237] = (N3)? mem[237] :
                         (N0)? mem[807] : 1'b0;
  assign r_data_o[236] = (N3)? mem[236] :
                         (N0)? mem[806] : 1'b0;
  assign r_data_o[235] = (N3)? mem[235] :
                         (N0)? mem[805] : 1'b0;
  assign r_data_o[234] = (N3)? mem[234] :
                         (N0)? mem[804] : 1'b0;
  assign r_data_o[233] = (N3)? mem[233] :
                         (N0)? mem[803] : 1'b0;
  assign r_data_o[232] = (N3)? mem[232] :
                         (N0)? mem[802] : 1'b0;
  assign r_data_o[231] = (N3)? mem[231] :
                         (N0)? mem[801] : 1'b0;
  assign r_data_o[230] = (N3)? mem[230] :
                         (N0)? mem[800] : 1'b0;
  assign r_data_o[229] = (N3)? mem[229] :
                         (N0)? mem[799] : 1'b0;
  assign r_data_o[228] = (N3)? mem[228] :
                         (N0)? mem[798] : 1'b0;
  assign r_data_o[227] = (N3)? mem[227] :
                         (N0)? mem[797] : 1'b0;
  assign r_data_o[226] = (N3)? mem[226] :
                         (N0)? mem[796] : 1'b0;
  assign r_data_o[225] = (N3)? mem[225] :
                         (N0)? mem[795] : 1'b0;
  assign r_data_o[224] = (N3)? mem[224] :
                         (N0)? mem[794] : 1'b0;
  assign r_data_o[223] = (N3)? mem[223] :
                         (N0)? mem[793] : 1'b0;
  assign r_data_o[222] = (N3)? mem[222] :
                         (N0)? mem[792] : 1'b0;
  assign r_data_o[221] = (N3)? mem[221] :
                         (N0)? mem[791] : 1'b0;
  assign r_data_o[220] = (N3)? mem[220] :
                         (N0)? mem[790] : 1'b0;
  assign r_data_o[219] = (N3)? mem[219] :
                         (N0)? mem[789] : 1'b0;
  assign r_data_o[218] = (N3)? mem[218] :
                         (N0)? mem[788] : 1'b0;
  assign r_data_o[217] = (N3)? mem[217] :
                         (N0)? mem[787] : 1'b0;
  assign r_data_o[216] = (N3)? mem[216] :
                         (N0)? mem[786] : 1'b0;
  assign r_data_o[215] = (N3)? mem[215] :
                         (N0)? mem[785] : 1'b0;
  assign r_data_o[214] = (N3)? mem[214] :
                         (N0)? mem[784] : 1'b0;
  assign r_data_o[213] = (N3)? mem[213] :
                         (N0)? mem[783] : 1'b0;
  assign r_data_o[212] = (N3)? mem[212] :
                         (N0)? mem[782] : 1'b0;
  assign r_data_o[211] = (N3)? mem[211] :
                         (N0)? mem[781] : 1'b0;
  assign r_data_o[210] = (N3)? mem[210] :
                         (N0)? mem[780] : 1'b0;
  assign r_data_o[209] = (N3)? mem[209] :
                         (N0)? mem[779] : 1'b0;
  assign r_data_o[208] = (N3)? mem[208] :
                         (N0)? mem[778] : 1'b0;
  assign r_data_o[207] = (N3)? mem[207] :
                         (N0)? mem[777] : 1'b0;
  assign r_data_o[206] = (N3)? mem[206] :
                         (N0)? mem[776] : 1'b0;
  assign r_data_o[205] = (N3)? mem[205] :
                         (N0)? mem[775] : 1'b0;
  assign r_data_o[204] = (N3)? mem[204] :
                         (N0)? mem[774] : 1'b0;
  assign r_data_o[203] = (N3)? mem[203] :
                         (N0)? mem[773] : 1'b0;
  assign r_data_o[202] = (N3)? mem[202] :
                         (N0)? mem[772] : 1'b0;
  assign r_data_o[201] = (N3)? mem[201] :
                         (N0)? mem[771] : 1'b0;
  assign r_data_o[200] = (N3)? mem[200] :
                         (N0)? mem[770] : 1'b0;
  assign r_data_o[199] = (N3)? mem[199] :
                         (N0)? mem[769] : 1'b0;
  assign r_data_o[198] = (N3)? mem[198] :
                         (N0)? mem[768] : 1'b0;
  assign r_data_o[197] = (N3)? mem[197] :
                         (N0)? mem[767] : 1'b0;
  assign r_data_o[196] = (N3)? mem[196] :
                         (N0)? mem[766] : 1'b0;
  assign r_data_o[195] = (N3)? mem[195] :
                         (N0)? mem[765] : 1'b0;
  assign r_data_o[194] = (N3)? mem[194] :
                         (N0)? mem[764] : 1'b0;
  assign r_data_o[193] = (N3)? mem[193] :
                         (N0)? mem[763] : 1'b0;
  assign r_data_o[192] = (N3)? mem[192] :
                         (N0)? mem[762] : 1'b0;
  assign r_data_o[191] = (N3)? mem[191] :
                         (N0)? mem[761] : 1'b0;
  assign r_data_o[190] = (N3)? mem[190] :
                         (N0)? mem[760] : 1'b0;
  assign r_data_o[189] = (N3)? mem[189] :
                         (N0)? mem[759] : 1'b0;
  assign r_data_o[188] = (N3)? mem[188] :
                         (N0)? mem[758] : 1'b0;
  assign r_data_o[187] = (N3)? mem[187] :
                         (N0)? mem[757] : 1'b0;
  assign r_data_o[186] = (N3)? mem[186] :
                         (N0)? mem[756] : 1'b0;
  assign r_data_o[185] = (N3)? mem[185] :
                         (N0)? mem[755] : 1'b0;
  assign r_data_o[184] = (N3)? mem[184] :
                         (N0)? mem[754] : 1'b0;
  assign r_data_o[183] = (N3)? mem[183] :
                         (N0)? mem[753] : 1'b0;
  assign r_data_o[182] = (N3)? mem[182] :
                         (N0)? mem[752] : 1'b0;
  assign r_data_o[181] = (N3)? mem[181] :
                         (N0)? mem[751] : 1'b0;
  assign r_data_o[180] = (N3)? mem[180] :
                         (N0)? mem[750] : 1'b0;
  assign r_data_o[179] = (N3)? mem[179] :
                         (N0)? mem[749] : 1'b0;
  assign r_data_o[178] = (N3)? mem[178] :
                         (N0)? mem[748] : 1'b0;
  assign r_data_o[177] = (N3)? mem[177] :
                         (N0)? mem[747] : 1'b0;
  assign r_data_o[176] = (N3)? mem[176] :
                         (N0)? mem[746] : 1'b0;
  assign r_data_o[175] = (N3)? mem[175] :
                         (N0)? mem[745] : 1'b0;
  assign r_data_o[174] = (N3)? mem[174] :
                         (N0)? mem[744] : 1'b0;
  assign r_data_o[173] = (N3)? mem[173] :
                         (N0)? mem[743] : 1'b0;
  assign r_data_o[172] = (N3)? mem[172] :
                         (N0)? mem[742] : 1'b0;
  assign r_data_o[171] = (N3)? mem[171] :
                         (N0)? mem[741] : 1'b0;
  assign r_data_o[170] = (N3)? mem[170] :
                         (N0)? mem[740] : 1'b0;
  assign r_data_o[169] = (N3)? mem[169] :
                         (N0)? mem[739] : 1'b0;
  assign r_data_o[168] = (N3)? mem[168] :
                         (N0)? mem[738] : 1'b0;
  assign r_data_o[167] = (N3)? mem[167] :
                         (N0)? mem[737] : 1'b0;
  assign r_data_o[166] = (N3)? mem[166] :
                         (N0)? mem[736] : 1'b0;
  assign r_data_o[165] = (N3)? mem[165] :
                         (N0)? mem[735] : 1'b0;
  assign r_data_o[164] = (N3)? mem[164] :
                         (N0)? mem[734] : 1'b0;
  assign r_data_o[163] = (N3)? mem[163] :
                         (N0)? mem[733] : 1'b0;
  assign r_data_o[162] = (N3)? mem[162] :
                         (N0)? mem[732] : 1'b0;
  assign r_data_o[161] = (N3)? mem[161] :
                         (N0)? mem[731] : 1'b0;
  assign r_data_o[160] = (N3)? mem[160] :
                         (N0)? mem[730] : 1'b0;
  assign r_data_o[159] = (N3)? mem[159] :
                         (N0)? mem[729] : 1'b0;
  assign r_data_o[158] = (N3)? mem[158] :
                         (N0)? mem[728] : 1'b0;
  assign r_data_o[157] = (N3)? mem[157] :
                         (N0)? mem[727] : 1'b0;
  assign r_data_o[156] = (N3)? mem[156] :
                         (N0)? mem[726] : 1'b0;
  assign r_data_o[155] = (N3)? mem[155] :
                         (N0)? mem[725] : 1'b0;
  assign r_data_o[154] = (N3)? mem[154] :
                         (N0)? mem[724] : 1'b0;
  assign r_data_o[153] = (N3)? mem[153] :
                         (N0)? mem[723] : 1'b0;
  assign r_data_o[152] = (N3)? mem[152] :
                         (N0)? mem[722] : 1'b0;
  assign r_data_o[151] = (N3)? mem[151] :
                         (N0)? mem[721] : 1'b0;
  assign r_data_o[150] = (N3)? mem[150] :
                         (N0)? mem[720] : 1'b0;
  assign r_data_o[149] = (N3)? mem[149] :
                         (N0)? mem[719] : 1'b0;
  assign r_data_o[148] = (N3)? mem[148] :
                         (N0)? mem[718] : 1'b0;
  assign r_data_o[147] = (N3)? mem[147] :
                         (N0)? mem[717] : 1'b0;
  assign r_data_o[146] = (N3)? mem[146] :
                         (N0)? mem[716] : 1'b0;
  assign r_data_o[145] = (N3)? mem[145] :
                         (N0)? mem[715] : 1'b0;
  assign r_data_o[144] = (N3)? mem[144] :
                         (N0)? mem[714] : 1'b0;
  assign r_data_o[143] = (N3)? mem[143] :
                         (N0)? mem[713] : 1'b0;
  assign r_data_o[142] = (N3)? mem[142] :
                         (N0)? mem[712] : 1'b0;
  assign r_data_o[141] = (N3)? mem[141] :
                         (N0)? mem[711] : 1'b0;
  assign r_data_o[140] = (N3)? mem[140] :
                         (N0)? mem[710] : 1'b0;
  assign r_data_o[139] = (N3)? mem[139] :
                         (N0)? mem[709] : 1'b0;
  assign r_data_o[138] = (N3)? mem[138] :
                         (N0)? mem[708] : 1'b0;
  assign r_data_o[137] = (N3)? mem[137] :
                         (N0)? mem[707] : 1'b0;
  assign r_data_o[136] = (N3)? mem[136] :
                         (N0)? mem[706] : 1'b0;
  assign r_data_o[135] = (N3)? mem[135] :
                         (N0)? mem[705] : 1'b0;
  assign r_data_o[134] = (N3)? mem[134] :
                         (N0)? mem[704] : 1'b0;
  assign r_data_o[133] = (N3)? mem[133] :
                         (N0)? mem[703] : 1'b0;
  assign r_data_o[132] = (N3)? mem[132] :
                         (N0)? mem[702] : 1'b0;
  assign r_data_o[131] = (N3)? mem[131] :
                         (N0)? mem[701] : 1'b0;
  assign r_data_o[130] = (N3)? mem[130] :
                         (N0)? mem[700] : 1'b0;
  assign r_data_o[129] = (N3)? mem[129] :
                         (N0)? mem[699] : 1'b0;
  assign r_data_o[128] = (N3)? mem[128] :
                         (N0)? mem[698] : 1'b0;
  assign r_data_o[127] = (N3)? mem[127] :
                         (N0)? mem[697] : 1'b0;
  assign r_data_o[126] = (N3)? mem[126] :
                         (N0)? mem[696] : 1'b0;
  assign r_data_o[125] = (N3)? mem[125] :
                         (N0)? mem[695] : 1'b0;
  assign r_data_o[124] = (N3)? mem[124] :
                         (N0)? mem[694] : 1'b0;
  assign r_data_o[123] = (N3)? mem[123] :
                         (N0)? mem[693] : 1'b0;
  assign r_data_o[122] = (N3)? mem[122] :
                         (N0)? mem[692] : 1'b0;
  assign r_data_o[121] = (N3)? mem[121] :
                         (N0)? mem[691] : 1'b0;
  assign r_data_o[120] = (N3)? mem[120] :
                         (N0)? mem[690] : 1'b0;
  assign r_data_o[119] = (N3)? mem[119] :
                         (N0)? mem[689] : 1'b0;
  assign r_data_o[118] = (N3)? mem[118] :
                         (N0)? mem[688] : 1'b0;
  assign r_data_o[117] = (N3)? mem[117] :
                         (N0)? mem[687] : 1'b0;
  assign r_data_o[116] = (N3)? mem[116] :
                         (N0)? mem[686] : 1'b0;
  assign r_data_o[115] = (N3)? mem[115] :
                         (N0)? mem[685] : 1'b0;
  assign r_data_o[114] = (N3)? mem[114] :
                         (N0)? mem[684] : 1'b0;
  assign r_data_o[113] = (N3)? mem[113] :
                         (N0)? mem[683] : 1'b0;
  assign r_data_o[112] = (N3)? mem[112] :
                         (N0)? mem[682] : 1'b0;
  assign r_data_o[111] = (N3)? mem[111] :
                         (N0)? mem[681] : 1'b0;
  assign r_data_o[110] = (N3)? mem[110] :
                         (N0)? mem[680] : 1'b0;
  assign r_data_o[109] = (N3)? mem[109] :
                         (N0)? mem[679] : 1'b0;
  assign r_data_o[108] = (N3)? mem[108] :
                         (N0)? mem[678] : 1'b0;
  assign r_data_o[107] = (N3)? mem[107] :
                         (N0)? mem[677] : 1'b0;
  assign r_data_o[106] = (N3)? mem[106] :
                         (N0)? mem[676] : 1'b0;
  assign r_data_o[105] = (N3)? mem[105] :
                         (N0)? mem[675] : 1'b0;
  assign r_data_o[104] = (N3)? mem[104] :
                         (N0)? mem[674] : 1'b0;
  assign r_data_o[103] = (N3)? mem[103] :
                         (N0)? mem[673] : 1'b0;
  assign r_data_o[102] = (N3)? mem[102] :
                         (N0)? mem[672] : 1'b0;
  assign r_data_o[101] = (N3)? mem[101] :
                         (N0)? mem[671] : 1'b0;
  assign r_data_o[100] = (N3)? mem[100] :
                         (N0)? mem[670] : 1'b0;
  assign r_data_o[99] = (N3)? mem[99] :
                        (N0)? mem[669] : 1'b0;
  assign r_data_o[98] = (N3)? mem[98] :
                        (N0)? mem[668] : 1'b0;
  assign r_data_o[97] = (N3)? mem[97] :
                        (N0)? mem[667] : 1'b0;
  assign r_data_o[96] = (N3)? mem[96] :
                        (N0)? mem[666] : 1'b0;
  assign r_data_o[95] = (N3)? mem[95] :
                        (N0)? mem[665] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] :
                        (N0)? mem[664] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] :
                        (N0)? mem[663] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] :
                        (N0)? mem[662] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] :
                        (N0)? mem[661] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] :
                        (N0)? mem[660] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] :
                        (N0)? mem[659] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] :
                        (N0)? mem[658] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] :
                        (N0)? mem[657] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] :
                        (N0)? mem[656] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] :
                        (N0)? mem[655] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] :
                        (N0)? mem[654] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] :
                        (N0)? mem[653] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] :
                        (N0)? mem[652] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] :
                        (N0)? mem[651] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] :
                        (N0)? mem[650] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] :
                        (N0)? mem[649] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] :
                        (N0)? mem[648] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] :
                        (N0)? mem[647] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] :
                        (N0)? mem[646] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] :
                        (N0)? mem[645] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] :
                        (N0)? mem[644] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] :
                        (N0)? mem[643] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] :
                        (N0)? mem[642] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] :
                        (N0)? mem[641] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] :
                        (N0)? mem[640] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] :
                        (N0)? mem[639] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] :
                        (N0)? mem[638] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] :
                        (N0)? mem[637] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] :
                        (N0)? mem[636] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] :
                        (N0)? mem[635] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] :
                        (N0)? mem[634] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] :
                        (N0)? mem[633] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] :
                        (N0)? mem[632] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] :
                        (N0)? mem[631] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] :
                        (N0)? mem[630] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] :
                        (N0)? mem[629] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] :
                        (N0)? mem[628] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] :
                        (N0)? mem[627] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] :
                        (N0)? mem[626] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] :
                        (N0)? mem[625] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] :
                        (N0)? mem[624] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] :
                        (N0)? mem[623] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] :
                        (N0)? mem[622] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] :
                        (N0)? mem[621] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] :
                        (N0)? mem[620] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] :
                        (N0)? mem[619] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] :
                        (N0)? mem[618] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] :
                        (N0)? mem[617] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] :
                        (N0)? mem[616] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] :
                        (N0)? mem[615] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] :
                        (N0)? mem[614] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] :
                        (N0)? mem[613] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] :
                        (N0)? mem[612] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] :
                        (N0)? mem[611] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] :
                        (N0)? mem[610] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] :
                        (N0)? mem[609] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] :
                        (N0)? mem[608] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] :
                        (N0)? mem[607] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] :
                        (N0)? mem[606] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] :
                        (N0)? mem[605] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] :
                        (N0)? mem[604] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] :
                        (N0)? mem[603] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] :
                        (N0)? mem[602] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] :
                        (N0)? mem[601] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] :
                        (N0)? mem[600] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] :
                        (N0)? mem[599] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] :
                        (N0)? mem[598] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] :
                        (N0)? mem[597] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] :
                        (N0)? mem[596] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] :
                        (N0)? mem[595] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] :
                        (N0)? mem[594] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] :
                        (N0)? mem[593] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] :
                        (N0)? mem[592] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] :
                        (N0)? mem[591] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] :
                        (N0)? mem[590] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] :
                        (N0)? mem[589] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] :
                        (N0)? mem[588] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] :
                        (N0)? mem[587] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] :
                        (N0)? mem[586] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] :
                        (N0)? mem[585] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] :
                        (N0)? mem[584] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] :
                        (N0)? mem[583] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] :
                        (N0)? mem[582] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] :
                        (N0)? mem[581] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] :
                        (N0)? mem[580] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] :
                       (N0)? mem[579] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] :
                       (N0)? mem[578] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] :
                       (N0)? mem[577] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] :
                       (N0)? mem[576] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] :
                       (N0)? mem[575] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] :
                       (N0)? mem[574] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] :
                       (N0)? mem[573] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] :
                       (N0)? mem[572] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] :
                       (N0)? mem[571] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] :
                       (N0)? mem[570] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], N5, N5, N5, N5, N5, N5 } :
                                                                       (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N13) begin
      { mem[1139:1041], mem[570:570] } <= { w_data_i[569:471], w_data_i[0:0] };
    end
    if(N14) begin
      { mem[1040:942], mem[571:571] } <= { w_data_i[470:372], w_data_i[1:1] };
    end
    if(N15) begin
      { mem[941:843], mem[572:572] } <= { w_data_i[371:273], w_data_i[2:2] };
    end
    if(N16) begin
      { mem[842:744], mem[573:573] } <= { w_data_i[272:174], w_data_i[3:3] };
    end
    if(N17) begin
      { mem[743:645], mem[574:574] } <= { w_data_i[173:75], w_data_i[4:4] };
    end
    if(N18) begin
      { mem[644:575] } <= { w_data_i[74:5] };
    end
    if(N7) begin
      { mem[569:471], mem[0:0] } <= { w_data_i[569:471], w_data_i[0:0] };
    end
    if(N8) begin
      { mem[470:372], mem[1:1] } <= { w_data_i[470:372], w_data_i[1:1] };
    end
    if(N9) begin
      { mem[371:273], mem[2:2] } <= { w_data_i[371:273], w_data_i[2:2] };
    end
    if(N10) begin
      { mem[272:174], mem[3:3] } <= { w_data_i[272:174], w_data_i[3:3] };
    end
    if(N11) begin
      { mem[173:75], mem[4:4] } <= { w_data_i[173:75], w_data_i[4:4] };
    end
    if(N12) begin
      { mem[74:5] } <= { w_data_i[74:5] };
    end
  end


endmodule



module bsg_mem_1r1w_width_p570_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [569:0] w_data_i;
  input [0:0] r_addr_i;
  output [569:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [569:0] r_data_o;

  bsg_mem_p570
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p570
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [569:0] data_i;
  output [569:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [569:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p570_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 :
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 :
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 :
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 :
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 :
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 :
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end
    if(N9) begin
      tail_r <= N10;
    end
    if(N11) begin
      head_r <= N12;
    end
  end


endmodule



module bsg_mem_1rw_sync_width_p96_els_p256
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_i,
  data_o
);

  input [95:0] data_i;
  input [7:0] addr_i;
  output [95:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [95:0] data_o;

  hard_mem_1rw_d256_w96_wrapper
  macro_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bp_cce_pc_inst_ram_els_p256_harden_p0
(
  clk_i,
  reset_i,
  alu_branch_res_i,
  pc_stall_i,
  pc_branch_target_i,
  inst_o,
  inst_v_o,
  boot_rom_addr_o,
  boot_rom_data_i
);

  input [7:0] pc_branch_target_i;
  output [95:0] inst_o;
  output [7:0] boot_rom_addr_o;
  input [95:0] boot_rom_data_i;
  input clk_i;
  input reset_i;
  input alu_branch_res_i;
  input pc_stall_i;
  output inst_v_o;
  wire [95:0] inst_o,ram_data_i_r_n;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,ram_w_r_n,inst_v_r_n,N9,N10,N11,N12,N13,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,
  N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,
  N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,
  N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,
  N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,
  N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,
  N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,
  N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,
  N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211,N212;
  wire [7:0] ram_addr_i,ram_addr_r_n,boot_rom_addr_r_n,ex_pc_r_n;
  wire [1:0] pc_state_n;
  reg inst_v_o,ram_v_r,ram_w_r;
  reg [1:0] pc_state;
  reg [7:0] ram_addr_r,boot_rom_addr_o,ex_pc_r;
  reg [95:0] ram_data_i_r;

  bsg_mem_1rw_sync_width_p96_els_p256
  cce_inst_ram
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(ram_data_i_r),
    .addr_i(ram_addr_i),
    .v_i(ram_v_r),
    .w_i(ram_w_r),
    .data_o(inst_o)
  );

  assign N135 = N133 & N134;
  assign N136 = pc_state[1] | N134;
  assign N138 = N133 | pc_state[0];
  assign N140 = pc_state[1] & pc_state[0];
  assign N206 = boot_rom_addr_o[6] & boot_rom_addr_o[7];
  assign N207 = boot_rom_addr_o[5] & N206;
  assign N208 = boot_rom_addr_o[4] & N207;
  assign N209 = boot_rom_addr_o[3] & N208;
  assign N210 = boot_rom_addr_o[2] & N209;
  assign N211 = boot_rom_addr_o[1] & N210;
  assign N212 = boot_rom_addr_o[0] & N211;
  assign { N176, N175, N174, N173, N172, N171, N170, N169 } = ram_addr_r + 1'b1;
  assign { N148, N147, N146, N145, N144, N143, N142, N141 } = boot_rom_addr_o + 1'b1;
  assign { N168, N167, N166, N165, N164, N163, N162, N161 } = pc_branch_target_i + 1'b1;
  assign { N156, N155, N154, N153, N152, N151, N150, N149 } = ram_addr_r + 1'b1;
  assign { N10, N9 } = (N0)? { 1'b0, 1'b0 } :
                       (N1)? pc_state_n : 1'b0;
  assign N0 = N8;
  assign N1 = N7;
  assign N11 = (N0)? 1'b0 :
               (N1)? ram_w_r_n : 1'b0;
  assign { N19, N18, N17, N16, N15, N14, N13, N12 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                      (N1)? ram_addr_r_n : 1'b0;
  assign { N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1)? ram_data_i_r_n : 1'b0;
  assign { N123, N122, N121, N120, N119, N118, N117, N116 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                              (N1)? boot_rom_addr_r_n : 1'b0;
  assign { N131, N130, N129, N128, N127, N126, N125, N124 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                              (N1)? ex_pc_r_n : 1'b0;
  assign N132 = (N0)? 1'b0 :
                (N1)? inst_v_r_n : 1'b0;
  assign { N184, N183, N182, N181, N180, N179, N178, N177 } = (N202)? pc_branch_target_i :
                                                              (N159)? ram_addr_r : 1'b0;
  assign { N192, N191, N190, N189, N188, N187, N186, N185 } = (N202)? { N168, N167, N166, N165, N164, N163, N162, N161 } :
                                                              (N159)? { N176, N175, N174, N173, N172, N171, N170, N169 } : 1'b0;
  assign { N200, N199, N198, N197, N196, N195, N194, N193 } = (N2)? ex_pc_r :
                                                              (N202)? pc_branch_target_i :
                                                              (N159)? ram_addr_r : 1'b0;
  assign N2 = pc_stall_i;
  assign pc_state_n = (N3)? { 1'b0, N212 } :
                      (N4)? { 1'b1, 1'b0 } :
                      (N5)? { 1'b1, 1'b1 } :
                      (N6)? { 1'b1, 1'b1 } : 1'b0;
  assign N3 = N135;
  assign N4 = N137;
  assign N5 = N139;
  assign N6 = N140;
  assign ram_w_r_n = (N3)? 1'b1 :
                     (N4)? 1'b0 :
                     (N5)? 1'b0 :
                     (N6)? 1'b0 : 1'b0;
  assign ram_addr_r_n = (N3)? boot_rom_addr_o :
                        (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                        (N5)? { N156, N155, N154, N153, N152, N151, N150, N149 } :
                        (N6)? { N192, N191, N190, N189, N188, N187, N186, N185 } : 1'b0;
  assign ram_data_i_r_n = (N3)? boot_rom_data_i :
                          (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                          (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                          (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign ex_pc_r_n = (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                     (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                     (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                     (N6)? { N184, N183, N182, N181, N180, N179, N178, N177 } : 1'b0;
  assign inst_v_r_n = (N3)? 1'b0 :
                      (N4)? 1'b0 :
                      (N5)? 1'b0 :
                      (N6)? 1'b1 : 1'b0;
  assign boot_rom_addr_r_n = (N3)? { N148, N147, N146, N145, N144, N143, N142, N141 } :
                             (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                             (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                             (N6)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign ram_addr_i = (N3)? ram_addr_r :
                      (N4)? ram_addr_r :
                      (N5)? ram_addr_r :
                      (N6)? { N200, N199, N198, N197, N196, N195, N194, N193 } : 1'b0;
  assign N7 = ~reset_i;
  assign N8 = reset_i;
  assign N133 = ~pc_state[1];
  assign N134 = ~pc_state[0];
  assign N137 = ~N136;
  assign N139 = ~N138;
  assign N157 = N140;
  assign N158 = alu_branch_res_i | pc_stall_i;
  assign N159 = ~N158;
  assign N160 = N157 & N202;
  assign N201 = ~pc_stall_i;
  assign N202 = alu_branch_res_i & N201;
  assign N203 = N140 & N7;
  assign N204 = pc_stall_i & N203;
  assign N205 = ~N204;

  always @(posedge clk_i) begin
    if(1'b1) begin
      inst_v_o <= N132;
      { pc_state[1:0] } <= { N10, N9 };
      ram_v_r <= N7;
      ram_w_r <= N11;
      { ram_data_i_r[95:0] } <= { N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20 };
      { boot_rom_addr_o[7:0] } <= { N123, N122, N121, N120, N119, N118, N117, N116 };
    end
    if(N205) begin
      { ram_addr_r[7:0] } <= { N19, N18, N17, N16, N15, N14, N13, N12 };
      { ex_pc_r[7:0] } <= { N131, N130, N129, N128, N127, N126, N125, N124 };
    end
  end


endmodule



module bp_cce_inst_decode_inst_width_p96_inst_addr_width_p8
(
  clk_i,
  reset_i,
  inst_i,
  inst_v_i,
  lce_req_v_i,
  lce_resp_v_i,
  lce_data_resp_v_i,
  mem_resp_v_i,
  mem_data_resp_v_i,
  pending_v_i,
  lce_cmd_ready_i,
  lce_data_cmd_ready_i,
  mem_cmd_ready_i,
  mem_data_cmd_ready_i,
  decoded_inst_o,
  decoded_inst_v_o,
  pc_stall_o,
  pc_branch_target_o
);

  input [95:0] inst_i;
  output [127:0] decoded_inst_o;
  output [7:0] pc_branch_target_o;
  input clk_i;
  input reset_i;
  input inst_v_i;
  input lce_req_v_i;
  input lce_resp_v_i;
  input lce_data_resp_v_i;
  input mem_resp_v_i;
  input mem_data_resp_v_i;
  input pending_v_i;
  input lce_cmd_ready_i;
  input lce_data_cmd_ready_i;
  input mem_cmd_ready_i;
  input mem_data_cmd_ready_i;
  output decoded_inst_v_o;
  output pc_stall_o;
  wire [127:0] decoded_inst_o;
  wire [7:0] pc_branch_target_o;
  wire decoded_inst_v_o,pc_stall_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,pushq_op,
  popq_op,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,
  N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,wfq_op,stall_op,wfq_q_ready,N42,N43,
  N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,
  N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,
  N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,
  N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,
  N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,
  N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,
  N151,N152,N153,N154,N155;
  assign N44 = N102 & N99;
  assign N45 = inst_i[63] | N99;
  assign N47 = N102 | inst_i[62];
  assign N49 = inst_i[63] & inst_i[62];
  assign N57 = inst_i[94] | inst_i[95];
  assign N58 = inst_i[93] | N57;
  assign N59 = ~N58;
  assign N60 = ~inst_i[93];
  assign N61 = N60 | N57;
  assign N62 = ~N61;
  assign N63 = ~inst_i[95];
  assign N64 = ~inst_i[94];
  assign N65 = N64 | N63;
  assign N66 = inst_i[93] | N65;
  assign N67 = ~N66;
  assign N68 = inst_i[91] | inst_i[92];
  assign N69 = inst_i[90] | N68;
  assign N70 = ~N69;
  assign N71 = inst_i[94] | N63;
  assign N72 = inst_i[93] | N71;
  assign N73 = ~N72;
  assign N74 = ~inst_i[90];
  assign N75 = N74 | N68;
  assign N76 = ~N75;
  assign N77 = ~inst_i[91];
  assign N78 = N77 | inst_i[92];
  assign N79 = inst_i[90] | N78;
  assign N80 = ~N79;
  assign N81 = inst_i[60] | inst_i[61];
  assign N82 = inst_i[59] | N81;
  assign N83 = ~N82;
  assign N84 = ~inst_i[60];
  assign N85 = N84 | inst_i[61];
  assign N86 = inst_i[59] | N85;
  assign N87 = ~N86;
  assign N88 = ~inst_i[61];
  assign N89 = inst_i[60] | N88;
  assign N90 = inst_i[59] | N89;
  assign N91 = ~N90;
  assign N92 = ~inst_i[59];
  assign N93 = N92 | N89;
  assign N94 = ~N93;
  assign N95 = N92 | N81;
  assign N96 = ~N95;
  assign N97 = inst_i[62] | inst_i[63];
  assign N98 = ~N97;
  assign N99 = ~inst_i[62];
  assign N100 = N99 | inst_i[63];
  assign N101 = ~N100;
  assign N102 = ~inst_i[63];
  assign N103 = inst_i[62] | N102;
  assign N104 = ~N103;
  assign N105 = inst_i[62] & inst_i[63];
  assign N106 = ~inst_i[76];
  assign N107 = ~inst_i[75];
  assign N108 = inst_i[78] | inst_i[79];
  assign N109 = inst_i[77] | N108;
  assign N110 = N106 | N109;
  assign N111 = N107 | N110;
  assign N112 = ~N111;
  assign N113 = inst_i[75] | N110;
  assign N114 = ~N113;
  assign N115 = inst_i[76] | N109;
  assign N116 = N107 | N115;
  assign N117 = ~N116;
  assign N118 = inst_i[75] | N115;
  assign N119 = ~N118;
  assign N120 = N64 | inst_i[95];
  assign N121 = inst_i[93] | N120;
  assign N122 = ~N121;
  assign N123 = inst_i[94] & inst_i[95];
  assign N124 = inst_i[93] & N123;
  assign N125 = N60 | N71;
  assign N126 = ~N125;
  assign N127 = inst_i[91] & inst_i[92];
  assign N128 = inst_i[90] & N127;
  assign { N18, N17, N16 } = (N0)? inst_i[92:90] :
                             (N1)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N73;
  assign N1 = N72;
  assign { N21, N20, N19 } = (N2)? inst_i[92:90] :
                             (N3)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2 = N126;
  assign N3 = N125;
  assign decoded_inst_v_o = (N4)? 1'b0 :
                            (N14)? inst_v_i : 1'b0;
  assign N4 = N13;
  assign decoded_inst_o = (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                          (N14)? { inst_i[92:59], N15, inst_i[58:29], N18, N17, N16, N73, N21, N20, N19, N126, inst_i[28:20], inst_i[61:59], inst_i[19:19], N122, N59, N22, N23, N24, N25, N26, inst_i[18:13], N27, N28, N29, inst_i[12:0], N39, N40, N41, inst_i[12:12], N30, N31, N32, N33, N34, N35, N36, N37, N38 } : 1'b0;
  assign N54 = (N5)? N50 :
               (N6)? N51 :
               (N7)? N52 :
               (N8)? N53 : 1'b0;
  assign N5 = N44;
  assign N6 = N46;
  assign N7 = N48;
  assign N8 = N49;
  assign N55 = (N9)? N54 :
               (N10)? N42 : 1'b0;
  assign N9 = pushq_op;
  assign N10 = N43;
  assign pc_stall_o = (N11)? 1'b0 :
                      (N12)? N55 : 1'b0;
  assign N11 = reset_i;
  assign N12 = N56;
  assign pc_branch_target_o = (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                              (N12)? inst_i[66:59] : 1'b0;
  assign pushq_op = N124 & N76;
  assign popq_op = N124 & N80;
  assign N13 = reset_i | N129;
  assign N129 = ~inst_v_i;
  assign N14 = ~N13;
  assign N15 = N59 | N62;
  assign N22 = N112 & N130;
  assign N130 = N122 | N59;
  assign N23 = N114 & N131;
  assign N131 = N122 | N59;
  assign N24 = N117 & N132;
  assign N132 = N122 | N59;
  assign N25 = N119 & N133;
  assign N133 = N122 | N59;
  assign N26 = N135 | N25;
  assign N135 = N134 | N24;
  assign N134 = N22 | N23;
  assign N27 = N67 & N70;
  assign N28 = N73 & N76;
  assign N29 = N73 & N80;
  assign N30 = popq_op & N83;
  assign N31 = popq_op & N91;
  assign N32 = popq_op & N94;
  assign N33 = popq_op & N96;
  assign N34 = popq_op & N87;
  assign N35 = N136 & N98;
  assign N136 = lce_cmd_ready_i & pushq_op;
  assign N36 = pushq_op & N101;
  assign N37 = N137 & N104;
  assign N137 = mem_cmd_ready_i & pushq_op;
  assign N38 = N138 & N105;
  assign N138 = mem_data_cmd_ready_i & pushq_op;
  assign N39 = popq_op & N83;
  assign N40 = popq_op & N87;
  assign N41 = popq_op & N139;
  assign N139 = N83 | N87;
  assign wfq_op = N124 & N70;
  assign stall_op = N67 & N128;
  assign wfq_q_ready = N148 | N149;
  assign N148 = N146 | N147;
  assign N146 = N144 | N145;
  assign N144 = N142 | N143;
  assign N142 = N140 | N141;
  assign N140 = inst_i[64] & lce_req_v_i;
  assign N141 = inst_i[63] & lce_resp_v_i;
  assign N143 = inst_i[62] & lce_data_resp_v_i;
  assign N145 = inst_i[61] & mem_resp_v_i;
  assign N147 = inst_i[60] & mem_data_resp_v_i;
  assign N149 = inst_i[59] & pending_v_i;
  assign N42 = stall_op | N151;
  assign N151 = wfq_op & N150;
  assign N150 = ~wfq_q_ready;
  assign N43 = ~pushq_op;
  assign N46 = ~N45;
  assign N48 = ~N47;
  assign N50 = N42 | N152;
  assign N152 = ~lce_cmd_ready_i;
  assign N51 = N42 | N153;
  assign N153 = ~lce_data_cmd_ready_i;
  assign N52 = N42 | N154;
  assign N154 = ~mem_cmd_ready_i;
  assign N53 = N42 | N155;
  assign N155 = ~mem_data_cmd_ready_i;
  assign N56 = ~reset_i;

endmodule



module bp_cce_alu_width_p16
(
  v_i,
  opd_a_i,
  opd_b_i,
  alu_op_i,
  v_o,
  res_o,
  branch_res_o
);

  input [15:0] opd_a_i;
  input [15:0] opd_b_i;
  input [2:0] alu_op_i;
  output [15:0] res_o;
  input v_i;
  output v_o;
  output branch_res_o;
  wire [15:0] res_o;
  wire v_o,branch_res_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,v_i,equal,less,N11,N12,N13,
  N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,
  N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,
  N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,
  N94,N95,N96,N97,N98,N99,N100,N101;
  assign v_o = v_i;
  assign equal = opd_a_i == opd_b_i;
  assign less = opd_a_i < opd_b_i;
  assign N12 = alu_op_i[2] | N28;
  assign N13 = N12 | alu_op_i[0];
  assign N16 = N12 | N15;
  assign N18 = N27 | alu_op_i[1];
  assign N19 = N18 | alu_op_i[0];
  assign N21 = N18 | N15;
  assign N23 = alu_op_i[2] & alu_op_i[1];
  assign N24 = N23 & alu_op_i[0];
  assign N25 = N27 | N28;
  assign N26 = N25 | alu_op_i[0];
  assign N29 = N27 & N28;
  assign { N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37 } = opd_a_i + opd_b_i;
  assign { N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53 } = opd_a_i - opd_b_i;
  assign N33 = (N0)? equal :
               (N1)? N31 :
               (N2)? less :
               (N3)? N32 :
               (N4)? 1'b1 :
               (N5)? 1'b0 : 1'b0;
  assign N0 = N14;
  assign N1 = N17;
  assign N2 = N20;
  assign N3 = N22;
  assign N4 = N24;
  assign N5 = N30;
  assign branch_res_o = (N6)? N33 :
                        (N7)? 1'b0 : 1'b0;
  assign N6 = v_i;
  assign N7 = N11;
  assign { N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69 } = (N8)? { N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37 } :
                                                                                              (N9)? { N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53 } : 1'b0;
  assign N8 = N15;
  assign N9 = alu_op_i[0];
  assign { N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85 } = (N10)? { N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69 } :
                                                                                               (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = N29;
  assign res_o = (N6)? { N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85 } :
                 (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = ~v_i;
  assign N14 = ~N13;
  assign N15 = ~alu_op_i[0];
  assign N17 = ~N16;
  assign N20 = ~N19;
  assign N22 = ~N21;
  assign N27 = ~alu_op_i[2];
  assign N28 = ~alu_op_i[1];
  assign N30 = N101 | N29;
  assign N101 = ~N26;
  assign N31 = ~equal;
  assign N32 = less | equal;
  assign N34 = v_i;
  assign N35 = ~N29;
  assign N36 = N34 & N29;

endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p192_els_p64
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [191:0] data_i;
  input [5:0] addr_i;
  input [191:0] w_mask_i;
  output [191:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [191:0] data_o;

  hard_mem_1rw_bit_mask_d64_w96_wrapper
  macro_mem0
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[95:0]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i[95:0]),
    .w_i(w_i),
    .data_o(data_o[95:0])
  );


  hard_mem_1rw_bit_mask_d64_w96_wrapper
  macro_mem1
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[191:96]),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i[191:96]),
    .w_i(w_i),
    .data_o(data_o[191:96])
  );


endmodule



module bp_cce_dir_num_way_groups_p64_num_lce_p2_lce_assoc_p8_tag_width_p10_harden_p0
(
  clk_i,
  reset_i,
  way_group_i,
  lce_i,
  way_i,
  r_cmd_i,
  r_v_i,
  tag_i,
  coh_state_i,
  pending_i,
  w_cmd_i,
  w_v_i,
  pending_o,
  pending_v_o,
  tag_o,
  coh_state_o,
  entry_v_o,
  way_group_o,
  way_group_v_o
);

  input [5:0] way_group_i;
  input [0:0] lce_i;
  input [2:0] way_i;
  input [2:0] r_cmd_i;
  input [9:0] tag_i;
  input [1:0] coh_state_i;
  input [2:0] w_cmd_i;
  output [9:0] tag_o;
  output [1:0] coh_state_o;
  output [191:0] way_group_o;
  input clk_i;
  input reset_i;
  input r_v_i;
  input pending_i;
  input w_v_i;
  output pending_o;
  output pending_v_o;
  output entry_v_o;
  output way_group_v_o;
  wire [9:0] tag_o;
  wire [1:0] coh_state_o;
  wire [191:0] way_group_o,wg_ram_w_mask,wg_ram_w_data;
  wire pending_o,pending_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,pending_w_v,N32,N33,
  N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,
  N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,
  N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,
  N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,
  N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,
  N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,
  N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,
  N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,
  N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
  N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,wg_ram_r_v,wg_ram_w_v,wg_ram_v,N291,N292,N293,N294,N295,N296,
  N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,
  N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,
  N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,
  N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,
  N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,
  N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,
  N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
  N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,
  N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,
  N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,
  N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,
  N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,
  N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,
  N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,
  N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,
  N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,
  N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,
  N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,
  N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,
  N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,
  N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,
  N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,
  N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,
  N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,
  N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,
  N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,
  N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,
  N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,
  N745,N746,N747,N748,N749,N750,N751,N752,N754,N755,N756,N757,N758,N759,N760,N761,
  N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,
  N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,
  N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,
  N810,N811,N812,N813,N814,N815,N816,N817,N818;
  wire [5:0] wg_ram_addr;
  wire [95:0] tag_set;
  reg [63:0] pending_bits_r;
  reg entry_v_o,way_group_v_o;
  assign pending_o = (N227)? pending_bits_r[0] :
                     (N229)? pending_bits_r[1] :
                     (N231)? pending_bits_r[2] :
                     (N233)? pending_bits_r[3] :
                     (N235)? pending_bits_r[4] :
                     (N237)? pending_bits_r[5] :
                     (N239)? pending_bits_r[6] :
                     (N241)? pending_bits_r[7] :
                     (N243)? pending_bits_r[8] :
                     (N245)? pending_bits_r[9] :
                     (N247)? pending_bits_r[10] :
                     (N249)? pending_bits_r[11] :
                     (N251)? pending_bits_r[12] :
                     (N253)? pending_bits_r[13] :
                     (N255)? pending_bits_r[14] :
                     (N257)? pending_bits_r[15] :
                     (N259)? pending_bits_r[16] :
                     (N261)? pending_bits_r[17] :
                     (N263)? pending_bits_r[18] :
                     (N265)? pending_bits_r[19] :
                     (N267)? pending_bits_r[20] :
                     (N269)? pending_bits_r[21] :
                     (N271)? pending_bits_r[22] :
                     (N273)? pending_bits_r[23] :
                     (N275)? pending_bits_r[24] :
                     (N277)? pending_bits_r[25] :
                     (N279)? pending_bits_r[26] :
                     (N281)? pending_bits_r[27] :
                     (N283)? pending_bits_r[28] :
                     (N285)? pending_bits_r[29] :
                     (N287)? pending_bits_r[30] :
                     (N289)? pending_bits_r[31] :
                     (N228)? pending_bits_r[32] :
                     (N230)? pending_bits_r[33] :
                     (N232)? pending_bits_r[34] :
                     (N234)? pending_bits_r[35] :
                     (N236)? pending_bits_r[36] :
                     (N238)? pending_bits_r[37] :
                     (N240)? pending_bits_r[38] :
                     (N242)? pending_bits_r[39] :
                     (N244)? pending_bits_r[40] :
                     (N246)? pending_bits_r[41] :
                     (N248)? pending_bits_r[42] :
                     (N250)? pending_bits_r[43] :
                     (N252)? pending_bits_r[44] :
                     (N254)? pending_bits_r[45] :
                     (N256)? pending_bits_r[46] :
                     (N258)? pending_bits_r[47] :
                     (N260)? pending_bits_r[48] :
                     (N262)? pending_bits_r[49] :
                     (N264)? pending_bits_r[50] :
                     (N266)? pending_bits_r[51] :
                     (N268)? pending_bits_r[52] :
                     (N270)? pending_bits_r[53] :
                     (N272)? pending_bits_r[54] :
                     (N274)? pending_bits_r[55] :
                     (N276)? pending_bits_r[56] :
                     (N278)? pending_bits_r[57] :
                     (N280)? pending_bits_r[58] :
                     (N282)? pending_bits_r[59] :
                     (N284)? pending_bits_r[60] :
                     (N286)? pending_bits_r[61] :
                     (N288)? pending_bits_r[62] :
                     (N290)? pending_bits_r[63] : 1'b0;
  assign { N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } << { N318, N317, N316, N315, N314, N313, N312, N311, N310 };
  assign { N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } << { N534, N533, N532, N531, N530, N529, N528, N527, N526 };
  assign wg_ram_w_data = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tag_i, coh_state_i } << { N750, N749, N748, N747, N746, N745, N744, N743, N742 };

  bsg_mem_1rw_sync_mask_write_bit_width_p192_els_p64
  wg_ram
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(wg_ram_w_data),
    .addr_i(wg_ram_addr),
    .v_i(wg_ram_v),
    .w_mask_i(wg_ram_w_mask),
    .w_i(wg_ram_w_v),
    .data_o(way_group_o)
  );

  assign N762 = r_cmd_i[1] | r_cmd_i[2];
  assign N763 = r_cmd_i[0] | N762;
  assign N764 = ~N763;
  assign N765 = ~w_cmd_i[0];
  assign N766 = N765 | N784;
  assign N767 = ~N766;
  assign N768 = ~w_cmd_i[1];
  assign N769 = N768 | w_cmd_i[2];
  assign N770 = w_cmd_i[0] | N769;
  assign N771 = ~N770;
  assign N772 = ~r_cmd_i[1];
  assign N773 = N772 | r_cmd_i[2];
  assign N774 = r_cmd_i[0] | N773;
  assign N775 = ~N774;
  assign N776 = ~r_cmd_i[0];
  assign N777 = N776 | N762;
  assign N778 = ~N777;
  assign N779 = N765 | N784;
  assign N780 = ~N779;
  assign N781 = N768 | w_cmd_i[2];
  assign N782 = w_cmd_i[0] | N781;
  assign N783 = ~N782;
  assign N784 = w_cmd_i[1] | w_cmd_i[2];
  assign N785 = w_cmd_i[0] | N784;
  assign N786 = ~N785;
  assign { N302, N301, N300, N299, N298, N297, N296, N295 } = lce_i[0] * { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign { N309, N308, N307, N306, N305, N304, N303 } = way_i * { 1'b1, 1'b1, 1'b0, 1'b0 };
  assign { N518, N517, N516, N515, N514, N513, N512, N511 } = lce_i[0] * { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign { N525, N524, N523, N522, N521, N520, N519 } = way_i * { 1'b1, 1'b1, 1'b0, 1'b0 };
  assign { N734, N733, N732, N731, N730, N729, N728, N727 } = lce_i[0] * { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign { N741, N740, N739, N738, N737, N736, N735 } = way_i * { 1'b1, 1'b1, 1'b0, 1'b0 };
  assign { N318, N317, N316, N315, N314, N313, N312, N311, N310 } = { N302, N301, N300, N299, N298, N297, N296, N295 } + { N309, N308, N307, N306, N305, N304, N303 };
  assign { N534, N533, N532, N531, N530, N529, N528, N527, N526 } = { N518, N517, N516, N515, N514, N513, N512, N511 } + { N525, N524, N523, N522, N521, N520, N519 };
  assign { N750, N749, N748, N747, N746, N745, N744, N743, N742 } = { N734, N733, N732, N731, N730, N729, N728, N727 } + { N741, N740, N739, N738, N737, N736, N735 };
  assign N787 = ~way_group_i[5];
  assign N788 = way_group_i[3] & way_group_i[4];
  assign N789 = N0 & way_group_i[4];
  assign N0 = ~way_group_i[3];
  assign N790 = way_group_i[3] & N1;
  assign N1 = ~way_group_i[4];
  assign N791 = N2 & N3;
  assign N2 = ~way_group_i[3];
  assign N3 = ~way_group_i[4];
  assign N792 = way_group_i[5] & N788;
  assign N793 = way_group_i[5] & N789;
  assign N794 = way_group_i[5] & N790;
  assign N795 = way_group_i[5] & N791;
  assign N796 = N787 & N788;
  assign N797 = N787 & N789;
  assign N798 = N787 & N790;
  assign N799 = N787 & N791;
  assign N800 = ~way_group_i[2];
  assign N801 = way_group_i[0] & way_group_i[1];
  assign N802 = N4 & way_group_i[1];
  assign N4 = ~way_group_i[0];
  assign N803 = way_group_i[0] & N5;
  assign N5 = ~way_group_i[1];
  assign N804 = N6 & N7;
  assign N6 = ~way_group_i[0];
  assign N7 = ~way_group_i[1];
  assign N805 = way_group_i[2] & N801;
  assign N806 = way_group_i[2] & N802;
  assign N807 = way_group_i[2] & N803;
  assign N808 = way_group_i[2] & N804;
  assign N809 = N800 & N801;
  assign N810 = N800 & N802;
  assign N811 = N800 & N803;
  assign N812 = N800 & N804;
  assign N96 = N792 & N805;
  assign N95 = N792 & N806;
  assign N94 = N792 & N807;
  assign N93 = N792 & N808;
  assign N92 = N792 & N809;
  assign N91 = N792 & N810;
  assign N90 = N792 & N811;
  assign N89 = N792 & N812;
  assign N88 = N793 & N805;
  assign N87 = N793 & N806;
  assign N86 = N793 & N807;
  assign N85 = N793 & N808;
  assign N84 = N793 & N809;
  assign N83 = N793 & N810;
  assign N82 = N793 & N811;
  assign N81 = N793 & N812;
  assign N80 = N794 & N805;
  assign N79 = N794 & N806;
  assign N78 = N794 & N807;
  assign N77 = N794 & N808;
  assign N76 = N794 & N809;
  assign N75 = N794 & N810;
  assign N74 = N794 & N811;
  assign N73 = N794 & N812;
  assign N72 = N795 & N805;
  assign N71 = N795 & N806;
  assign N70 = N795 & N807;
  assign N69 = N795 & N808;
  assign N68 = N795 & N809;
  assign N67 = N795 & N810;
  assign N66 = N795 & N811;
  assign N65 = N795 & N812;
  assign N64 = N796 & N805;
  assign N63 = N796 & N806;
  assign N62 = N796 & N807;
  assign N61 = N796 & N808;
  assign N60 = N796 & N809;
  assign N59 = N796 & N810;
  assign N58 = N796 & N811;
  assign N57 = N796 & N812;
  assign N56 = N797 & N805;
  assign N55 = N797 & N806;
  assign N54 = N797 & N807;
  assign N53 = N797 & N808;
  assign N52 = N797 & N809;
  assign N51 = N797 & N810;
  assign N50 = N797 & N811;
  assign N49 = N797 & N812;
  assign N48 = N798 & N805;
  assign N47 = N798 & N806;
  assign N46 = N798 & N807;
  assign N45 = N798 & N808;
  assign N44 = N798 & N809;
  assign N43 = N798 & N810;
  assign N42 = N798 & N811;
  assign N41 = N798 & N812;
  assign N40 = N799 & N805;
  assign N39 = N799 & N806;
  assign N38 = N799 & N807;
  assign N37 = N799 & N808;
  assign N36 = N799 & N809;
  assign N35 = N799 & N810;
  assign N34 = N799 & N811;
  assign N33 = N799 & N812;
  assign N752 = ~lce_i[0];
  assign N813 = way_i[0] & way_i[1];
  assign N761 = N813 & way_i[2];
  assign N814 = N8 & way_i[1];
  assign N8 = ~way_i[0];
  assign N760 = N814 & way_i[2];
  assign N815 = way_i[0] & N9;
  assign N9 = ~way_i[1];
  assign N759 = N815 & way_i[2];
  assign N816 = N10 & N11;
  assign N10 = ~way_i[0];
  assign N11 = ~way_i[1];
  assign N758 = N816 & way_i[2];
  assign N757 = N813 & N12;
  assign N12 = ~way_i[2];
  assign N756 = N814 & N13;
  assign N13 = ~way_i[2];
  assign N755 = N815 & N14;
  assign N14 = ~way_i[2];
  assign N754 = N816 & N15;
  assign N15 = ~way_i[2];
  assign { N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97 } = (N16)? { N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33 } :
                                                                                                                                                                                                                                                                                                                                                                                                           (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = pending_w_v;
  assign N17 = N32;
  assign wg_ram_addr = (N18)? way_group_i :
                       (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N18 = N292;
  assign N19 = N291;
  assign wg_ram_w_mask = (N20)? { N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319 } :
                         (N21)? { N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535 } :
                         (N294)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N20 = N780;
  assign N21 = N783;
  assign tag_set = (N22)? way_group_o[191:96] :
                   (N23)? way_group_o[95:0] : 1'b0;
  assign N22 = lce_i[0];
  assign N23 = N752;
  assign { tag_o, coh_state_o } = (N24)? tag_set[95:84] :
                                  (N25)? tag_set[83:72] :
                                  (N26)? tag_set[71:60] :
                                  (N27)? tag_set[59:48] :
                                  (N28)? tag_set[47:36] :
                                  (N29)? tag_set[35:24] :
                                  (N30)? tag_set[23:12] :
                                  (N31)? tag_set[11:0] : 1'b0;
  assign N24 = N761;
  assign N25 = N760;
  assign N26 = N759;
  assign N27 = N758;
  assign N28 = N757;
  assign N29 = N756;
  assign N30 = N755;
  assign N31 = N754;
  assign pending_w_v = w_v_i & N786;
  assign pending_v_o = r_v_i & N764;
  assign N32 = ~pending_w_v;
  assign N161 = ~way_group_i[0];
  assign N162 = ~way_group_i[1];
  assign N163 = N161 & N162;
  assign N164 = N161 & way_group_i[1];
  assign N165 = way_group_i[0] & N162;
  assign N166 = way_group_i[0] & way_group_i[1];
  assign N167 = ~way_group_i[2];
  assign N168 = N163 & N167;
  assign N169 = N163 & way_group_i[2];
  assign N170 = N165 & N167;
  assign N171 = N165 & way_group_i[2];
  assign N172 = N164 & N167;
  assign N173 = N164 & way_group_i[2];
  assign N174 = N166 & N167;
  assign N175 = N166 & way_group_i[2];
  assign N176 = ~way_group_i[3];
  assign N177 = N168 & N176;
  assign N178 = N168 & way_group_i[3];
  assign N179 = N170 & N176;
  assign N180 = N170 & way_group_i[3];
  assign N181 = N172 & N176;
  assign N182 = N172 & way_group_i[3];
  assign N183 = N174 & N176;
  assign N184 = N174 & way_group_i[3];
  assign N185 = N169 & N176;
  assign N186 = N169 & way_group_i[3];
  assign N187 = N171 & N176;
  assign N188 = N171 & way_group_i[3];
  assign N189 = N173 & N176;
  assign N190 = N173 & way_group_i[3];
  assign N191 = N175 & N176;
  assign N192 = N175 & way_group_i[3];
  assign N193 = ~way_group_i[4];
  assign N194 = N177 & N193;
  assign N195 = N177 & way_group_i[4];
  assign N196 = N179 & N193;
  assign N197 = N179 & way_group_i[4];
  assign N198 = N181 & N193;
  assign N199 = N181 & way_group_i[4];
  assign N200 = N183 & N193;
  assign N201 = N183 & way_group_i[4];
  assign N202 = N185 & N193;
  assign N203 = N185 & way_group_i[4];
  assign N204 = N187 & N193;
  assign N205 = N187 & way_group_i[4];
  assign N206 = N189 & N193;
  assign N207 = N189 & way_group_i[4];
  assign N208 = N191 & N193;
  assign N209 = N191 & way_group_i[4];
  assign N210 = N178 & N193;
  assign N211 = N178 & way_group_i[4];
  assign N212 = N180 & N193;
  assign N213 = N180 & way_group_i[4];
  assign N214 = N182 & N193;
  assign N215 = N182 & way_group_i[4];
  assign N216 = N184 & N193;
  assign N217 = N184 & way_group_i[4];
  assign N218 = N186 & N193;
  assign N219 = N186 & way_group_i[4];
  assign N220 = N188 & N193;
  assign N221 = N188 & way_group_i[4];
  assign N222 = N190 & N193;
  assign N223 = N190 & way_group_i[4];
  assign N224 = N192 & N193;
  assign N225 = N192 & way_group_i[4];
  assign N226 = ~way_group_i[5];
  assign N227 = N194 & N226;
  assign N228 = N194 & way_group_i[5];
  assign N229 = N196 & N226;
  assign N230 = N196 & way_group_i[5];
  assign N231 = N198 & N226;
  assign N232 = N198 & way_group_i[5];
  assign N233 = N200 & N226;
  assign N234 = N200 & way_group_i[5];
  assign N235 = N202 & N226;
  assign N236 = N202 & way_group_i[5];
  assign N237 = N204 & N226;
  assign N238 = N204 & way_group_i[5];
  assign N239 = N206 & N226;
  assign N240 = N206 & way_group_i[5];
  assign N241 = N208 & N226;
  assign N242 = N208 & way_group_i[5];
  assign N243 = N210 & N226;
  assign N244 = N210 & way_group_i[5];
  assign N245 = N212 & N226;
  assign N246 = N212 & way_group_i[5];
  assign N247 = N214 & N226;
  assign N248 = N214 & way_group_i[5];
  assign N249 = N216 & N226;
  assign N250 = N216 & way_group_i[5];
  assign N251 = N218 & N226;
  assign N252 = N218 & way_group_i[5];
  assign N253 = N220 & N226;
  assign N254 = N220 & way_group_i[5];
  assign N255 = N222 & N226;
  assign N256 = N222 & way_group_i[5];
  assign N257 = N224 & N226;
  assign N258 = N224 & way_group_i[5];
  assign N259 = N195 & N226;
  assign N260 = N195 & way_group_i[5];
  assign N261 = N197 & N226;
  assign N262 = N197 & way_group_i[5];
  assign N263 = N199 & N226;
  assign N264 = N199 & way_group_i[5];
  assign N265 = N201 & N226;
  assign N266 = N201 & way_group_i[5];
  assign N267 = N203 & N226;
  assign N268 = N203 & way_group_i[5];
  assign N269 = N205 & N226;
  assign N270 = N205 & way_group_i[5];
  assign N271 = N207 & N226;
  assign N272 = N207 & way_group_i[5];
  assign N273 = N209 & N226;
  assign N274 = N209 & way_group_i[5];
  assign N275 = N211 & N226;
  assign N276 = N211 & way_group_i[5];
  assign N277 = N213 & N226;
  assign N278 = N213 & way_group_i[5];
  assign N279 = N215 & N226;
  assign N280 = N215 & way_group_i[5];
  assign N281 = N217 & N226;
  assign N282 = N217 & way_group_i[5];
  assign N283 = N219 & N226;
  assign N284 = N219 & way_group_i[5];
  assign N285 = N221 & N226;
  assign N286 = N221 & way_group_i[5];
  assign N287 = N223 & N226;
  assign N288 = N223 & way_group_i[5];
  assign N289 = N225 & N226;
  assign N290 = N225 & way_group_i[5];
  assign wg_ram_r_v = r_v_i & N817;
  assign N817 = N778 | N775;
  assign wg_ram_w_v = w_v_i & N818;
  assign N818 = N767 | N771;
  assign wg_ram_v = wg_ram_r_v | wg_ram_w_v;
  assign N291 = ~wg_ram_v;
  assign N292 = wg_ram_v;
  assign N293 = N783 | N780;
  assign N294 = ~N293;
  assign N751 = r_v_i & N775;

  always @(posedge clk_i) begin
    if(N160) begin
      { pending_bits_r[63:63] } <= { pending_i };
    end
    if(N159) begin
      { pending_bits_r[62:62] } <= { pending_i };
    end
    if(N158) begin
      { pending_bits_r[61:61] } <= { pending_i };
    end
    if(N157) begin
      { pending_bits_r[60:60] } <= { pending_i };
    end
    if(N156) begin
      { pending_bits_r[59:59] } <= { pending_i };
    end
    if(N155) begin
      { pending_bits_r[58:58] } <= { pending_i };
    end
    if(N154) begin
      { pending_bits_r[57:57] } <= { pending_i };
    end
    if(N153) begin
      { pending_bits_r[56:56] } <= { pending_i };
    end
    if(N152) begin
      { pending_bits_r[55:55] } <= { pending_i };
    end
    if(N151) begin
      { pending_bits_r[54:54] } <= { pending_i };
    end
    if(N150) begin
      { pending_bits_r[53:53] } <= { pending_i };
    end
    if(N149) begin
      { pending_bits_r[52:52] } <= { pending_i };
    end
    if(N148) begin
      { pending_bits_r[51:51] } <= { pending_i };
    end
    if(N147) begin
      { pending_bits_r[50:50] } <= { pending_i };
    end
    if(N146) begin
      { pending_bits_r[49:49] } <= { pending_i };
    end
    if(N145) begin
      { pending_bits_r[48:48] } <= { pending_i };
    end
    if(N144) begin
      { pending_bits_r[47:47] } <= { pending_i };
    end
    if(N143) begin
      { pending_bits_r[46:46] } <= { pending_i };
    end
    if(N142) begin
      { pending_bits_r[45:45] } <= { pending_i };
    end
    if(N141) begin
      { pending_bits_r[44:44] } <= { pending_i };
    end
    if(N140) begin
      { pending_bits_r[43:43] } <= { pending_i };
    end
    if(N139) begin
      { pending_bits_r[42:42] } <= { pending_i };
    end
    if(N138) begin
      { pending_bits_r[41:41] } <= { pending_i };
    end
    if(N137) begin
      { pending_bits_r[40:40] } <= { pending_i };
    end
    if(N136) begin
      { pending_bits_r[39:39] } <= { pending_i };
    end
    if(N135) begin
      { pending_bits_r[38:38] } <= { pending_i };
    end
    if(N134) begin
      { pending_bits_r[37:37] } <= { pending_i };
    end
    if(N133) begin
      { pending_bits_r[36:36] } <= { pending_i };
    end
    if(N132) begin
      { pending_bits_r[35:35] } <= { pending_i };
    end
    if(N131) begin
      { pending_bits_r[34:34] } <= { pending_i };
    end
    if(N130) begin
      { pending_bits_r[33:33] } <= { pending_i };
    end
    if(N129) begin
      { pending_bits_r[32:32] } <= { pending_i };
    end
    if(N128) begin
      { pending_bits_r[31:31] } <= { pending_i };
    end
    if(N127) begin
      { pending_bits_r[30:30] } <= { pending_i };
    end
    if(N126) begin
      { pending_bits_r[29:29] } <= { pending_i };
    end
    if(N125) begin
      { pending_bits_r[28:28] } <= { pending_i };
    end
    if(N124) begin
      { pending_bits_r[27:27] } <= { pending_i };
    end
    if(N123) begin
      { pending_bits_r[26:26] } <= { pending_i };
    end
    if(N122) begin
      { pending_bits_r[25:25] } <= { pending_i };
    end
    if(N121) begin
      { pending_bits_r[24:24] } <= { pending_i };
    end
    if(N120) begin
      { pending_bits_r[23:23] } <= { pending_i };
    end
    if(N119) begin
      { pending_bits_r[22:22] } <= { pending_i };
    end
    if(N118) begin
      { pending_bits_r[21:21] } <= { pending_i };
    end
    if(N117) begin
      { pending_bits_r[20:20] } <= { pending_i };
    end
    if(N116) begin
      { pending_bits_r[19:19] } <= { pending_i };
    end
    if(N115) begin
      { pending_bits_r[18:18] } <= { pending_i };
    end
    if(N114) begin
      { pending_bits_r[17:17] } <= { pending_i };
    end
    if(N113) begin
      { pending_bits_r[16:16] } <= { pending_i };
    end
    if(N112) begin
      { pending_bits_r[15:15] } <= { pending_i };
    end
    if(N111) begin
      { pending_bits_r[14:14] } <= { pending_i };
    end
    if(N110) begin
      { pending_bits_r[13:13] } <= { pending_i };
    end
    if(N109) begin
      { pending_bits_r[12:12] } <= { pending_i };
    end
    if(N108) begin
      { pending_bits_r[11:11] } <= { pending_i };
    end
    if(N107) begin
      { pending_bits_r[10:10] } <= { pending_i };
    end
    if(N106) begin
      { pending_bits_r[9:9] } <= { pending_i };
    end
    if(N105) begin
      { pending_bits_r[8:8] } <= { pending_i };
    end
    if(N104) begin
      { pending_bits_r[7:7] } <= { pending_i };
    end
    if(N103) begin
      { pending_bits_r[6:6] } <= { pending_i };
    end
    if(N102) begin
      { pending_bits_r[5:5] } <= { pending_i };
    end
    if(N101) begin
      { pending_bits_r[4:4] } <= { pending_i };
    end
    if(N100) begin
      { pending_bits_r[3:3] } <= { pending_i };
    end
    if(N99) begin
      { pending_bits_r[2:2] } <= { pending_i };
    end
    if(N98) begin
      { pending_bits_r[1:1] } <= { pending_i };
    end
    if(N97) begin
      { pending_bits_r[0:0] } <= { pending_i };
    end
    if(1'b1) begin
      entry_v_o <= N751;
      way_group_v_o <= wg_ram_r_v;
    end
  end


endmodule



module bsg_decode_num_out_p2
(
  i,
  o
);

  input [0:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o = { 1'b0, 1'b1 } << i[0];

endmodule



module bp_cce_gad_num_way_groups_p64_num_lce_p2_lce_assoc_p8_tag_width_p10_harden_p0
(
  clk_i,
  reset_i,
  way_group_i,
  req_lce_i,
  req_tag_i,
  lru_way_i,
  req_type_flag_i,
  lru_dirty_flag_i,
  gad_v_i,
  req_addr_way_o,
  coh_state_o,
  lru_tag_o,
  transfer_flag_o,
  transfer_lce_o,
  transfer_way_o,
  replacement_flag_o,
  upgrade_flag_o,
  invalidate_flag_o,
  exclusive_flag_o,
  sharers_hits_o,
  sharers_ways_o,
  sharers_coh_states_o
);

  input [191:0] way_group_i;
  input [0:0] req_lce_i;
  input [9:0] req_tag_i;
  input [2:0] lru_way_i;
  output [2:0] req_addr_way_o;
  output [1:0] coh_state_o;
  output [9:0] lru_tag_o;
  output [0:0] transfer_lce_o;
  output [2:0] transfer_way_o;
  output [1:0] sharers_hits_o;
  output [5:0] sharers_ways_o;
  output [3:0] sharers_coh_states_o;
  input clk_i;
  input reset_i;
  input req_type_flag_i;
  input lru_dirty_flag_i;
  input gad_v_i;
  output transfer_flag_o;
  output replacement_flag_o;
  output upgrade_flag_o;
  output invalidate_flag_o;
  output exclusive_flag_o;
  wire [2:0] req_addr_way_o,transfer_way_o;
  wire [1:0] coh_state_o,sharers_hits_o,lce_id_one_hot,lru_coh_state,excl_bits,
  sharers_cached,inv_hits,transfer_lce_one_hot;
  wire [9:0] lru_tag_o;
  wire [0:0] transfer_lce_o,transfer_lce_n;
  wire [5:0] sharers_ways_o;
  wire [3:0] sharers_coh_states_o;
  wire transfer_flag_o,replacement_flag_o,upgrade_flag_o,invalidate_flag_o,
  exclusive_flag_o,N0,N1,N2,N3,N4,exclusive_flag_o,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,
  N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,
  N57,N58,N59,hit,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,
  N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,
  N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,
  N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,
  N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,
  N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,
  N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,
  N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,
  N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,
  N208,N209,N210,N211,transfer_lce_v,N212,N213,N214,N215,N216,N217,N218,N219,N220,
  N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,
  N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,
  N253,N254,N255,N256;
  wire [15:0] tag_set_hits;
  assign transfer_flag_o = exclusive_flag_o;

  bsg_decode_num_out_p2
  lce_id_to_one_hot
  (
    .i(req_lce_i[0]),
    .o(lce_id_one_hot)
  );

  assign N5 = way_group_i[11:2] == req_tag_i;
  assign N6 = way_group_i[23:14] == req_tag_i;
  assign N7 = way_group_i[35:26] == req_tag_i;
  assign N8 = way_group_i[47:38] == req_tag_i;
  assign N9 = way_group_i[59:50] == req_tag_i;
  assign N10 = way_group_i[71:62] == req_tag_i;
  assign N11 = way_group_i[83:74] == req_tag_i;
  assign N12 = way_group_i[95:86] == req_tag_i;
  assign N13 = way_group_i[107:98] == req_tag_i;
  assign N14 = way_group_i[119:110] == req_tag_i;
  assign N15 = way_group_i[131:122] == req_tag_i;
  assign N16 = way_group_i[143:134] == req_tag_i;
  assign N17 = way_group_i[155:146] == req_tag_i;
  assign N18 = way_group_i[167:158] == req_tag_i;
  assign N19 = way_group_i[179:170] == req_tag_i;
  assign N20 = way_group_i[191:182] == req_tag_i;

  bsg_encode_one_hot_width_p8
  hit_vec_to_way_id_gen_0__tag_set_hits_to_way_id
  (
    .i(tag_set_hits[7:0]),
    .addr_o(sharers_ways_o[2:0]),
    .v_o(sharers_hits_o[0])
  );


  bsg_encode_one_hot_width_p8
  hit_vec_to_way_id_gen_1__tag_set_hits_to_way_id
  (
    .i(tag_set_hits[15:8]),
    .addr_o(sharers_ways_o[5:3]),
    .v_o(sharers_hits_o[1])
  );

  assign sharers_coh_states_o[1] = (N28)? way_group_i[1] :
                                   (N30)? way_group_i[13] :
                                   (N32)? way_group_i[25] :
                                   (N34)? way_group_i[37] :
                                   (N29)? way_group_i[49] :
                                   (N31)? way_group_i[61] :
                                   (N33)? way_group_i[73] :
                                   (N35)? way_group_i[85] : 1'b0;
  assign sharers_coh_states_o[0] = (N28)? way_group_i[0] :
                                   (N30)? way_group_i[12] :
                                   (N32)? way_group_i[24] :
                                   (N34)? way_group_i[36] :
                                   (N29)? way_group_i[48] :
                                   (N31)? way_group_i[60] :
                                   (N33)? way_group_i[72] :
                                   (N35)? way_group_i[84] : 1'b0;
  assign sharers_coh_states_o[3] = (N43)? way_group_i[97] :
                                   (N45)? way_group_i[109] :
                                   (N47)? way_group_i[121] :
                                   (N49)? way_group_i[133] :
                                   (N44)? way_group_i[145] :
                                   (N46)? way_group_i[157] :
                                   (N48)? way_group_i[169] :
                                   (N50)? way_group_i[181] : 1'b0;
  assign sharers_coh_states_o[2] = (N43)? way_group_i[96] :
                                   (N45)? way_group_i[108] :
                                   (N47)? way_group_i[120] :
                                   (N49)? way_group_i[132] :
                                   (N44)? way_group_i[144] :
                                   (N46)? way_group_i[156] :
                                   (N48)? way_group_i[168] :
                                   (N50)? way_group_i[180] : 1'b0;
  assign N52 = (N51)? tag_set_hits[7] :
               (N0)? tag_set_hits[15] : 1'b0;
  assign N0 = req_lce_i[0];
  assign N53 = (N51)? tag_set_hits[6] :
               (N0)? tag_set_hits[14] : 1'b0;
  assign N54 = (N51)? tag_set_hits[5] :
               (N0)? tag_set_hits[13] : 1'b0;
  assign N55 = (N51)? tag_set_hits[4] :
               (N0)? tag_set_hits[12] : 1'b0;
  assign N56 = (N51)? tag_set_hits[3] :
               (N0)? tag_set_hits[11] : 1'b0;
  assign N57 = (N51)? tag_set_hits[2] :
               (N0)? tag_set_hits[10] : 1'b0;
  assign N58 = (N51)? tag_set_hits[1] :
               (N0)? tag_set_hits[9] : 1'b0;
  assign N59 = (N51)? tag_set_hits[0] :
               (N0)? tag_set_hits[8] : 1'b0;
  assign N62 = (N61)? sharers_ways_o[2] :
               (N0)? sharers_ways_o[5] : 1'b0;
  assign N63 = (N61)? sharers_ways_o[1] :
               (N0)? sharers_ways_o[4] : 1'b0;
  assign N64 = (N61)? sharers_ways_o[0] :
               (N0)? sharers_ways_o[3] : 1'b0;
  assign N66 = (N65)? way_group_i[85] :
               (N0)? way_group_i[181] : 1'b0;
  assign N67 = (N65)? way_group_i[84] :
               (N0)? way_group_i[180] : 1'b0;
  assign N68 = (N65)? way_group_i[73] :
               (N0)? way_group_i[169] : 1'b0;
  assign N69 = (N65)? way_group_i[72] :
               (N0)? way_group_i[168] : 1'b0;
  assign N70 = (N65)? way_group_i[61] :
               (N0)? way_group_i[157] : 1'b0;
  assign N71 = (N65)? way_group_i[60] :
               (N0)? way_group_i[156] : 1'b0;
  assign N72 = (N65)? way_group_i[49] :
               (N0)? way_group_i[145] : 1'b0;
  assign N73 = (N65)? way_group_i[48] :
               (N0)? way_group_i[144] : 1'b0;
  assign N74 = (N65)? way_group_i[37] :
               (N0)? way_group_i[133] : 1'b0;
  assign N75 = (N65)? way_group_i[36] :
               (N0)? way_group_i[132] : 1'b0;
  assign N76 = (N65)? way_group_i[25] :
               (N0)? way_group_i[121] : 1'b0;
  assign N77 = (N65)? way_group_i[24] :
               (N0)? way_group_i[120] : 1'b0;
  assign N78 = (N65)? way_group_i[13] :
               (N0)? way_group_i[109] : 1'b0;
  assign N79 = (N65)? way_group_i[12] :
               (N0)? way_group_i[108] : 1'b0;
  assign N80 = (N65)? way_group_i[1] :
               (N0)? way_group_i[97] : 1'b0;
  assign N81 = (N65)? way_group_i[0] :
               (N0)? way_group_i[96] : 1'b0;
  assign N97 = (N89)? N80 :
               (N91)? N78 :
               (N93)? N76 :
               (N95)? N74 :
               (N90)? N72 :
               (N92)? N70 :
               (N94)? N68 :
               (N96)? N66 : 1'b0;
  assign N98 = (N89)? N81 :
               (N91)? N79 :
               (N93)? N77 :
               (N95)? N75 :
               (N90)? N73 :
               (N92)? N71 :
               (N94)? N69 :
               (N96)? N67 : 1'b0;
  assign N100 = (N99)? way_group_i[95] :
                (N0)? way_group_i[191] : 1'b0;
  assign N101 = (N99)? way_group_i[94] :
                (N0)? way_group_i[190] : 1'b0;
  assign N102 = (N99)? way_group_i[93] :
                (N0)? way_group_i[189] : 1'b0;
  assign N103 = (N99)? way_group_i[92] :
                (N0)? way_group_i[188] : 1'b0;
  assign N104 = (N99)? way_group_i[91] :
                (N0)? way_group_i[187] : 1'b0;
  assign N105 = (N99)? way_group_i[90] :
                (N0)? way_group_i[186] : 1'b0;
  assign N106 = (N99)? way_group_i[89] :
                (N0)? way_group_i[185] : 1'b0;
  assign N107 = (N99)? way_group_i[88] :
                (N0)? way_group_i[184] : 1'b0;
  assign N108 = (N99)? way_group_i[87] :
                (N0)? way_group_i[183] : 1'b0;
  assign N109 = (N99)? way_group_i[86] :
                (N0)? way_group_i[182] : 1'b0;
  assign N110 = (N99)? way_group_i[83] :
                (N0)? way_group_i[179] : 1'b0;
  assign N111 = (N99)? way_group_i[82] :
                (N0)? way_group_i[178] : 1'b0;
  assign N112 = (N99)? way_group_i[81] :
                (N0)? way_group_i[177] : 1'b0;
  assign N113 = (N99)? way_group_i[80] :
                (N0)? way_group_i[176] : 1'b0;
  assign N114 = (N99)? way_group_i[79] :
                (N0)? way_group_i[175] : 1'b0;
  assign N115 = (N99)? way_group_i[78] :
                (N0)? way_group_i[174] : 1'b0;
  assign N116 = (N99)? way_group_i[77] :
                (N0)? way_group_i[173] : 1'b0;
  assign N117 = (N99)? way_group_i[76] :
                (N0)? way_group_i[172] : 1'b0;
  assign N118 = (N99)? way_group_i[75] :
                (N0)? way_group_i[171] : 1'b0;
  assign N119 = (N99)? way_group_i[74] :
                (N0)? way_group_i[170] : 1'b0;
  assign N120 = (N99)? way_group_i[71] :
                (N0)? way_group_i[167] : 1'b0;
  assign N121 = (N99)? way_group_i[70] :
                (N0)? way_group_i[166] : 1'b0;
  assign N122 = (N99)? way_group_i[69] :
                (N0)? way_group_i[165] : 1'b0;
  assign N123 = (N99)? way_group_i[68] :
                (N0)? way_group_i[164] : 1'b0;
  assign N124 = (N99)? way_group_i[67] :
                (N0)? way_group_i[163] : 1'b0;
  assign N125 = (N99)? way_group_i[66] :
                (N0)? way_group_i[162] : 1'b0;
  assign N126 = (N99)? way_group_i[65] :
                (N0)? way_group_i[161] : 1'b0;
  assign N127 = (N99)? way_group_i[64] :
                (N0)? way_group_i[160] : 1'b0;
  assign N128 = (N99)? way_group_i[63] :
                (N0)? way_group_i[159] : 1'b0;
  assign N129 = (N99)? way_group_i[62] :
                (N0)? way_group_i[158] : 1'b0;
  assign N130 = (N99)? way_group_i[59] :
                (N0)? way_group_i[155] : 1'b0;
  assign N131 = (N99)? way_group_i[58] :
                (N0)? way_group_i[154] : 1'b0;
  assign N132 = (N99)? way_group_i[57] :
                (N0)? way_group_i[153] : 1'b0;
  assign N133 = (N99)? way_group_i[56] :
                (N0)? way_group_i[152] : 1'b0;
  assign N134 = (N99)? way_group_i[55] :
                (N0)? way_group_i[151] : 1'b0;
  assign N135 = (N99)? way_group_i[54] :
                (N0)? way_group_i[150] : 1'b0;
  assign N136 = (N99)? way_group_i[53] :
                (N0)? way_group_i[149] : 1'b0;
  assign N137 = (N99)? way_group_i[52] :
                (N0)? way_group_i[148] : 1'b0;
  assign N138 = (N99)? way_group_i[51] :
                (N0)? way_group_i[147] : 1'b0;
  assign N139 = (N99)? way_group_i[50] :
                (N0)? way_group_i[146] : 1'b0;
  assign N140 = (N99)? way_group_i[47] :
                (N0)? way_group_i[143] : 1'b0;
  assign N141 = (N99)? way_group_i[46] :
                (N0)? way_group_i[142] : 1'b0;
  assign N142 = (N99)? way_group_i[45] :
                (N0)? way_group_i[141] : 1'b0;
  assign N143 = (N99)? way_group_i[44] :
                (N0)? way_group_i[140] : 1'b0;
  assign N144 = (N99)? way_group_i[43] :
                (N0)? way_group_i[139] : 1'b0;
  assign N145 = (N99)? way_group_i[42] :
                (N0)? way_group_i[138] : 1'b0;
  assign N146 = (N99)? way_group_i[41] :
                (N0)? way_group_i[137] : 1'b0;
  assign N147 = (N99)? way_group_i[40] :
                (N0)? way_group_i[136] : 1'b0;
  assign N148 = (N99)? way_group_i[39] :
                (N0)? way_group_i[135] : 1'b0;
  assign N149 = (N99)? way_group_i[38] :
                (N0)? way_group_i[134] : 1'b0;
  assign N150 = (N99)? way_group_i[35] :
                (N0)? way_group_i[131] : 1'b0;
  assign N151 = (N99)? way_group_i[34] :
                (N0)? way_group_i[130] : 1'b0;
  assign N152 = (N99)? way_group_i[33] :
                (N0)? way_group_i[129] : 1'b0;
  assign N153 = (N99)? way_group_i[32] :
                (N0)? way_group_i[128] : 1'b0;
  assign N154 = (N99)? way_group_i[31] :
                (N0)? way_group_i[127] : 1'b0;
  assign N155 = (N99)? way_group_i[30] :
                (N0)? way_group_i[126] : 1'b0;
  assign N156 = (N99)? way_group_i[29] :
                (N0)? way_group_i[125] : 1'b0;
  assign N157 = (N99)? way_group_i[28] :
                (N0)? way_group_i[124] : 1'b0;
  assign N158 = (N99)? way_group_i[27] :
                (N0)? way_group_i[123] : 1'b0;
  assign N159 = (N99)? way_group_i[26] :
                (N0)? way_group_i[122] : 1'b0;
  assign N160 = (N99)? way_group_i[23] :
                (N0)? way_group_i[119] : 1'b0;
  assign N161 = (N99)? way_group_i[22] :
                (N0)? way_group_i[118] : 1'b0;
  assign N162 = (N99)? way_group_i[21] :
                (N0)? way_group_i[117] : 1'b0;
  assign N163 = (N99)? way_group_i[20] :
                (N0)? way_group_i[116] : 1'b0;
  assign N164 = (N99)? way_group_i[19] :
                (N0)? way_group_i[115] : 1'b0;
  assign N165 = (N99)? way_group_i[18] :
                (N0)? way_group_i[114] : 1'b0;
  assign N166 = (N99)? way_group_i[17] :
                (N0)? way_group_i[113] : 1'b0;
  assign N167 = (N99)? way_group_i[16] :
                (N0)? way_group_i[112] : 1'b0;
  assign N168 = (N99)? way_group_i[15] :
                (N0)? way_group_i[111] : 1'b0;
  assign N169 = (N99)? way_group_i[14] :
                (N0)? way_group_i[110] : 1'b0;
  assign N170 = (N99)? way_group_i[11] :
                (N0)? way_group_i[107] : 1'b0;
  assign N171 = (N99)? way_group_i[10] :
                (N0)? way_group_i[106] : 1'b0;
  assign N172 = (N99)? way_group_i[9] :
                (N0)? way_group_i[105] : 1'b0;
  assign N173 = (N99)? way_group_i[8] :
                (N0)? way_group_i[104] : 1'b0;
  assign N174 = (N99)? way_group_i[7] :
                (N0)? way_group_i[103] : 1'b0;
  assign N175 = (N99)? way_group_i[6] :
                (N0)? way_group_i[102] : 1'b0;
  assign N176 = (N99)? way_group_i[5] :
                (N0)? way_group_i[101] : 1'b0;
  assign N177 = (N99)? way_group_i[4] :
                (N0)? way_group_i[100] : 1'b0;
  assign N178 = (N99)? way_group_i[3] :
                (N0)? way_group_i[99] : 1'b0;
  assign N179 = (N99)? way_group_i[2] :
                (N0)? way_group_i[98] : 1'b0;
  assign lru_tag_o[9] = (N187)? N170 :
                        (N189)? N160 :
                        (N191)? N150 :
                        (N193)? N140 :
                        (N188)? N130 :
                        (N190)? N120 :
                        (N192)? N110 :
                        (N194)? N100 : 1'b0;
  assign lru_tag_o[8] = (N187)? N171 :
                        (N189)? N161 :
                        (N191)? N151 :
                        (N193)? N141 :
                        (N188)? N131 :
                        (N190)? N121 :
                        (N192)? N111 :
                        (N194)? N101 : 1'b0;
  assign lru_tag_o[7] = (N187)? N172 :
                        (N189)? N162 :
                        (N191)? N152 :
                        (N193)? N142 :
                        (N188)? N132 :
                        (N190)? N122 :
                        (N192)? N112 :
                        (N194)? N102 : 1'b0;
  assign lru_tag_o[6] = (N187)? N173 :
                        (N189)? N163 :
                        (N191)? N153 :
                        (N193)? N143 :
                        (N188)? N133 :
                        (N190)? N123 :
                        (N192)? N113 :
                        (N194)? N103 : 1'b0;
  assign lru_tag_o[5] = (N187)? N174 :
                        (N189)? N164 :
                        (N191)? N154 :
                        (N193)? N144 :
                        (N188)? N134 :
                        (N190)? N124 :
                        (N192)? N114 :
                        (N194)? N104 : 1'b0;
  assign lru_tag_o[4] = (N187)? N175 :
                        (N189)? N165 :
                        (N191)? N155 :
                        (N193)? N145 :
                        (N188)? N135 :
                        (N190)? N125 :
                        (N192)? N115 :
                        (N194)? N105 : 1'b0;
  assign lru_tag_o[3] = (N187)? N176 :
                        (N189)? N166 :
                        (N191)? N156 :
                        (N193)? N146 :
                        (N188)? N136 :
                        (N190)? N126 :
                        (N192)? N116 :
                        (N194)? N106 : 1'b0;
  assign lru_tag_o[2] = (N187)? N177 :
                        (N189)? N167 :
                        (N191)? N157 :
                        (N193)? N147 :
                        (N188)? N137 :
                        (N190)? N127 :
                        (N192)? N117 :
                        (N194)? N107 : 1'b0;
  assign lru_tag_o[1] = (N187)? N178 :
                        (N189)? N168 :
                        (N191)? N158 :
                        (N193)? N148 :
                        (N188)? N138 :
                        (N190)? N128 :
                        (N192)? N118 :
                        (N194)? N108 : 1'b0;
  assign lru_tag_o[0] = (N187)? N179 :
                        (N189)? N169 :
                        (N191)? N159 :
                        (N193)? N149 :
                        (N188)? N139 :
                        (N190)? N129 :
                        (N192)? N119 :
                        (N194)? N109 : 1'b0;
  assign N196 = (N195)? way_group_i[85] :
                (N0)? way_group_i[181] : 1'b0;
  assign N197 = (N195)? way_group_i[84] :
                (N0)? way_group_i[180] : 1'b0;
  assign N198 = (N195)? way_group_i[73] :
                (N0)? way_group_i[169] : 1'b0;
  assign N199 = (N195)? way_group_i[72] :
                (N0)? way_group_i[168] : 1'b0;
  assign N200 = (N195)? way_group_i[61] :
                (N0)? way_group_i[157] : 1'b0;
  assign N201 = (N195)? way_group_i[60] :
                (N0)? way_group_i[156] : 1'b0;
  assign N202 = (N195)? way_group_i[49] :
                (N0)? way_group_i[145] : 1'b0;
  assign N203 = (N195)? way_group_i[48] :
                (N0)? way_group_i[144] : 1'b0;
  assign N204 = (N195)? way_group_i[37] :
                (N0)? way_group_i[133] : 1'b0;
  assign N205 = (N195)? way_group_i[36] :
                (N0)? way_group_i[132] : 1'b0;
  assign N206 = (N195)? way_group_i[25] :
                (N0)? way_group_i[121] : 1'b0;
  assign N207 = (N195)? way_group_i[24] :
                (N0)? way_group_i[120] : 1'b0;
  assign N208 = (N195)? way_group_i[13] :
                (N0)? way_group_i[109] : 1'b0;
  assign N209 = (N195)? way_group_i[12] :
                (N0)? way_group_i[108] : 1'b0;
  assign N210 = (N195)? way_group_i[1] :
                (N0)? way_group_i[97] : 1'b0;
  assign N211 = (N195)? way_group_i[0] :
                (N0)? way_group_i[96] : 1'b0;
  assign lru_coh_state[1] = (N187)? N210 :
                            (N189)? N208 :
                            (N191)? N206 :
                            (N193)? N204 :
                            (N188)? N202 :
                            (N190)? N200 :
                            (N192)? N198 :
                            (N194)? N196 : 1'b0;
  assign lru_coh_state[0] = (N187)? N211 :
                            (N189)? N209 :
                            (N191)? N207 :
                            (N193)? N205 :
                            (N188)? N203 :
                            (N190)? N201 :
                            (N192)? N199 :
                            (N194)? N197 : 1'b0;

  bsg_encode_one_hot_width_p2
  tag_set_hits_to_way_id
  (
    .i(transfer_lce_one_hot),
    .addr_o(transfer_lce_n[0]),
    .v_o(transfer_lce_v)
  );

  assign N215 = (N214)? sharers_ways_o[2] :
                (N1)? sharers_ways_o[5] : 1'b0;
  assign N1 = transfer_lce_n[0];
  assign N216 = (N214)? sharers_ways_o[1] :
                (N1)? sharers_ways_o[4] : 1'b0;
  assign N217 = (N214)? sharers_ways_o[0] :
                (N1)? sharers_ways_o[3] : 1'b0;
  assign N218 = ~lru_coh_state[1];
  assign N219 = lru_coh_state[0] | N218;
  assign N220 = ~N219;
  assign N221 = lru_coh_state[0] & lru_coh_state[1];
  assign N222 = ~coh_state_o[0];
  assign N223 = N222 | coh_state_o[1];
  assign N224 = ~N223;
  assign req_addr_way_o = (N2)? { N62, N63, N64 } :
                          (N3)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2 = hit;
  assign N3 = N60;
  assign coh_state_o = (N2)? { N97, N98 } :
                       (N3)? { 1'b0, 1'b0 } : 1'b0;
  assign transfer_lce_o[0] = (N4)? transfer_lce_n[0] :
                             (N213)? 1'b0 : 1'b0;
  assign N4 = N212;
  assign transfer_way_o = (N4)? { N215, N216, N217 } :
                          (N213)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_set_hits[0] = N5 & N225;
  assign N225 = way_group_i[1] | way_group_i[0];
  assign tag_set_hits[1] = N6 & N226;
  assign N226 = way_group_i[13] | way_group_i[12];
  assign tag_set_hits[2] = N7 & N227;
  assign N227 = way_group_i[25] | way_group_i[24];
  assign tag_set_hits[3] = N8 & N228;
  assign N228 = way_group_i[37] | way_group_i[36];
  assign tag_set_hits[4] = N9 & N229;
  assign N229 = way_group_i[49] | way_group_i[48];
  assign tag_set_hits[5] = N10 & N230;
  assign N230 = way_group_i[61] | way_group_i[60];
  assign tag_set_hits[6] = N11 & N231;
  assign N231 = way_group_i[73] | way_group_i[72];
  assign tag_set_hits[7] = N12 & N232;
  assign N232 = way_group_i[85] | way_group_i[84];
  assign tag_set_hits[8] = N13 & N233;
  assign N233 = way_group_i[97] | way_group_i[96];
  assign tag_set_hits[9] = N14 & N234;
  assign N234 = way_group_i[109] | way_group_i[108];
  assign tag_set_hits[10] = N15 & N235;
  assign N235 = way_group_i[121] | way_group_i[120];
  assign tag_set_hits[11] = N16 & N236;
  assign N236 = way_group_i[133] | way_group_i[132];
  assign tag_set_hits[12] = N17 & N237;
  assign N237 = way_group_i[145] | way_group_i[144];
  assign tag_set_hits[13] = N18 & N238;
  assign N238 = way_group_i[157] | way_group_i[156];
  assign tag_set_hits[14] = N19 & N239;
  assign N239 = way_group_i[169] | way_group_i[168];
  assign tag_set_hits[15] = N20 & N240;
  assign N240 = way_group_i[181] | way_group_i[180];
  assign N21 = ~sharers_ways_o[0];
  assign N22 = ~sharers_ways_o[1];
  assign N23 = N21 & N22;
  assign N24 = N21 & sharers_ways_o[1];
  assign N25 = sharers_ways_o[0] & N22;
  assign N26 = sharers_ways_o[0] & sharers_ways_o[1];
  assign N27 = ~sharers_ways_o[2];
  assign N28 = N23 & N27;
  assign N29 = N23 & sharers_ways_o[2];
  assign N30 = N25 & N27;
  assign N31 = N25 & sharers_ways_o[2];
  assign N32 = N24 & N27;
  assign N33 = N24 & sharers_ways_o[2];
  assign N34 = N26 & N27;
  assign N35 = N26 & sharers_ways_o[2];
  assign N36 = ~sharers_ways_o[3];
  assign N37 = ~sharers_ways_o[4];
  assign N38 = N36 & N37;
  assign N39 = N36 & sharers_ways_o[4];
  assign N40 = sharers_ways_o[3] & N37;
  assign N41 = sharers_ways_o[3] & sharers_ways_o[4];
  assign N42 = ~sharers_ways_o[5];
  assign N43 = N38 & N42;
  assign N44 = N38 & sharers_ways_o[5];
  assign N45 = N40 & N42;
  assign N46 = N40 & sharers_ways_o[5];
  assign N47 = N39 & N42;
  assign N48 = N39 & sharers_ways_o[5];
  assign N49 = N41 & N42;
  assign N50 = N41 & sharers_ways_o[5];
  assign N51 = ~req_lce_i[0];
  assign hit = N246 | N59;
  assign N246 = N245 | N58;
  assign N245 = N244 | N57;
  assign N244 = N243 | N56;
  assign N243 = N242 | N55;
  assign N242 = N241 | N54;
  assign N241 = N52 | N53;
  assign N60 = ~hit;
  assign N61 = ~req_lce_i[0];
  assign N65 = ~req_lce_i[0];
  assign N82 = ~N64;
  assign N83 = ~N63;
  assign N84 = N82 & N83;
  assign N85 = N82 & N63;
  assign N86 = N64 & N83;
  assign N87 = N64 & N63;
  assign N88 = ~N62;
  assign N89 = N84 & N88;
  assign N90 = N84 & N62;
  assign N91 = N86 & N88;
  assign N92 = N86 & N62;
  assign N93 = N85 & N88;
  assign N94 = N85 & N62;
  assign N95 = N87 & N88;
  assign N96 = N87 & N62;
  assign N99 = ~req_lce_i[0];
  assign N180 = ~lru_way_i[0];
  assign N181 = ~lru_way_i[1];
  assign N182 = N180 & N181;
  assign N183 = N180 & lru_way_i[1];
  assign N184 = lru_way_i[0] & N181;
  assign N185 = lru_way_i[0] & lru_way_i[1];
  assign N186 = ~lru_way_i[2];
  assign N187 = N182 & N186;
  assign N188 = N182 & lru_way_i[2];
  assign N189 = N184 & N186;
  assign N190 = N184 & lru_way_i[2];
  assign N191 = N183 & N186;
  assign N192 = N183 & lru_way_i[2];
  assign N193 = N185 & N186;
  assign N194 = N185 & lru_way_i[2];
  assign N195 = ~req_lce_i[0];
  assign excl_bits[0] = sharers_coh_states_o[1] & sharers_hits_o[0];
  assign excl_bits[1] = sharers_coh_states_o[3] & sharers_hits_o[1];
  assign exclusive_flag_o = N248 | N250;
  assign N248 = excl_bits[1] & N247;
  assign N247 = ~lce_id_one_hot[1];
  assign N250 = excl_bits[0] & N249;
  assign N249 = ~lce_id_one_hot[0];
  assign upgrade_flag_o = N251 & N224;
  assign N251 = hit & req_type_flag_i;
  assign sharers_cached[0] = sharers_coh_states_o[1] | sharers_coh_states_o[0];
  assign sharers_cached[1] = sharers_coh_states_o[3] | sharers_coh_states_o[2];
  assign inv_hits[1] = sharers_hits_o[1] & N247;
  assign inv_hits[0] = sharers_hits_o[0] & N249;
  assign invalidate_flag_o = N255 | exclusive_flag_o;
  assign N255 = req_type_flag_i & N254;
  assign N254 = N252 | N253;
  assign N252 = inv_hits[1] & sharers_cached[1];
  assign N253 = inv_hits[0] & sharers_cached[0];
  assign replacement_flag_o = N256 & lru_dirty_flag_i;
  assign N256 = N220 | N221;
  assign transfer_lce_one_hot[1] = N247 & sharers_hits_o[1];
  assign transfer_lce_one_hot[0] = N249 & sharers_hits_o[0];
  assign N212 = gad_v_i & exclusive_flag_o;
  assign N213 = ~N212;
  assign N214 = ~transfer_lce_n[0];

endmodule



module bp_cce_reg_num_lce_p2_num_cce_p1_addr_width_p22_lce_assoc_p8_lce_sets_p64_block_size_in_bytes_p64_lce_req_data_width_p64
(
  clk_i,
  reset_i,
  decoded_inst_i,
  lce_req_i,
  lce_data_resp_i,
  lce_resp_i,
  mem_resp_i,
  mem_data_resp_i,
  alu_res_i,
  mov_src_i,
  dir_way_group_o_i,
  dir_way_group_v_o_i,
  dir_coh_state_o_i,
  dir_entry_v_o_i,
  dir_pending_o_i,
  dir_pending_v_o_i,
  gad_sharers_hits_i,
  gad_sharers_ways_i,
  gad_sharers_coh_states_i,
  gad_req_addr_way_i,
  gad_coh_state_i,
  gad_lru_tag_i,
  gad_transfer_lce_i,
  gad_transfer_lce_way_i,
  gad_transfer_flag_i,
  gad_replacement_flag_i,
  gad_upgrade_flag_i,
  gad_invalidate_flag_i,
  gad_exclusive_flag_i,
  req_lce_o,
  req_addr_o,
  req_tag_o,
  req_addr_way_o,
  req_coh_state_o,
  lru_way_o,
  lru_addr_o,
  transfer_lce_o,
  transfer_lce_way_o,
  next_coh_state_o,
  cache_block_data_o,
  flags_o,
  gpr_o,
  ack_type_o,
  way_group_o,
  sharers_hits_o,
  sharers_ways_o,
  sharers_coh_states_o,
  nc_req_size_o,
  nc_data_o
);

  input [127:0] decoded_inst_i;
  input [96:0] lce_req_i;
  input [536:0] lce_data_resp_i;
  input [25:0] lce_resp_i;
  input [57:0] mem_resp_i;
  input [541:0] mem_data_resp_i;
  input [15:0] alu_res_i;
  input [15:0] mov_src_i;
  input [191:0] dir_way_group_o_i;
  input [1:0] dir_coh_state_o_i;
  input [1:0] gad_sharers_hits_i;
  input [5:0] gad_sharers_ways_i;
  input [3:0] gad_sharers_coh_states_i;
  input [2:0] gad_req_addr_way_i;
  input [1:0] gad_coh_state_i;
  input [9:0] gad_lru_tag_i;
  input [0:0] gad_transfer_lce_i;
  input [2:0] gad_transfer_lce_way_i;
  output [0:0] req_lce_o;
  output [21:0] req_addr_o;
  output [9:0] req_tag_o;
  output [2:0] req_addr_way_o;
  output [1:0] req_coh_state_o;
  output [2:0] lru_way_o;
  output [21:0] lru_addr_o;
  output [0:0] transfer_lce_o;
  output [2:0] transfer_lce_way_o;
  output [1:0] next_coh_state_o;
  output [511:0] cache_block_data_o;
  output [12:0] flags_o;
  output [63:0] gpr_o;
  output [1:0] ack_type_o;
  output [191:0] way_group_o;
  output [1:0] sharers_hits_o;
  output [5:0] sharers_ways_o;
  output [3:0] sharers_coh_states_o;
  output [1:0] nc_req_size_o;
  output [63:0] nc_data_o;
  input clk_i;
  input reset_i;
  input dir_way_group_v_o_i;
  input dir_entry_v_o_i;
  input dir_pending_o_i;
  input dir_pending_v_o_i;
  input gad_transfer_flag_i;
  input gad_replacement_flag_i;
  input gad_upgrade_flag_i;
  input gad_invalidate_flag_i;
  input gad_exclusive_flag_i;
  wire [9:0] req_tag_o;
  wire [1:0] req_coh_state_o,req_coh_state_n,nc_req_size_n;
  wire [191:0] way_group_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,flags_n_12,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,
  N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,
  N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,
  N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,
  N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,
  N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
  N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,
  N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,
  N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,
  N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,
  N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,
  N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,
  N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
  N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,
  N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,
  N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,
  N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,
  N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,
  N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,
  N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,
  N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,
  N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,
  N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,
  N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,
  N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,
  N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,
  N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,
  N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,
  N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,
  N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,
  N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,
  N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,
  N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,
  N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,
  N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,
  N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,
  N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,
  N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,
  N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,
  N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,
  N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,
  N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,
  N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,
  N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
  N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,
  N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,
  N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,
  N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,
  N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,
  N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,
  N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,
  N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,
  N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,
  N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,
  N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,
  N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,
  N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,
  N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,
  N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,
  N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,
  N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,
  N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,
  N1103,N1104,N1105;
  wire [0:0] req_lce_n,transfer_lce_n;
  wire [21:0] req_addr_n;
  wire [2:0] req_addr_way_n,lru_way_n,transfer_lce_way_n;
  wire [21:6] lru_addr_n;
  wire [511:0] cache_block_data_n;
  wire [10:0] flags_n;
  wire [63:0] gpr_n,nc_data_n;
  reg [1:0] nc_req_size_o,req_coh_state_r,next_coh_state_o,ack_type_o,sharers_hits_o;
  reg [0:0] req_lce_o,transfer_lce_o;
  reg [21:0] req_addr_o,lru_addr_o;
  reg [2:0] req_addr_way_o,lru_way_o,transfer_lce_way_o;
  reg [511:0] cache_block_data_o;
  reg [12:0] flags_o;
  reg [63:0] gpr_o,nc_data_o;
  reg [191:0] way_group_r;
  reg [5:0] sharers_ways_o;
  reg [3:0] sharers_coh_states_o;
  assign req_tag_o[9] = req_addr_o[21];
  assign req_tag_o[8] = req_addr_o[20];
  assign req_tag_o[7] = req_addr_o[19];
  assign req_tag_o[6] = req_addr_o[18];
  assign req_tag_o[5] = req_addr_o[17];
  assign req_tag_o[4] = req_addr_o[16];
  assign req_tag_o[3] = req_addr_o[15];
  assign req_tag_o[2] = req_addr_o[14];
  assign req_tag_o[1] = req_addr_o[13];
  assign req_tag_o[0] = req_addr_o[12];
  assign N64 = N62 & N63;
  assign N65 = decoded_inst_i[92] | N63;
  assign N67 = N62 | decoded_inst_i[91];
  assign N69 = decoded_inst_i[92] & decoded_inst_i[91];
  assign N72 = N70 & N71;
  assign N73 = decoded_inst_i[90] | N71;
  assign N75 = N70 | decoded_inst_i[89];
  assign N77 = decoded_inst_i[90] & decoded_inst_i[89];
  assign N82 = N80 & N81;
  assign N83 = decoded_inst_i[88] | N81;
  assign N85 = N80 | decoded_inst_i[87];
  assign N87 = decoded_inst_i[88] & decoded_inst_i[87];
  assign N94 = N91 & N92;
  assign N95 = N94 & N93;
  assign N96 = decoded_inst_i[84] | decoded_inst_i[83];
  assign N97 = N96 | N93;
  assign N99 = decoded_inst_i[84] | N92;
  assign N100 = N99 | decoded_inst_i[82];
  assign N102 = N99 | N93;
  assign N104 = N91 | decoded_inst_i[83];
  assign N105 = N104 | decoded_inst_i[82];
  assign N107 = decoded_inst_i[84] & decoded_inst_i[82];
  assign N108 = decoded_inst_i[84] & decoded_inst_i[83];
  assign N112 = N110 & N111;
  assign N113 = decoded_inst_i[81] | N111;
  assign N115 = N110 | decoded_inst_i[80];
  assign N117 = decoded_inst_i[81] & decoded_inst_i[80];
  assign N121 = N119 & N120;
  assign N122 = decoded_inst_i[78] | N120;
  assign N124 = N119 | decoded_inst_i[77];
  assign N126 = decoded_inst_i[78] & decoded_inst_i[77];
  assign N1099 = ~decoded_inst_i[114];
  assign N1100 = ~decoded_inst_i[110];
  assign N1101 = decoded_inst_i[113] | N1099;
  assign N1102 = decoded_inst_i[112] | N1101;
  assign N1103 = decoded_inst_i[111] | N1102;
  assign N1104 = N1100 | N1103;
  assign N1105 = ~N1104;
  assign req_coh_state_o = (N0)? dir_coh_state_o_i :
                           (N1)? req_coh_state_r : 1'b0;
  assign N0 = dir_entry_v_o_i;
  assign N1 = N60;
  assign way_group_o = (N2)? dir_way_group_o_i :
                       (N3)? way_group_r : 1'b0;
  assign N2 = dir_way_group_v_o_i;
  assign N3 = N61;
  assign req_lce_n[0] = (N4)? lce_req_i[31] :
                        (N5)? mem_resp_i[34] :
                        (N6)? mem_data_resp_i[518] :
                        (N7)? 1'b0 : 1'b0;
  assign N4 = N64;
  assign N5 = N66;
  assign N6 = N68;
  assign N7 = N69;
  assign req_addr_n = (N4)? lce_req_i[28:7] :
                      (N5)? mem_resp_i[30:9] :
                      (N6)? mem_data_resp_i[540:519] :
                      (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign req_addr_way_n = (N8)? gad_req_addr_way_i :
                          (N9)? mem_resp_i[33:31] :
                          (N10)? mem_data_resp_i[517:515] :
                          (N11)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = N72;
  assign N9 = N74;
  assign N10 = N76;
  assign N11 = N77;
  assign req_coh_state_n = (N12)? gad_coh_state_i :
                           (N211)? dir_coh_state_o_i :
                           (N79)? { 1'b0, 1'b0 } : 1'b0;
  assign N12 = decoded_inst_i[28];
  assign lru_way_n = (N13)? lce_req_i[6:4] :
                     (N14)? mem_resp_i[33:31] :
                     (N15)? mem_data_resp_i[517:515] :
                     (N16)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = N82;
  assign N14 = N84;
  assign N15 = N86;
  assign N16 = N87;
  assign lru_addr_n = (N12)? { gad_lru_tag_i, req_addr_o[11:6] } :
                      (N88)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign transfer_lce_n[0] = (N17)? gad_transfer_lce_i[0] :
                             (N18)? mem_resp_i[8] : 1'b0;
  assign N17 = N89;
  assign N18 = decoded_inst_i[86];
  assign transfer_lce_way_n = (N17)? gad_transfer_lce_way_i :
                              (N18)? mem_resp_i[7:5] : 1'b0;
  assign cache_block_data_n = (N19)? lce_data_resp_i[536:25] :
                              (N20)? mem_data_resp_i[511:0] : 1'b0;
  assign N19 = N90;
  assign N20 = decoded_inst_i[85];
  assign { flags_n_12, flags_n[0:0] } = (N21)? { lce_req_i[2:2], lce_req_i[30:30] } :
                                        (N22)? { mem_resp_i[2:2], mem_resp_i[57:57] } :
                                        (N23)? { mem_data_resp_i[514:514], mem_data_resp_i[541:541] } :
                                        (N24)? { 1'b0, 1'b0 } :
                                        (N25)? { decoded_inst_i[94:94], decoded_inst_i[94:94] } :
                                        (N26)? { 1'b0, 1'b0 } : 1'b0;
  assign N21 = N95;
  assign N22 = N98;
  assign N23 = N101;
  assign N24 = N103;
  assign N25 = N106;
  assign N26 = N109;
  assign nc_req_size_n = (N21)? lce_req_i[1:0] :
                         (N22)? mem_resp_i[1:0] :
                         (N23)? mem_data_resp_i[513:512] :
                         (N24)? { 1'b0, 1'b0 } :
                         (N25)? { 1'b0, 1'b0 } :
                         (N26)? { 1'b0, 1'b0 } : 1'b0;
  assign flags_n[2:1] = (N27)? { lce_req_i[3:3], lce_req_i[29:29] } :
                        (N28)? { 1'b0, 1'b0 } :
                        (N29)? { decoded_inst_i[94:94], decoded_inst_i[94:94] } :
                        (N30)? { 1'b0, 1'b0 } : 1'b0;
  assign N27 = N112;
  assign N28 = N114;
  assign N29 = N116;
  assign N30 = N117;
  assign flags_n[3] = (N31)? lce_data_resp_i[22] :
                      (N32)? decoded_inst_i[94] : 1'b0;
  assign N31 = N118;
  assign N32 = decoded_inst_i[79];
  assign flags_n[4] = (N33)? gad_transfer_flag_i :
                      (N34)? mem_resp_i[4] :
                      (N35)? decoded_inst_i[94] :
                      (N36)? 1'b0 : 1'b0;
  assign N33 = N121;
  assign N34 = N123;
  assign N35 = N125;
  assign N36 = N126;
  assign { flags_n[10:7], flags_n[5:5] } = (N37)? { gad_exclusive_flag_i, gad_invalidate_flag_i, gad_upgrade_flag_i, dir_pending_o_i, gad_replacement_flag_i } :
                                           (N38)? { decoded_inst_i[94:94], decoded_inst_i[94:94], decoded_inst_i[94:94], decoded_inst_i[94:94], decoded_inst_i[94:94] } : 1'b0;
  assign N37 = N127;
  assign N38 = decoded_inst_i[76];
  assign flags_n[6] = (N39)? mem_resp_i[3] :
                      (N40)? decoded_inst_i[94] : 1'b0;
  assign N39 = N128;
  assign N40 = decoded_inst_i[75];
  assign { N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133 } = (N41)? mov_src_i :
                                                                                                              (N42)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N41 = N131;
  assign N42 = N132;
  assign gpr_n[15:0] = (N43)? alu_res_i :
                       (N44)? { N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133 } : 1'b0;
  assign N43 = N129;
  assign N44 = N130;
  assign { N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153 } = (N45)? mov_src_i :
                                                                                                              (N46)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N45 = N151;
  assign N46 = N152;
  assign gpr_n[31:16] = (N47)? alu_res_i :
                        (N48)? { N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153 } : 1'b0;
  assign N47 = N149;
  assign N48 = N150;
  assign { N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173 } = (N49)? mov_src_i :
                                                                                                              (N50)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N49 = N171;
  assign N50 = N172;
  assign gpr_n[47:32] = (N51)? alu_res_i :
                        (N52)? { N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173 } : 1'b0;
  assign N51 = N169;
  assign N52 = N170;
  assign { N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193 } = (N53)? mov_src_i :
                                                                                                              (N54)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N53 = N191;
  assign N54 = N192;
  assign gpr_n[63:48] = (N55)? alu_res_i :
                        (N56)? { N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193 } : 1'b0;
  assign N55 = N189;
  assign N56 = N190;
  assign nc_data_n = (N57)? lce_req_i[96:33] :
                     (N213)? mem_data_resp_i[63:0] :
                     (N210)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N57 = decoded_inst_i[12];
  assign N217 = (N58)? 1'b1 :
                (N59)? decoded_inst_i[34] : 1'b0;
  assign N58 = reset_i;
  assign N59 = N214;
  assign N218 = (N58)? 1'b0 :
                (N59)? req_lce_n[0] : 1'b0;
  assign { N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219 } = (N58)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                  (N59)? req_addr_n : 1'b0;
  assign N241 = (N58)? 1'b1 :
                (N59)? decoded_inst_i[33] : 1'b0;
  assign { N244, N243, N242 } = (N58)? { 1'b0, 1'b0, 1'b0 } :
                                (N59)? req_addr_way_n : 1'b0;
  assign N245 = (N58)? 1'b1 :
                (N59)? N215 : 1'b0;
  assign { N247, N246 } = (N58)? { 1'b0, 1'b0 } :
                          (N59)? req_coh_state_n : 1'b0;
  assign N248 = (N58)? 1'b1 :
                (N59)? decoded_inst_i[32] : 1'b0;
  assign { N251, N250, N249 } = (N58)? { 1'b0, 1'b0, 1'b0 } :
                                (N59)? lru_way_n : 1'b0;
  assign N252 = (N58)? 1'b1 :
                (N59)? decoded_inst_i[28] : 1'b0;
  assign { N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253 } = (N58)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                              (N59)? lru_addr_n : 1'b0;
  assign N269 = (N58)? 1'b1 :
                (N59)? decoded_inst_i[31] : 1'b0;
  assign N270 = (N58)? 1'b0 :
                (N59)? transfer_lce_n[0] : 1'b0;
  assign { N273, N272, N271 } = (N58)? { 1'b0, 1'b0, 1'b0 } :
                                (N59)? transfer_lce_way_n : 1'b0;
  assign N274 = (N58)? 1'b1 :
                (N59)? N216 : 1'b0;
  assign { N276, N275 } = (N58)? { 1'b0, 1'b0 } :
                          (N59)? decoded_inst_i[95:94] : 1'b0;
  assign { N287, N285, N283, N281, N279, N277 } = (N58)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } :
                                                  (N59)? { decoded_inst_i[30:30], decoded_inst_i[30:30], decoded_inst_i[30:30], decoded_inst_i[30:30], decoded_inst_i[30:30], decoded_inst_i[30:30] } : 1'b0;
  assign { N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N286, N284, N282, N280, N278 } = (N58)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N59)? cache_block_data_n : 1'b0;
  assign { N818, N817, N815, N813, N811, N809, N807, N805, N803, N801, N799, N797, N795 } = (N58)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } :
                                                                                            (N59)? decoded_inst_i[25:13] : 1'b0;
  assign { N819, N816, N814, N812, N810, N808, N806, N804, N802, N800, N798, N796 } = (N58)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                      (N59)? { flags_n_12, flags_n } : 1'b0;
  assign { N871, N854, N837, N820 } = (N58)? { 1'b1, 1'b1, 1'b1, 1'b1 } :
                                      (N59)? decoded_inst_i[39:36] : 1'b0;
  assign { N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821 } = (N58)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                                                                                                                                                                                                                                                                              (N59)? gpr_n : 1'b0;
  assign N888 = (N58)? 1'b1 :
                (N59)? decoded_inst_i[29] : 1'b0;
  assign { N890, N889 } = (N58)? { 1'b0, 1'b0 } :
                          (N59)? lce_resp_i[23:22] : 1'b0;
  assign { N893, N891 } = (N58)? { 1'b1, 1'b1 } :
                          (N59)? { dir_way_group_v_o_i, dir_way_group_v_o_i } : 1'b0;
  assign { N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N892 } = (N58)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   (N59)? dir_way_group_o_i : 1'b0;
  assign { N1086, N1085 } = (N58)? { 1'b0, 1'b0 } :
                            (N59)? gad_sharers_hits_i : 1'b0;
  assign { N1092, N1091, N1090, N1089, N1088, N1087 } = (N58)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                        (N59)? gad_sharers_ways_i : 1'b0;
  assign { N1096, N1095, N1094, N1093 } = (N58)? { 1'b0, 1'b0, 1'b0, 1'b0 } :
                                          (N59)? gad_sharers_coh_states_i : 1'b0;
  assign N1097 = (N58)? 1'b0 :
                 (N59)? decoded_inst_i[10] : 1'b0;
  assign N1098 = (N58)? 1'b0 :
                 (N59)? decoded_inst_i[9] : 1'b0;
  assign N60 = ~dir_entry_v_o_i;
  assign N61 = ~dir_way_group_v_o_i;
  assign N62 = ~decoded_inst_i[92];
  assign N63 = ~decoded_inst_i[91];
  assign N66 = ~N65;
  assign N68 = ~N67;
  assign N70 = ~decoded_inst_i[90];
  assign N71 = ~decoded_inst_i[89];
  assign N74 = ~N73;
  assign N76 = ~N75;
  assign N78 = dir_entry_v_o_i | decoded_inst_i[28];
  assign N79 = ~N78;
  assign N80 = ~decoded_inst_i[88];
  assign N81 = ~decoded_inst_i[87];
  assign N84 = ~N83;
  assign N86 = ~N85;
  assign N88 = ~decoded_inst_i[28];
  assign N89 = ~decoded_inst_i[86];
  assign N90 = ~decoded_inst_i[85];
  assign N91 = ~decoded_inst_i[84];
  assign N92 = ~decoded_inst_i[83];
  assign N93 = ~decoded_inst_i[82];
  assign N98 = ~N97;
  assign N101 = ~N100;
  assign N103 = ~N102;
  assign N106 = ~N105;
  assign N109 = N107 | N108;
  assign N110 = ~decoded_inst_i[81];
  assign N111 = ~decoded_inst_i[80];
  assign N114 = ~N113;
  assign N116 = ~N115;
  assign N118 = ~decoded_inst_i[79];
  assign N119 = ~decoded_inst_i[78];
  assign N120 = ~decoded_inst_i[77];
  assign N123 = ~N122;
  assign N125 = ~N124;
  assign N127 = ~decoded_inst_i[76];
  assign N128 = ~decoded_inst_i[75];
  assign N129 = decoded_inst_i[40] & decoded_inst_i[36];
  assign N130 = ~N129;
  assign N131 = decoded_inst_i[41] & decoded_inst_i[36];
  assign N132 = ~N131;
  assign N149 = decoded_inst_i[40] & decoded_inst_i[37];
  assign N150 = ~N149;
  assign N151 = decoded_inst_i[41] & decoded_inst_i[37];
  assign N152 = ~N151;
  assign N169 = decoded_inst_i[40] & decoded_inst_i[38];
  assign N170 = ~N169;
  assign N171 = decoded_inst_i[41] & decoded_inst_i[38];
  assign N172 = ~N171;
  assign N189 = decoded_inst_i[40] & decoded_inst_i[39];
  assign N190 = ~N189;
  assign N191 = decoded_inst_i[41] & decoded_inst_i[39];
  assign N192 = ~N191;
  assign N209 = decoded_inst_i[11] | decoded_inst_i[12];
  assign N210 = ~N209;
  assign N211 = dir_entry_v_o_i & N88;
  assign N212 = ~decoded_inst_i[12];
  assign N213 = decoded_inst_i[11] & N212;
  assign N214 = ~reset_i;
  assign N215 = decoded_inst_i[28] | dir_entry_v_o_i;
  assign N216 = decoded_inst_i[41] & N1105;

  always @(posedge clk_i) begin
    if(N1098) begin
      { nc_req_size_o[1:0] } <= { nc_req_size_n[1:0] };
    end
    if(N217) begin
      { req_lce_o[0:0] } <= { N218 };
      { req_addr_o[21:0] } <= { N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219 };
    end
    if(N241) begin
      { req_addr_way_o[2:0] } <= { N244, N243, N242 };
    end
    if(N245) begin
      { req_coh_state_r[1:0] } <= { N247, N246 };
    end
    if(N248) begin
      { lru_way_o[2:0] } <= { N251, N250, N249 };
    end
    if(N252) begin
      { lru_addr_o[21:0] } <= { N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
      { sharers_hits_o[1:0] } <= { N1086, N1085 };
      { sharers_ways_o[5:0] } <= { N1092, N1091, N1090, N1089, N1088, N1087 };
      { sharers_coh_states_o[3:0] } <= { N1096, N1095, N1094, N1093 };
    end
    if(N269) begin
      { transfer_lce_o[0:0] } <= { N270 };
      { transfer_lce_way_o[2:0] } <= { N273, N272, N271 };
    end
    if(N274) begin
      { next_coh_state_o[1:0] } <= { N276, N275 };
    end
    if(N277) begin
      { cache_block_data_o[511:413], cache_block_data_o[0:0] } <= { N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N278 };
    end
    if(N279) begin
      { cache_block_data_o[412:314], cache_block_data_o[1:1] } <= { N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N280 };
    end
    if(N281) begin
      { cache_block_data_o[313:215], cache_block_data_o[2:2] } <= { N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N282 };
    end
    if(N283) begin
      { cache_block_data_o[214:116], cache_block_data_o[3:3] } <= { N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N284 };
    end
    if(N285) begin
      { cache_block_data_o[115:17], cache_block_data_o[4:4] } <= { N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N286 };
    end
    if(N287) begin
      { cache_block_data_o[16:5] } <= { N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288 };
    end
    if(N818) begin
      { flags_o[12:12] } <= { N819 };
    end
    if(N817) begin
      { flags_o[11:11] } <= { N275 };
    end
    if(N815) begin
      { flags_o[10:10] } <= { N816 };
    end
    if(N813) begin
      { flags_o[9:9] } <= { N814 };
    end
    if(N811) begin
      { flags_o[8:8] } <= { N812 };
    end
    if(N809) begin
      { flags_o[7:7] } <= { N810 };
    end
    if(N807) begin
      { flags_o[6:6] } <= { N808 };
    end
    if(N805) begin
      { flags_o[5:5] } <= { N806 };
    end
    if(N803) begin
      { flags_o[4:4] } <= { N804 };
    end
    if(N801) begin
      { flags_o[3:3] } <= { N802 };
    end
    if(N799) begin
      { flags_o[2:2] } <= { N800 };
    end
    if(N797) begin
      { flags_o[1:1] } <= { N798 };
    end
    if(N795) begin
      { flags_o[0:0] } <= { N796 };
    end
    if(N871) begin
      { gpr_o[63:48] } <= { N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872 };
    end
    if(N854) begin
      { gpr_o[47:32] } <= { N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855 };
    end
    if(N837) begin
      { gpr_o[31:16] } <= { N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838 };
    end
    if(N820) begin
      { gpr_o[15:0] } <= { N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821 };
    end
    if(N888) begin
      { ack_type_o[1:0] } <= { N890, N889 };
    end
    if(N891) begin
      { way_group_r[191:93], way_group_r[0:0] } <= { N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N892 };
    end
    if(N893) begin
      { way_group_r[92:1] } <= { N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894 };
    end
    if(N1097) begin
      { nc_data_o[63:0] } <= { nc_data_n[63:0] };
    end
  end


endmodule



module bp_cce_num_lce_p2_num_cce_p1_paddr_width_p22_lce_assoc_p8_lce_sets_p64_block_size_in_bytes_p64_num_cce_inst_ram_els_p256_lce_req_data_width_p64
(
  clk_i,
  reset_i,
  lce_req_i,
  lce_req_v_i,
  lce_req_yumi_o,
  lce_resp_i,
  lce_resp_v_i,
  lce_resp_yumi_o,
  lce_data_resp_i,
  lce_data_resp_v_i,
  lce_data_resp_yumi_o,
  lce_cmd_o,
  lce_cmd_v_o,
  lce_cmd_ready_i,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i,
  mem_resp_i,
  mem_resp_v_i,
  mem_resp_yumi_o,
  mem_data_resp_i,
  mem_data_resp_v_i,
  mem_data_resp_yumi_o,
  mem_cmd_o,
  mem_cmd_v_o,
  mem_cmd_ready_i,
  mem_data_cmd_o,
  mem_data_cmd_v_o,
  mem_data_cmd_ready_i,
  cce_id_i,
  boot_rom_addr_o,
  boot_rom_data_i
);

  input [96:0] lce_req_i;
  input [25:0] lce_resp_i;
  input [536:0] lce_data_resp_i;
  output [35:0] lce_cmd_o;
  output [517:0] lce_data_cmd_o;
  input [57:0] mem_resp_i;
  input [541:0] mem_data_resp_i;
  output [29:0] mem_cmd_o;
  output [569:0] mem_data_cmd_o;
  input [0:0] cce_id_i;
  output [7:0] boot_rom_addr_o;
  input [95:0] boot_rom_data_i;
  input clk_i;
  input reset_i;
  input lce_req_v_i;
  input lce_resp_v_i;
  input lce_data_resp_v_i;
  input lce_cmd_ready_i;
  input lce_data_cmd_ready_i;
  input mem_resp_v_i;
  input mem_data_resp_v_i;
  input mem_cmd_ready_i;
  input mem_data_cmd_ready_i;
  output lce_req_yumi_o;
  output lce_resp_yumi_o;
  output lce_data_resp_yumi_o;
  output lce_cmd_v_o;
  output lce_data_cmd_v_o;
  output mem_resp_yumi_o;
  output mem_data_resp_yumi_o;
  output mem_cmd_v_o;
  output mem_data_cmd_v_o;
  wire [35:0] lce_cmd_o;
  wire [517:0] lce_data_cmd_o;
  wire [29:0] mem_cmd_o;
  wire [569:0] mem_data_cmd_o;
  wire [7:0] boot_rom_addr_o,decode_branch_target_o;
  wire lce_req_yumi_o,lce_resp_yumi_o,lce_data_resp_yumi_o,lce_cmd_v_o,
  lce_data_cmd_v_o,mem_resp_yumi_o,mem_data_resp_yumi_o,mem_cmd_v_o,mem_data_cmd_v_o,N0,N1,N2,N3,
  N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,
  N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,
  N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,
  N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,
  N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,
  N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,
  alu_branch_res_o,decode_stall_o,pc_inst_v_o,decoded_inst_o_minor_op_u__2_,
  decoded_inst_o_minor_op_u__1_,decoded_inst_o_minor_op_u__0_,decoded_inst_o_src_a__4_,
  decoded_inst_o_src_a__3_,decoded_inst_o_src_a__2_,decoded_inst_o_src_a__1_,
  decoded_inst_o_src_a__0_,decoded_inst_o_src_b__4_,decoded_inst_o_src_b__3_,
  decoded_inst_o_src_b__2_,decoded_inst_o_src_b__1_,decoded_inst_o_src_b__0_,decoded_inst_o_dst__4_,
  decoded_inst_o_dst__3_,decoded_inst_o_dst__2_,decoded_inst_o_dst__1_,
  decoded_inst_o_dst__0_,decoded_inst_o_imm__15_,decoded_inst_o_imm__14_,
  decoded_inst_o_imm__13_,decoded_inst_o_imm__12_,decoded_inst_o_imm__11_,decoded_inst_o_imm__10_,
  decoded_inst_o_imm__9_,decoded_inst_o_imm__8_,decoded_inst_o_imm__7_,
  decoded_inst_o_imm__6_,decoded_inst_o_imm__5_,decoded_inst_o_imm__4_,decoded_inst_o_imm__3_,
  decoded_inst_o_imm__2_,decoded_inst_o_imm__1_,decoded_inst_o_imm__0_,
  decoded_inst_o_alu_v_,decoded_inst_o_req_sel__1_,decoded_inst_o_req_sel__0_,
  decoded_inst_o_req_addr_way_sel__1_,decoded_inst_o_req_addr_way_sel__0_,
  decoded_inst_o_lru_way_sel__1_,decoded_inst_o_lru_way_sel__0_,decoded_inst_o_transfer_lce_sel_,
  decoded_inst_o_cache_block_data_sel_,decoded_inst_o_rqf_sel__2_,decoded_inst_o_rqf_sel__1_,
  decoded_inst_o_rqf_sel__0_,decoded_inst_o_nerldf_sel__1_,
  decoded_inst_o_nerldf_sel__0_,decoded_inst_o_nwbf_sel_,decoded_inst_o_tf_sel__1_,
  decoded_inst_o_tf_sel__0_,decoded_inst_o_pruief_sel_,decoded_inst_o_rwbf_sel_,
  decoded_inst_o_dir_way_group_sel__2_,decoded_inst_o_dir_way_group_sel__1_,
  decoded_inst_o_dir_way_group_sel__0_,decoded_inst_o_dir_lce_sel__2_,decoded_inst_o_dir_lce_sel__1_,
  decoded_inst_o_dir_lce_sel__0_,decoded_inst_o_dir_way_sel__2_,
  decoded_inst_o_dir_way_sel__1_,decoded_inst_o_dir_way_sel__0_,decoded_inst_o_dir_coh_state_sel_,
  decoded_inst_o_dir_tag_sel__1_,decoded_inst_o_dir_tag_sel__0_,decoded_inst_o_dir_r_cmd__2_,
  decoded_inst_o_dir_r_cmd__1_,decoded_inst_o_dir_r_cmd__0_,decoded_inst_o_dir_r_v_,
  decoded_inst_o_dir_w_cmd__2_,decoded_inst_o_dir_w_cmd__1_,
  decoded_inst_o_dir_w_cmd__0_,decoded_inst_o_dir_w_v_,decoded_inst_o_lce_cmd_lce_sel__2_,
  decoded_inst_o_lce_cmd_lce_sel__1_,decoded_inst_o_lce_cmd_lce_sel__0_,
  decoded_inst_o_lce_cmd_addr_sel__2_,decoded_inst_o_lce_cmd_addr_sel__1_,
  decoded_inst_o_lce_cmd_addr_sel__0_,decoded_inst_o_lce_cmd_way_sel__2_,decoded_inst_o_lce_cmd_way_sel__1_,
  decoded_inst_o_lce_cmd_way_sel__0_,decoded_inst_o_mem_data_cmd_addr_sel_,
  decoded_inst_o_mov_dst_w_v_,decoded_inst_o_alu_dst_w_v_,decoded_inst_o_gpr_w_mask__3_,
  decoded_inst_o_gpr_w_mask__2_,decoded_inst_o_gpr_w_mask__1_,
  decoded_inst_o_gpr_w_mask__0_,decoded_inst_o_gpr_w_v_,decoded_inst_o_req_w_v_,
  decoded_inst_o_req_addr_way_w_v_,decoded_inst_o_lru_way_w_v_,decoded_inst_o_transfer_lce_w_v_,
  decoded_inst_o_cache_block_data_w_v_,decoded_inst_o_ack_type_w_v_,decoded_inst_o_gad_op_w_v_,
  decoded_inst_o_rdw_op_w_v_,decoded_inst_o_rde_op_w_v_,
  decoded_inst_o_flag_mask_w_v__12_,decoded_inst_o_flag_mask_w_v__11_,decoded_inst_o_flag_mask_w_v__10_,
  decoded_inst_o_flag_mask_w_v__9_,decoded_inst_o_flag_mask_w_v__8_,
  decoded_inst_o_flag_mask_w_v__7_,decoded_inst_o_flag_mask_w_v__6_,decoded_inst_o_flag_mask_w_v__5_,
  decoded_inst_o_flag_mask_w_v__4_,decoded_inst_o_flag_mask_w_v__3_,
  decoded_inst_o_flag_mask_w_v__2_,decoded_inst_o_flag_mask_w_v__1_,
  decoded_inst_o_flag_mask_w_v__0_,decoded_inst_o_nc_data_lce_req_,decoded_inst_o_nc_data_mem_data_resp_,
  decoded_inst_o_nc_data_w_v_,decoded_inst_o_nc_req_size_w_v_,decoded_inst_v_o,alu_v_o,
  dir_pending_o,dir_pending_v_o,dir_entry_v_o,dir_way_group_v_o,gad_v_i,flags_r_o_3,
  flags_r_o_2,flags_r_o_1,gad_transfer_flag_o,gad_replacement_flag_o,
  gad_upgrade_flag_o,gad_invalidate_flag_o,gad_exclusive_flag_o,N119,N120,N121,N122,N123,N124,
  N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,
  N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,
  N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,
  N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,
  N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,
  N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,
  N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,
  N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,
  N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,
  N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,
  N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,
  N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,
  N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,
  N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
  N349,N350,N351,N352,N353,N354,sharers_hits_r0,N355,N356,N357,N358,N359,N360,N361,
  N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,
  N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,
  N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,
  N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,
  N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,
  N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,
  N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,
  N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,
  N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,
  N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,
  N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,
  N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,
  N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,
  N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,
  N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,
  N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,
  N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,
  N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,
  N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,
  N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,
  N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,
  N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
  N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,
  N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,
  N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,
  N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,
  N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,
  N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,
  N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,
  N826,N827,N828,N829,N830,N831;
  wire [95:0] pc_inst_o;
  wire [15:0] alu_opd_a_i,alu_opd_b_i,alu_res_o,mov_src;
  wire [5:0] dir_way_group_i,gad_sharers_ways_o,sharers_ways_r_o;
  wire [0:0] dir_lce_i,gad_transfer_lce_o;
  wire [2:0] dir_way_i,gad_req_addr_way_o,gad_transfer_lce_way_o,req_addr_way_r_o;
  wire [9:0] dir_tag_i,dir_tag_o,req_tag_r_o,gad_lru_tag_o;
  wire [1:0] dir_coh_state_i,dir_coh_state_o,gad_coh_state_o,gad_sharers_hits_o,
  req_coh_state_r_o,next_coh_state_r_o,ack_type_r_o,sharers_hits_r_o;
  wire [191:0] dir_way_group_o,way_group_r_o;
  wire [11:6] flags_r_o;
  wire [3:0] gad_sharers_coh_states_o,sharers_coh_states_r_o;
  wire [21:0] lru_addr_r_o;
  wire [511:0] cache_block_data_r_o;
  wire [63:0] gpr_r_o,nc_data_r_o;
  assign lce_cmd_o[34] = cce_id_i[0];
  assign mem_data_cmd_o[546] = lce_data_cmd_o[5];
  assign mem_cmd_o[6] = lce_data_cmd_o[5];
  assign mem_data_cmd_o[569] = mem_cmd_o[29];
  assign mem_data_cmd_o[542] = mem_cmd_o[28];
  assign mem_data_cmd_o[541] = mem_cmd_o[27];
  assign mem_data_cmd_o[540] = mem_cmd_o[26];
  assign mem_data_cmd_o[539] = mem_cmd_o[25];
  assign mem_data_cmd_o[538] = mem_cmd_o[24];
  assign mem_data_cmd_o[537] = mem_cmd_o[23];
  assign mem_data_cmd_o[536] = mem_cmd_o[22];
  assign mem_data_cmd_o[535] = mem_cmd_o[21];
  assign mem_data_cmd_o[534] = mem_cmd_o[20];
  assign mem_data_cmd_o[533] = mem_cmd_o[19];
  assign mem_data_cmd_o[532] = mem_cmd_o[18];
  assign mem_data_cmd_o[531] = mem_cmd_o[17];
  assign mem_data_cmd_o[530] = mem_cmd_o[16];
  assign mem_data_cmd_o[529] = mem_cmd_o[15];
  assign mem_data_cmd_o[528] = mem_cmd_o[14];
  assign mem_data_cmd_o[527] = mem_cmd_o[13];
  assign mem_data_cmd_o[526] = mem_cmd_o[12];
  assign mem_data_cmd_o[525] = mem_cmd_o[11];
  assign mem_data_cmd_o[524] = mem_cmd_o[10];
  assign mem_data_cmd_o[523] = mem_cmd_o[9];
  assign mem_data_cmd_o[522] = mem_cmd_o[8];
  assign mem_data_cmd_o[521] = mem_cmd_o[7];
  assign mem_data_cmd_o[545] = mem_cmd_o[5];
  assign mem_data_cmd_o[544] = mem_cmd_o[4];
  assign mem_data_cmd_o[543] = mem_cmd_o[3];
  assign mem_data_cmd_o[514] = mem_cmd_o[2];
  assign mem_data_cmd_o[513] = mem_cmd_o[1];
  assign mem_data_cmd_o[512] = mem_cmd_o[0];

  bp_cce_pc_inst_ram_els_p256_harden_p0
  pc_inst_ram
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .alu_branch_res_i(alu_branch_res_o),
    .pc_stall_i(decode_stall_o),
    .pc_branch_target_i(decode_branch_target_o),
    .inst_o(pc_inst_o),
    .inst_v_o(pc_inst_v_o),
    .boot_rom_addr_o(boot_rom_addr_o),
    .boot_rom_data_i(boot_rom_data_i)
  );


  bp_cce_inst_decode_inst_width_p96_inst_addr_width_p8
  inst_decode
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .inst_i(pc_inst_o),
    .inst_v_i(pc_inst_v_o),
    .lce_req_v_i(lce_req_v_i),
    .lce_resp_v_i(lce_resp_v_i),
    .lce_data_resp_v_i(lce_data_resp_v_i),
    .mem_resp_v_i(mem_resp_v_i),
    .mem_data_resp_v_i(mem_data_resp_v_i),
    .pending_v_i(1'b0),
    .lce_cmd_ready_i(lce_cmd_ready_i),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_i),
    .mem_cmd_ready_i(mem_cmd_ready_i),
    .mem_data_cmd_ready_i(mem_data_cmd_ready_i),
    .decoded_inst_o({ decoded_inst_o_minor_op_u__2_, decoded_inst_o_minor_op_u__1_, decoded_inst_o_minor_op_u__0_, decoded_inst_o_src_a__4_, decoded_inst_o_src_a__3_, decoded_inst_o_src_a__2_, decoded_inst_o_src_a__1_, decoded_inst_o_src_a__0_, decoded_inst_o_src_b__4_, decoded_inst_o_src_b__3_, decoded_inst_o_src_b__2_, decoded_inst_o_src_b__1_, decoded_inst_o_src_b__0_, decoded_inst_o_dst__4_, decoded_inst_o_dst__3_, decoded_inst_o_dst__2_, decoded_inst_o_dst__1_, decoded_inst_o_dst__0_, decoded_inst_o_imm__15_, decoded_inst_o_imm__14_, decoded_inst_o_imm__13_, decoded_inst_o_imm__12_, decoded_inst_o_imm__11_, decoded_inst_o_imm__10_, decoded_inst_o_imm__9_, decoded_inst_o_imm__8_, decoded_inst_o_imm__7_, decoded_inst_o_imm__6_, decoded_inst_o_imm__5_, decoded_inst_o_imm__4_, decoded_inst_o_imm__3_, decoded_inst_o_imm__2_, decoded_inst_o_imm__1_, decoded_inst_o_imm__0_, decoded_inst_o_alu_v_, decoded_inst_o_req_sel__1_, decoded_inst_o_req_sel__0_, decoded_inst_o_req_addr_way_sel__1_, decoded_inst_o_req_addr_way_sel__0_, decoded_inst_o_lru_way_sel__1_, decoded_inst_o_lru_way_sel__0_, decoded_inst_o_transfer_lce_sel_, decoded_inst_o_cache_block_data_sel_, decoded_inst_o_rqf_sel__2_, decoded_inst_o_rqf_sel__1_, decoded_inst_o_rqf_sel__0_, decoded_inst_o_nerldf_sel__1_, decoded_inst_o_nerldf_sel__0_, decoded_inst_o_nwbf_sel_, decoded_inst_o_tf_sel__1_, decoded_inst_o_tf_sel__0_, decoded_inst_o_pruief_sel_, decoded_inst_o_rwbf_sel_, decoded_inst_o_dir_way_group_sel__2_, decoded_inst_o_dir_way_group_sel__1_, decoded_inst_o_dir_way_group_sel__0_, decoded_inst_o_dir_lce_sel__2_, decoded_inst_o_dir_lce_sel__1_, decoded_inst_o_dir_lce_sel__0_, decoded_inst_o_dir_way_sel__2_, decoded_inst_o_dir_way_sel__1_, decoded_inst_o_dir_way_sel__0_, decoded_inst_o_dir_coh_state_sel_, decoded_inst_o_dir_tag_sel__1_, decoded_inst_o_dir_tag_sel__0_, decoded_inst_o_dir_r_cmd__2_, decoded_inst_o_dir_r_cmd__1_, decoded_inst_o_dir_r_cmd__0_, decoded_inst_o_dir_r_v_, decoded_inst_o_dir_w_cmd__2_, decoded_inst_o_dir_w_cmd__1_, decoded_inst_o_dir_w_cmd__0_, decoded_inst_o_dir_w_v_, decoded_inst_o_lce_cmd_lce_sel__2_, decoded_inst_o_lce_cmd_lce_sel__1_, decoded_inst_o_lce_cmd_lce_sel__0_, decoded_inst_o_lce_cmd_addr_sel__2_, decoded_inst_o_lce_cmd_addr_sel__1_, decoded_inst_o_lce_cmd_addr_sel__0_, decoded_inst_o_lce_cmd_way_sel__2_, decoded_inst_o_lce_cmd_way_sel__1_, decoded_inst_o_lce_cmd_way_sel__0_, lce_cmd_o[33:31], decoded_inst_o_mem_data_cmd_addr_sel_, decoded_inst_o_mov_dst_w_v_, decoded_inst_o_alu_dst_w_v_, decoded_inst_o_gpr_w_mask__3_, decoded_inst_o_gpr_w_mask__2_, decoded_inst_o_gpr_w_mask__1_, decoded_inst_o_gpr_w_mask__0_, decoded_inst_o_gpr_w_v_, decoded_inst_o_req_w_v_, decoded_inst_o_req_addr_way_w_v_, decoded_inst_o_lru_way_w_v_, decoded_inst_o_transfer_lce_w_v_, decoded_inst_o_cache_block_data_w_v_, decoded_inst_o_ack_type_w_v_, decoded_inst_o_gad_op_w_v_, decoded_inst_o_rdw_op_w_v_, decoded_inst_o_rde_op_w_v_, decoded_inst_o_flag_mask_w_v__12_, decoded_inst_o_flag_mask_w_v__11_, decoded_inst_o_flag_mask_w_v__10_, decoded_inst_o_flag_mask_w_v__9_, decoded_inst_o_flag_mask_w_v__8_, decoded_inst_o_flag_mask_w_v__7_, decoded_inst_o_flag_mask_w_v__6_, decoded_inst_o_flag_mask_w_v__5_, decoded_inst_o_flag_mask_w_v__4_, decoded_inst_o_flag_mask_w_v__3_, decoded_inst_o_flag_mask_w_v__2_, decoded_inst_o_flag_mask_w_v__1_, decoded_inst_o_flag_mask_w_v__0_, decoded_inst_o_nc_data_lce_req_, decoded_inst_o_nc_data_mem_data_resp_, decoded_inst_o_nc_data_w_v_, decoded_inst_o_nc_req_size_w_v_, lce_req_yumi_o, lce_resp_yumi_o, lce_data_resp_yumi_o, mem_resp_yumi_o, mem_data_resp_yumi_o, lce_cmd_v_o, lce_data_cmd_v_o, mem_cmd_v_o, mem_data_cmd_v_o }),
    .decoded_inst_v_o(decoded_inst_v_o),
    .pc_stall_o(decode_stall_o),
    .pc_branch_target_o(decode_branch_target_o)
  );


  bp_cce_alu_width_p16
  alu
  (
    .v_i(decoded_inst_o_alu_v_),
    .opd_a_i(alu_opd_a_i),
    .opd_b_i(alu_opd_b_i),
    .alu_op_i({ decoded_inst_o_minor_op_u__2_, decoded_inst_o_minor_op_u__1_, decoded_inst_o_minor_op_u__0_ }),
    .v_o(alu_v_o),
    .res_o(alu_res_o),
    .branch_res_o(alu_branch_res_o)
  );


  bp_cce_dir_num_way_groups_p64_num_lce_p2_lce_assoc_p8_tag_width_p10_harden_p0
  directory
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .way_group_i(dir_way_group_i),
    .lce_i(dir_lce_i[0]),
    .way_i(dir_way_i),
    .r_cmd_i({ decoded_inst_o_dir_r_cmd__2_, decoded_inst_o_dir_r_cmd__1_, decoded_inst_o_dir_r_cmd__0_ }),
    .r_v_i(decoded_inst_o_dir_r_v_),
    .tag_i(dir_tag_i),
    .coh_state_i(dir_coh_state_i),
    .pending_i(decoded_inst_o_imm__0_),
    .w_cmd_i({ decoded_inst_o_dir_w_cmd__2_, decoded_inst_o_dir_w_cmd__1_, decoded_inst_o_dir_w_cmd__0_ }),
    .w_v_i(decoded_inst_o_dir_w_v_),
    .pending_o(dir_pending_o),
    .pending_v_o(dir_pending_v_o),
    .tag_o(dir_tag_o),
    .coh_state_o(dir_coh_state_o),
    .entry_v_o(dir_entry_v_o),
    .way_group_o(dir_way_group_o),
    .way_group_v_o(dir_way_group_v_o)
  );


  bp_cce_gad_num_way_groups_p64_num_lce_p2_lce_assoc_p8_tag_width_p10_harden_p0
  gad
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .way_group_i(way_group_r_o),
    .req_lce_i(lce_data_cmd_o[5]),
    .req_tag_i(req_tag_r_o),
    .lru_way_i(mem_cmd_o[5:3]),
    .req_type_flag_i(mem_cmd_o[29]),
    .lru_dirty_flag_i(flags_r_o_2),
    .gad_v_i(gad_v_i),
    .req_addr_way_o(gad_req_addr_way_o),
    .coh_state_o(gad_coh_state_o),
    .lru_tag_o(gad_lru_tag_o),
    .transfer_flag_o(gad_transfer_flag_o),
    .transfer_lce_o(gad_transfer_lce_o[0]),
    .transfer_way_o(gad_transfer_lce_way_o),
    .replacement_flag_o(gad_replacement_flag_o),
    .upgrade_flag_o(gad_upgrade_flag_o),
    .invalidate_flag_o(gad_invalidate_flag_o),
    .exclusive_flag_o(gad_exclusive_flag_o),
    .sharers_hits_o(gad_sharers_hits_o),
    .sharers_ways_o(gad_sharers_ways_o),
    .sharers_coh_states_o(gad_sharers_coh_states_o)
  );


  bp_cce_reg_num_lce_p2_num_cce_p1_addr_width_p22_lce_assoc_p8_lce_sets_p64_block_size_in_bytes_p64_lce_req_data_width_p64
  cce_reg
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .decoded_inst_i({ decoded_inst_o_minor_op_u__2_, decoded_inst_o_minor_op_u__1_, decoded_inst_o_minor_op_u__0_, decoded_inst_o_src_a__4_, decoded_inst_o_src_a__3_, decoded_inst_o_src_a__2_, decoded_inst_o_src_a__1_, decoded_inst_o_src_a__0_, decoded_inst_o_src_b__4_, decoded_inst_o_src_b__3_, decoded_inst_o_src_b__2_, decoded_inst_o_src_b__1_, decoded_inst_o_src_b__0_, decoded_inst_o_dst__4_, decoded_inst_o_dst__3_, decoded_inst_o_dst__2_, decoded_inst_o_dst__1_, decoded_inst_o_dst__0_, decoded_inst_o_imm__15_, decoded_inst_o_imm__14_, decoded_inst_o_imm__13_, decoded_inst_o_imm__12_, decoded_inst_o_imm__11_, decoded_inst_o_imm__10_, decoded_inst_o_imm__9_, decoded_inst_o_imm__8_, decoded_inst_o_imm__7_, decoded_inst_o_imm__6_, decoded_inst_o_imm__5_, decoded_inst_o_imm__4_, decoded_inst_o_imm__3_, decoded_inst_o_imm__2_, decoded_inst_o_imm__1_, decoded_inst_o_imm__0_, decoded_inst_o_alu_v_, decoded_inst_o_req_sel__1_, decoded_inst_o_req_sel__0_, decoded_inst_o_req_addr_way_sel__1_, decoded_inst_o_req_addr_way_sel__0_, decoded_inst_o_lru_way_sel__1_, decoded_inst_o_lru_way_sel__0_, decoded_inst_o_transfer_lce_sel_, decoded_inst_o_cache_block_data_sel_, decoded_inst_o_rqf_sel__2_, decoded_inst_o_rqf_sel__1_, decoded_inst_o_rqf_sel__0_, decoded_inst_o_nerldf_sel__1_, decoded_inst_o_nerldf_sel__0_, decoded_inst_o_nwbf_sel_, decoded_inst_o_tf_sel__1_, decoded_inst_o_tf_sel__0_, decoded_inst_o_pruief_sel_, decoded_inst_o_rwbf_sel_, decoded_inst_o_dir_way_group_sel__2_, decoded_inst_o_dir_way_group_sel__1_, decoded_inst_o_dir_way_group_sel__0_, decoded_inst_o_dir_lce_sel__2_, decoded_inst_o_dir_lce_sel__1_, decoded_inst_o_dir_lce_sel__0_, decoded_inst_o_dir_way_sel__2_, decoded_inst_o_dir_way_sel__1_, decoded_inst_o_dir_way_sel__0_, decoded_inst_o_dir_coh_state_sel_, decoded_inst_o_dir_tag_sel__1_, decoded_inst_o_dir_tag_sel__0_, decoded_inst_o_dir_r_cmd__2_, decoded_inst_o_dir_r_cmd__1_, decoded_inst_o_dir_r_cmd__0_, decoded_inst_o_dir_r_v_, decoded_inst_o_dir_w_cmd__2_, decoded_inst_o_dir_w_cmd__1_, decoded_inst_o_dir_w_cmd__0_, decoded_inst_o_dir_w_v_, decoded_inst_o_lce_cmd_lce_sel__2_, decoded_inst_o_lce_cmd_lce_sel__1_, decoded_inst_o_lce_cmd_lce_sel__0_, decoded_inst_o_lce_cmd_addr_sel__2_, decoded_inst_o_lce_cmd_addr_sel__1_, decoded_inst_o_lce_cmd_addr_sel__0_, decoded_inst_o_lce_cmd_way_sel__2_, decoded_inst_o_lce_cmd_way_sel__1_, decoded_inst_o_lce_cmd_way_sel__0_, lce_cmd_o[33:31], decoded_inst_o_mem_data_cmd_addr_sel_, decoded_inst_o_mov_dst_w_v_, decoded_inst_o_alu_dst_w_v_, decoded_inst_o_gpr_w_mask__3_, decoded_inst_o_gpr_w_mask__2_, decoded_inst_o_gpr_w_mask__1_, decoded_inst_o_gpr_w_mask__0_, decoded_inst_o_gpr_w_v_, decoded_inst_o_req_w_v_, decoded_inst_o_req_addr_way_w_v_, decoded_inst_o_lru_way_w_v_, decoded_inst_o_transfer_lce_w_v_, decoded_inst_o_cache_block_data_w_v_, decoded_inst_o_ack_type_w_v_, decoded_inst_o_gad_op_w_v_, decoded_inst_o_rdw_op_w_v_, decoded_inst_o_rde_op_w_v_, decoded_inst_o_flag_mask_w_v__12_, decoded_inst_o_flag_mask_w_v__11_, decoded_inst_o_flag_mask_w_v__10_, decoded_inst_o_flag_mask_w_v__9_, decoded_inst_o_flag_mask_w_v__8_, decoded_inst_o_flag_mask_w_v__7_, decoded_inst_o_flag_mask_w_v__6_, decoded_inst_o_flag_mask_w_v__5_, decoded_inst_o_flag_mask_w_v__4_, decoded_inst_o_flag_mask_w_v__3_, decoded_inst_o_flag_mask_w_v__2_, decoded_inst_o_flag_mask_w_v__1_, decoded_inst_o_flag_mask_w_v__0_, decoded_inst_o_nc_data_lce_req_, decoded_inst_o_nc_data_mem_data_resp_, decoded_inst_o_nc_data_w_v_, decoded_inst_o_nc_req_size_w_v_, lce_req_yumi_o, lce_resp_yumi_o, lce_data_resp_yumi_o, mem_resp_yumi_o, mem_data_resp_yumi_o, lce_cmd_v_o, lce_data_cmd_v_o, mem_cmd_v_o, mem_data_cmd_v_o }),
    .lce_req_i(lce_req_i),
    .lce_data_resp_i(lce_data_resp_i),
    .lce_resp_i(lce_resp_i),
    .mem_resp_i(mem_resp_i),
    .mem_data_resp_i(mem_data_resp_i),
    .alu_res_i(alu_res_o),
    .mov_src_i(mov_src),
    .dir_way_group_o_i(dir_way_group_o),
    .dir_way_group_v_o_i(dir_way_group_v_o),
    .dir_coh_state_o_i(dir_coh_state_o),
    .dir_entry_v_o_i(dir_entry_v_o),
    .dir_pending_o_i(dir_pending_o),
    .dir_pending_v_o_i(dir_pending_v_o),
    .gad_sharers_hits_i(gad_sharers_hits_o),
    .gad_sharers_ways_i(gad_sharers_ways_o),
    .gad_sharers_coh_states_i(gad_sharers_coh_states_o),
    .gad_req_addr_way_i(gad_req_addr_way_o),
    .gad_coh_state_i(gad_coh_state_o),
    .gad_lru_tag_i(gad_lru_tag_o),
    .gad_transfer_lce_i(gad_transfer_lce_o[0]),
    .gad_transfer_lce_way_i(gad_transfer_lce_way_o),
    .gad_transfer_flag_i(gad_transfer_flag_o),
    .gad_replacement_flag_i(gad_replacement_flag_o),
    .gad_upgrade_flag_i(gad_upgrade_flag_o),
    .gad_invalidate_flag_i(gad_invalidate_flag_o),
    .gad_exclusive_flag_i(gad_exclusive_flag_o),
    .req_lce_o(lce_data_cmd_o[5]),
    .req_addr_o(mem_cmd_o[28:7]),
    .req_tag_o(req_tag_r_o),
    .req_addr_way_o(req_addr_way_r_o),
    .req_coh_state_o(req_coh_state_r_o),
    .lru_way_o(mem_cmd_o[5:3]),
    .lru_addr_o(lru_addr_r_o),
    .transfer_lce_o(mem_data_cmd_o[520]),
    .transfer_lce_way_o(mem_data_cmd_o[519:517]),
    .next_coh_state_o(next_coh_state_r_o),
    .cache_block_data_o(cache_block_data_r_o),
    .flags_o({ mem_cmd_o[2:2], flags_r_o, mem_data_cmd_o[515:515], mem_data_cmd_o[516:516], flags_r_o_3, flags_r_o_2, flags_r_o_1, mem_cmd_o[29:29] }),
    .gpr_o(gpr_r_o),
    .ack_type_o(ack_type_r_o),
    .way_group_o(way_group_r_o),
    .sharers_hits_o(sharers_hits_r_o),
    .sharers_ways_o(sharers_ways_r_o),
    .sharers_coh_states_o(sharers_coh_states_r_o),
    .nc_req_size_o(mem_cmd_o[1:0]),
    .nc_data_o(nc_data_r_o)
  );

  assign N122 = N119 & N120;
  assign N123 = N122 & N121;
  assign N125 = decoded_inst_o_lce_cmd_lce_sel__2_ | decoded_inst_o_lce_cmd_lce_sel__1_;
  assign N126 = N125 | N124;
  assign N129 = decoded_inst_o_lce_cmd_lce_sel__2_ | N128;
  assign N130 = N129 | decoded_inst_o_lce_cmd_lce_sel__0_;
  assign N134 = decoded_inst_o_lce_cmd_lce_sel__2_ | N132;
  assign N135 = N134 | N133;
  assign N138 = N137 | decoded_inst_o_lce_cmd_lce_sel__1_;
  assign N139 = N138 | decoded_inst_o_lce_cmd_lce_sel__0_;
  assign N143 = N141 | decoded_inst_o_lce_cmd_lce_sel__1_;
  assign N144 = N143 | N142;
  assign N148 = N146 | N147;
  assign N149 = N148 | decoded_inst_o_lce_cmd_lce_sel__0_;
  assign N151 = decoded_inst_o_lce_cmd_lce_sel__2_ & decoded_inst_o_lce_cmd_lce_sel__1_;
  assign N152 = N151 & decoded_inst_o_lce_cmd_lce_sel__0_;
  assign N156 = N153 & N154;
  assign N157 = N156 & N155;
  assign N159 = decoded_inst_o_lce_cmd_addr_sel__2_ | decoded_inst_o_lce_cmd_addr_sel__1_;
  assign N160 = N159 | N158;
  assign N163 = decoded_inst_o_lce_cmd_addr_sel__2_ | N162;
  assign N164 = N163 | decoded_inst_o_lce_cmd_addr_sel__0_;
  assign N168 = decoded_inst_o_lce_cmd_addr_sel__2_ | N166;
  assign N169 = N168 | N167;
  assign N172 = N171 | decoded_inst_o_lce_cmd_addr_sel__1_;
  assign N173 = N172 | decoded_inst_o_lce_cmd_addr_sel__0_;
  assign N177 = N175 | decoded_inst_o_lce_cmd_addr_sel__1_;
  assign N178 = N177 | N176;
  assign N182 = N180 | N181;
  assign N183 = N182 | decoded_inst_o_lce_cmd_addr_sel__0_;
  assign N185 = decoded_inst_o_lce_cmd_addr_sel__2_ & decoded_inst_o_lce_cmd_addr_sel__1_;
  assign N186 = N185 & decoded_inst_o_lce_cmd_addr_sel__0_;
  assign N218 = N215 & N216;
  assign N219 = N218 & N217;
  assign N221 = decoded_inst_o_lce_cmd_way_sel__2_ | decoded_inst_o_lce_cmd_way_sel__1_;
  assign N222 = N221 | N220;
  assign N225 = decoded_inst_o_lce_cmd_way_sel__2_ | N224;
  assign N226 = N225 | decoded_inst_o_lce_cmd_way_sel__0_;
  assign N230 = decoded_inst_o_lce_cmd_way_sel__2_ | N228;
  assign N231 = N230 | N229;
  assign N234 = N233 | decoded_inst_o_lce_cmd_way_sel__1_;
  assign N235 = N234 | decoded_inst_o_lce_cmd_way_sel__0_;
  assign N237 = decoded_inst_o_lce_cmd_way_sel__2_ & decoded_inst_o_lce_cmd_way_sel__0_;
  assign N238 = decoded_inst_o_lce_cmd_way_sel__2_ & decoded_inst_o_lce_cmd_way_sel__1_;
  assign N241 = (N240)? sharers_ways_r_o[2] :
                (N0)? sharers_ways_r_o[5] : 1'b0;
  assign N0 = gpr_r_o[0];
  assign N242 = (N240)? sharers_ways_r_o[1] :
                (N0)? sharers_ways_r_o[4] : 1'b0;
  assign N243 = (N240)? sharers_ways_r_o[0] :
                (N0)? sharers_ways_r_o[3] : 1'b0;
  assign N253 = N250 & N251;
  assign N254 = N253 & N252;
  assign N256 = decoded_inst_o_dir_way_group_sel__2_ | decoded_inst_o_dir_way_group_sel__1_;
  assign N257 = N256 | N255;
  assign N260 = decoded_inst_o_dir_way_group_sel__2_ | N259;
  assign N261 = N260 | decoded_inst_o_dir_way_group_sel__0_;
  assign N265 = decoded_inst_o_dir_way_group_sel__2_ | N263;
  assign N266 = N265 | N264;
  assign N269 = N268 | decoded_inst_o_dir_way_group_sel__1_;
  assign N270 = N269 | decoded_inst_o_dir_way_group_sel__0_;
  assign N274 = N272 | decoded_inst_o_dir_way_group_sel__1_;
  assign N275 = N274 | N273;
  assign N277 = decoded_inst_o_dir_way_group_sel__2_ & decoded_inst_o_dir_way_group_sel__1_;
  assign N281 = N278 & N279;
  assign N282 = N281 & N280;
  assign N284 = decoded_inst_o_dir_lce_sel__2_ | decoded_inst_o_dir_lce_sel__1_;
  assign N285 = N284 | N283;
  assign N288 = decoded_inst_o_dir_lce_sel__2_ | N287;
  assign N289 = N288 | decoded_inst_o_dir_lce_sel__0_;
  assign N293 = decoded_inst_o_dir_lce_sel__2_ | N291;
  assign N294 = N293 | N292;
  assign N297 = N296 | decoded_inst_o_dir_lce_sel__1_;
  assign N298 = N297 | decoded_inst_o_dir_lce_sel__0_;
  assign N302 = N300 | decoded_inst_o_dir_lce_sel__1_;
  assign N303 = N302 | N301;
  assign N305 = decoded_inst_o_dir_lce_sel__2_ & decoded_inst_o_dir_lce_sel__1_;
  assign N309 = N306 & N307;
  assign N310 = N309 & N308;
  assign N312 = decoded_inst_o_dir_way_sel__2_ | decoded_inst_o_dir_way_sel__1_;
  assign N313 = N312 | N311;
  assign N316 = decoded_inst_o_dir_way_sel__2_ | N315;
  assign N317 = N316 | decoded_inst_o_dir_way_sel__0_;
  assign N321 = decoded_inst_o_dir_way_sel__2_ | N319;
  assign N322 = N321 | N320;
  assign N325 = N324 | decoded_inst_o_dir_way_sel__1_;
  assign N326 = N325 | decoded_inst_o_dir_way_sel__0_;
  assign N330 = N328 | decoded_inst_o_dir_way_sel__1_;
  assign N331 = N330 | N329;
  assign N335 = N333 | N334;
  assign N336 = N335 | decoded_inst_o_dir_way_sel__0_;
  assign N338 = decoded_inst_o_dir_way_sel__2_ & decoded_inst_o_dir_way_sel__1_;
  assign N339 = N338 & decoded_inst_o_dir_way_sel__0_;
  assign N340 = (N240)? sharers_ways_r_o[2] :
                (N0)? sharers_ways_r_o[5] : 1'b0;
  assign N341 = (N240)? sharers_ways_r_o[1] :
                (N0)? sharers_ways_r_o[4] : 1'b0;
  assign N342 = (N240)? sharers_ways_r_o[0] :
                (N0)? sharers_ways_r_o[3] : 1'b0;
  assign N347 = N345 & N346;
  assign N349 = decoded_inst_o_dir_tag_sel__1_ | N348;
  assign N352 = N351 | decoded_inst_o_dir_tag_sel__0_;
  assign N354 = decoded_inst_o_dir_tag_sel__1_ & decoded_inst_o_dir_tag_sel__0_;
  assign sharers_hits_r0 = (N240)? sharers_hits_r_o[0] :
                           (N0)? sharers_hits_r_o[1] : 1'b0;
  assign N360 = N355 & N356;
  assign N361 = N357 & N358;
  assign N362 = N360 & N361;
  assign N363 = N362 & N359;
  assign N365 = decoded_inst_o_src_a__4_ | decoded_inst_o_src_a__3_;
  assign N366 = decoded_inst_o_src_a__2_ | decoded_inst_o_src_a__1_;
  assign N367 = N365 | N366;
  assign N368 = N367 | N364;
  assign N371 = decoded_inst_o_src_a__4_ | decoded_inst_o_src_a__3_;
  assign N372 = decoded_inst_o_src_a__2_ | N370;
  assign N373 = N371 | N372;
  assign N374 = N373 | decoded_inst_o_src_a__0_;
  assign N378 = decoded_inst_o_src_a__4_ | decoded_inst_o_src_a__3_;
  assign N379 = decoded_inst_o_src_a__2_ | N376;
  assign N380 = N378 | N379;
  assign N381 = N380 | N377;
  assign N384 = decoded_inst_o_src_a__4_ | decoded_inst_o_src_a__3_;
  assign N385 = N383 | decoded_inst_o_src_a__1_;
  assign N386 = N384 | N385;
  assign N387 = N386 | decoded_inst_o_src_a__0_;
  assign N391 = decoded_inst_o_src_a__4_ | decoded_inst_o_src_a__3_;
  assign N392 = N389 | decoded_inst_o_src_a__1_;
  assign N393 = N391 | N392;
  assign N394 = N393 | N390;
  assign N398 = decoded_inst_o_src_a__4_ | decoded_inst_o_src_a__3_;
  assign N399 = N396 | N397;
  assign N400 = N398 | N399;
  assign N401 = N400 | decoded_inst_o_src_a__0_;
  assign N406 = decoded_inst_o_src_a__4_ | decoded_inst_o_src_a__3_;
  assign N407 = N403 | N404;
  assign N408 = N406 | N407;
  assign N409 = N408 | N405;
  assign N412 = decoded_inst_o_src_a__4_ | N411;
  assign N413 = decoded_inst_o_src_a__2_ | decoded_inst_o_src_a__1_;
  assign N414 = N412 | N413;
  assign N415 = N414 | decoded_inst_o_src_a__0_;
  assign N419 = decoded_inst_o_src_a__4_ | N417;
  assign N420 = decoded_inst_o_src_a__2_ | decoded_inst_o_src_a__1_;
  assign N421 = N419 | N420;
  assign N422 = N421 | N418;
  assign N426 = decoded_inst_o_src_a__4_ | N424;
  assign N427 = decoded_inst_o_src_a__2_ | N425;
  assign N428 = N426 | N427;
  assign N429 = N428 | decoded_inst_o_src_a__0_;
  assign N434 = decoded_inst_o_src_a__4_ | N431;
  assign N435 = decoded_inst_o_src_a__2_ | N432;
  assign N436 = N434 | N435;
  assign N437 = N436 | N433;
  assign N441 = decoded_inst_o_src_a__4_ | N439;
  assign N442 = N440 | decoded_inst_o_src_a__1_;
  assign N443 = N441 | N442;
  assign N444 = N443 | decoded_inst_o_src_a__0_;
  assign N449 = decoded_inst_o_src_a__4_ | N446;
  assign N450 = N447 | decoded_inst_o_src_a__1_;
  assign N451 = N449 | N450;
  assign N452 = N451 | N448;
  assign N457 = decoded_inst_o_src_a__4_ | N454;
  assign N458 = N455 | N456;
  assign N459 = N457 | N458;
  assign N460 = N459 | decoded_inst_o_src_a__0_;
  assign N466 = decoded_inst_o_src_a__4_ | N462;
  assign N467 = N463 | N464;
  assign N468 = N466 | N467;
  assign N469 = N468 | N465;
  assign N472 = N471 | decoded_inst_o_src_a__3_;
  assign N473 = decoded_inst_o_src_a__2_ | decoded_inst_o_src_a__1_;
  assign N474 = N472 | N473;
  assign N475 = N474 | decoded_inst_o_src_a__0_;
  assign N479 = N477 | decoded_inst_o_src_a__3_;
  assign N480 = decoded_inst_o_src_a__2_ | decoded_inst_o_src_a__1_;
  assign N481 = N479 | N480;
  assign N482 = N481 | N478;
  assign N486 = N484 | decoded_inst_o_src_a__3_;
  assign N487 = decoded_inst_o_src_a__2_ | N485;
  assign N488 = N486 | N487;
  assign N489 = N488 | decoded_inst_o_src_a__0_;
  assign N494 = N491 | decoded_inst_o_src_a__3_;
  assign N495 = decoded_inst_o_src_a__2_ | N492;
  assign N496 = N494 | N495;
  assign N497 = N496 | N493;
  assign N501 = N499 | decoded_inst_o_src_a__3_;
  assign N502 = N500 | decoded_inst_o_src_a__1_;
  assign N503 = N501 | N502;
  assign N504 = N503 | decoded_inst_o_src_a__0_;
  assign N509 = N506 | decoded_inst_o_src_a__3_;
  assign N510 = N507 | decoded_inst_o_src_a__1_;
  assign N511 = N509 | N510;
  assign N512 = N511 | N508;
  assign N517 = N514 | decoded_inst_o_src_a__3_;
  assign N518 = N515 | N516;
  assign N519 = N517 | N518;
  assign N520 = N519 | decoded_inst_o_src_a__0_;
  assign N524 = N522 | N523;
  assign N525 = decoded_inst_o_src_a__2_ | decoded_inst_o_src_a__1_;
  assign N526 = N524 | N525;
  assign N527 = N526 | decoded_inst_o_src_a__0_;
  assign N532 = N529 | N530;
  assign N533 = decoded_inst_o_src_a__2_ | decoded_inst_o_src_a__1_;
  assign N534 = N532 | N533;
  assign N535 = N534 | N531;
  assign N540 = N537 | N538;
  assign N541 = decoded_inst_o_src_a__2_ | N539;
  assign N542 = N540 | N541;
  assign N543 = N542 | decoded_inst_o_src_a__0_;
  assign N549 = N545 | N546;
  assign N550 = decoded_inst_o_src_a__2_ | N547;
  assign N551 = N549 | N550;
  assign N552 = N551 | N548;
  assign N557 = N554 | N555;
  assign N558 = N556 | decoded_inst_o_src_a__1_;
  assign N559 = N557 | N558;
  assign N560 = N559 | decoded_inst_o_src_a__0_;
  assign N566 = N562 | N563;
  assign N567 = N564 | decoded_inst_o_src_a__1_;
  assign N568 = N566 | N567;
  assign N569 = N568 | N565;
  assign N571 = decoded_inst_o_src_a__4_ & decoded_inst_o_src_a__2_;
  assign N572 = decoded_inst_o_src_a__1_ & decoded_inst_o_src_a__0_;
  assign N573 = N571 & N572;
  assign N574 = decoded_inst_o_src_a__4_ & decoded_inst_o_src_a__3_;
  assign N575 = decoded_inst_o_src_a__2_ & decoded_inst_o_src_a__1_;
  assign N576 = N574 & N575;
  assign N601 = N596 & N597;
  assign N602 = N598 & N599;
  assign N603 = N601 & N602;
  assign N604 = N603 & N600;
  assign N606 = decoded_inst_o_src_b__4_ | decoded_inst_o_src_b__3_;
  assign N607 = decoded_inst_o_src_b__2_ | decoded_inst_o_src_b__1_;
  assign N608 = N606 | N607;
  assign N609 = N608 | N605;
  assign N612 = decoded_inst_o_src_b__4_ | decoded_inst_o_src_b__3_;
  assign N613 = decoded_inst_o_src_b__2_ | N611;
  assign N614 = N612 | N613;
  assign N615 = N614 | decoded_inst_o_src_b__0_;
  assign N619 = decoded_inst_o_src_b__4_ | decoded_inst_o_src_b__3_;
  assign N620 = decoded_inst_o_src_b__2_ | N617;
  assign N621 = N619 | N620;
  assign N622 = N621 | N618;
  assign N625 = decoded_inst_o_src_b__4_ | decoded_inst_o_src_b__3_;
  assign N626 = N624 | decoded_inst_o_src_b__1_;
  assign N627 = N625 | N626;
  assign N628 = N627 | decoded_inst_o_src_b__0_;
  assign N632 = decoded_inst_o_src_b__4_ | decoded_inst_o_src_b__3_;
  assign N633 = N630 | decoded_inst_o_src_b__1_;
  assign N634 = N632 | N633;
  assign N635 = N634 | N631;
  assign N639 = decoded_inst_o_src_b__4_ | decoded_inst_o_src_b__3_;
  assign N640 = N637 | N638;
  assign N641 = N639 | N640;
  assign N642 = N641 | decoded_inst_o_src_b__0_;
  assign N647 = decoded_inst_o_src_b__4_ | decoded_inst_o_src_b__3_;
  assign N648 = N644 | N645;
  assign N649 = N647 | N648;
  assign N650 = N649 | N646;
  assign N653 = decoded_inst_o_src_b__4_ | N652;
  assign N654 = decoded_inst_o_src_b__2_ | decoded_inst_o_src_b__1_;
  assign N655 = N653 | N654;
  assign N656 = N655 | decoded_inst_o_src_b__0_;
  assign N660 = decoded_inst_o_src_b__4_ | N658;
  assign N661 = decoded_inst_o_src_b__2_ | decoded_inst_o_src_b__1_;
  assign N662 = N660 | N661;
  assign N663 = N662 | N659;
  assign N667 = decoded_inst_o_src_b__4_ | N665;
  assign N668 = decoded_inst_o_src_b__2_ | N666;
  assign N669 = N667 | N668;
  assign N670 = N669 | decoded_inst_o_src_b__0_;
  assign N675 = decoded_inst_o_src_b__4_ | N672;
  assign N676 = decoded_inst_o_src_b__2_ | N673;
  assign N677 = N675 | N676;
  assign N678 = N677 | N674;
  assign N682 = decoded_inst_o_src_b__4_ | N680;
  assign N683 = N681 | decoded_inst_o_src_b__1_;
  assign N684 = N682 | N683;
  assign N685 = N684 | decoded_inst_o_src_b__0_;
  assign N690 = decoded_inst_o_src_b__4_ | N687;
  assign N691 = N688 | decoded_inst_o_src_b__1_;
  assign N692 = N690 | N691;
  assign N693 = N692 | N689;
  assign N698 = decoded_inst_o_src_b__4_ | N695;
  assign N699 = N696 | N697;
  assign N700 = N698 | N699;
  assign N701 = N700 | decoded_inst_o_src_b__0_;
  assign N707 = decoded_inst_o_src_b__4_ | N703;
  assign N708 = N704 | N705;
  assign N709 = N707 | N708;
  assign N710 = N709 | N706;
  assign N713 = N712 | decoded_inst_o_src_b__3_;
  assign N714 = decoded_inst_o_src_b__2_ | decoded_inst_o_src_b__1_;
  assign N715 = N713 | N714;
  assign N716 = N715 | decoded_inst_o_src_b__0_;
  assign N720 = N718 | decoded_inst_o_src_b__3_;
  assign N721 = decoded_inst_o_src_b__2_ | decoded_inst_o_src_b__1_;
  assign N722 = N720 | N721;
  assign N723 = N722 | N719;
  assign N727 = N725 | decoded_inst_o_src_b__3_;
  assign N728 = decoded_inst_o_src_b__2_ | N726;
  assign N729 = N727 | N728;
  assign N730 = N729 | decoded_inst_o_src_b__0_;
  assign N735 = N732 | decoded_inst_o_src_b__3_;
  assign N736 = decoded_inst_o_src_b__2_ | N733;
  assign N737 = N735 | N736;
  assign N738 = N737 | N734;
  assign N742 = N740 | decoded_inst_o_src_b__3_;
  assign N743 = N741 | decoded_inst_o_src_b__1_;
  assign N744 = N742 | N743;
  assign N745 = N744 | decoded_inst_o_src_b__0_;
  assign N750 = N747 | decoded_inst_o_src_b__3_;
  assign N751 = N748 | decoded_inst_o_src_b__1_;
  assign N752 = N750 | N751;
  assign N753 = N752 | N749;
  assign N758 = N755 | decoded_inst_o_src_b__3_;
  assign N759 = N756 | N757;
  assign N760 = N758 | N759;
  assign N761 = N760 | decoded_inst_o_src_b__0_;
  assign N765 = N763 | N764;
  assign N766 = decoded_inst_o_src_b__2_ | decoded_inst_o_src_b__1_;
  assign N767 = N765 | N766;
  assign N768 = N767 | decoded_inst_o_src_b__0_;
  assign N773 = N770 | N771;
  assign N774 = decoded_inst_o_src_b__2_ | decoded_inst_o_src_b__1_;
  assign N775 = N773 | N774;
  assign N776 = N775 | N772;
  assign N781 = N778 | N779;
  assign N782 = decoded_inst_o_src_b__2_ | N780;
  assign N783 = N781 | N782;
  assign N784 = N783 | decoded_inst_o_src_b__0_;
  assign N790 = N786 | N787;
  assign N791 = decoded_inst_o_src_b__2_ | N788;
  assign N792 = N790 | N791;
  assign N793 = N792 | N789;
  assign N798 = N795 | N796;
  assign N799 = N797 | decoded_inst_o_src_b__1_;
  assign N800 = N798 | N799;
  assign N801 = N800 | decoded_inst_o_src_b__0_;
  assign N807 = N803 | N804;
  assign N808 = N805 | decoded_inst_o_src_b__1_;
  assign N809 = N807 | N808;
  assign N810 = N809 | N806;
  assign N812 = decoded_inst_o_src_b__4_ & decoded_inst_o_src_b__2_;
  assign N813 = decoded_inst_o_src_b__1_ & decoded_inst_o_src_b__0_;
  assign N814 = N812 & N813;
  assign N815 = decoded_inst_o_src_b__4_ & decoded_inst_o_src_b__3_;
  assign N816 = decoded_inst_o_src_b__2_ & decoded_inst_o_src_b__1_;
  assign N817 = N815 & N816;
  assign N819 = ~lce_cmd_o[32];
  assign N820 = N819 | lce_cmd_o[33];
  assign N821 = lce_cmd_o[31] | N820;
  assign N822 = ~N821;
  assign N823 = ~lce_cmd_o[33];
  assign N824 = lce_cmd_o[32] | N823;
  assign N825 = lce_cmd_o[31] | N824;
  assign N826 = ~N825;
  assign N827 = ~lce_cmd_o[33];
  assign N828 = ~lce_cmd_o[31];
  assign N829 = lce_cmd_o[32] | N827;
  assign N830 = N828 | N829;
  assign N831 = ~N830;
  assign { N193, N192, N191, N190, N189, N188, N187 } = gpr_r_o[5:0] + cce_id_i[0];
  assign { N200, N199, N198, N197, N196, N195, N194 } = gpr_r_o[21:16] + cce_id_i[0];
  assign { N207, N206, N205, N204, N203, N202, N201 } = gpr_r_o[37:32] + cce_id_i[0];
  assign { N214, N213, N212, N211, N210, N209, N208 } = gpr_r_o[53:48] + cce_id_i[0];
  assign lce_cmd_o[35] = (N1)? gpr_r_o[0] :
                         (N2)? gpr_r_o[16] :
                         (N3)? gpr_r_o[32] :
                         (N4)? gpr_r_o[48] :
                         (N5)? lce_data_cmd_o[5] :
                         (N6)? mem_data_cmd_o[520] :
                         (N7)? 1'b0 :
                         (N8)? 1'b0 : 1'b0;
  assign N1 = N123;
  assign N2 = N127;
  assign N3 = N131;
  assign N4 = N136;
  assign N5 = N140;
  assign N6 = N145;
  assign N7 = N150;
  assign N8 = N152;
  assign lce_cmd_o[30:9] = (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N193, N192, N191, N190, N189, N188, N187, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                           (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N200, N199, N198, N197, N196, N195, N194, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                           (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N207, N206, N205, N204, N203, N202, N201, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                           (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N214, N213, N212, N211, N210, N209, N208, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                           (N13)? mem_cmd_o[28:7] :
                           (N14)? lru_addr_r_o :
                           (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                           (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N9 = N157;
  assign N10 = N161;
  assign N11 = N165;
  assign N12 = N170;
  assign N13 = N174;
  assign N14 = N179;
  assign N15 = N184;
  assign N16 = N186;
  assign lce_cmd_o[8:6] = (N17)? req_addr_way_r_o :
                          (N18)? mem_data_cmd_o[519:517] :
                          (N19)? { N241, N242, N243 } :
                          (N20)? mem_cmd_o[5:3] :
                          (N21)? { 1'b0, 1'b0, 1'b0 } :
                          (N22)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N17 = N219;
  assign N18 = N223;
  assign N19 = N227;
  assign N20 = N232;
  assign N21 = N236;
  assign N22 = N239;
  assign mem_data_cmd_o[568:547] = (N23)? lru_addr_r_o :
                                   (N24)? mem_cmd_o[28:7] : 1'b0;
  assign N23 = N244;
  assign N24 = N245;
  assign lce_cmd_o[5:4] = (N25)? next_coh_state_r_o :
                          (N247)? { 1'b0, 1'b0 } : 1'b0;
  assign N25 = N246;
  assign lce_cmd_o[3:0] = (N26)? { lce_data_cmd_o[5:5], mem_cmd_o[5:3] } :
                          (N27)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N26 = N822;
  assign N27 = N821;
  assign lce_data_cmd_o[3] = ~lce_data_cmd_o[4];
  assign { lce_data_cmd_o[517:6], lce_data_cmd_o[2:0] } = (N28)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, nc_data_r_o, 1'b0, 1'b0, 1'b0 } :
                                                          (N248)? { cache_block_data_r_o, mem_cmd_o[5:3] } : 1'b0;
  assign N28 = lce_data_cmd_o[4];
  assign mem_data_cmd_o[511:0] = (N29)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, nc_data_r_o } :
                                 (N249)? cache_block_data_r_o : 1'b0;
  assign N29 = mem_cmd_o[2];
  assign dir_way_group_i = (N30)? gpr_r_o[5:0] :
                           (N31)? gpr_r_o[21:16] :
                           (N32)? gpr_r_o[37:32] :
                           (N33)? gpr_r_o[53:48] :
                           (N34)? mem_cmd_o[18:13] :
                           (N35)? lru_addr_r_o[11:6] :
                           (N36)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N30 = N254;
  assign N31 = N258;
  assign N32 = N262;
  assign N33 = N267;
  assign N34 = N271;
  assign N35 = N276;
  assign N36 = N277;
  assign dir_lce_i[0] = (N37)? gpr_r_o[0] :
                        (N38)? gpr_r_o[16] :
                        (N39)? gpr_r_o[32] :
                        (N40)? gpr_r_o[48] :
                        (N41)? lce_data_cmd_o[5] :
                        (N42)? mem_data_cmd_o[520] :
                        (N43)? 1'b0 : 1'b0;
  assign N37 = N282;
  assign N38 = N286;
  assign N39 = N290;
  assign N40 = N295;
  assign N41 = N299;
  assign N42 = N304;
  assign N43 = N305;
  assign dir_way_i = (N44)? gpr_r_o[2:0] :
                     (N45)? gpr_r_o[18:16] :
                     (N46)? gpr_r_o[34:32] :
                     (N47)? gpr_r_o[50:48] :
                     (N48)? req_addr_way_r_o :
                     (N49)? mem_cmd_o[5:3] :
                     (N50)? { N340, N341, N342 } :
                     (N51)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N44 = N310;
  assign N45 = N314;
  assign N46 = N318;
  assign N47 = N323;
  assign N48 = N327;
  assign N49 = N332;
  assign N50 = N337;
  assign N51 = N339;
  assign dir_coh_state_i = (N52)? next_coh_state_r_o :
                           (N53)? { decoded_inst_o_imm__1_, decoded_inst_o_imm__0_ } : 1'b0;
  assign N52 = N343;
  assign N53 = N344;
  assign dir_tag_i = (N54)? mem_cmd_o[28:19] :
                     (N55)? lru_addr_r_o[21:12] :
                     (N56)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                     (N57)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N54 = N347;
  assign N55 = N350;
  assign N56 = N353;
  assign N57 = N354;
  assign { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } = (N58)? gpr_r_o[15:0] :
                                                                                                              (N59)? gpr_r_o[31:16] :
                                                                                                              (N60)? gpr_r_o[47:32] :
                                                                                                              (N61)? gpr_r_o[63:48] :
                                                                                                              (N62)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_cmd_o[29:29] } :
                                                                                                              (N63)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o_1 } :
                                                                                                              (N64)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o_2 } :
                                                                                                              (N65)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o_3 } :
                                                                                                              (N66)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_data_cmd_o[516:516] } :
                                                                                                              (N67)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_data_cmd_o[515:515] } :
                                                                                                              (N68)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o[6:6] } :
                                                                                                              (N69)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o[7:7] } :
                                                                                                              (N70)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o[8:8] } :
                                                                                                              (N71)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o[9:9] } :
                                                                                                              (N72)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o[10:10] } :
                                                                                                              (N73)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o[11:11] } :
                                                                                                              (N74)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_cmd_o[2:2] } :
                                                                                                              (N75)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                              (N76)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } :
                                                                                                              (N77)? { decoded_inst_o_imm__15_, decoded_inst_o_imm__14_, decoded_inst_o_imm__13_, decoded_inst_o_imm__12_, decoded_inst_o_imm__11_, decoded_inst_o_imm__10_, decoded_inst_o_imm__9_, decoded_inst_o_imm__8_, decoded_inst_o_imm__7_, decoded_inst_o_imm__6_, decoded_inst_o_imm__5_, decoded_inst_o_imm__4_, decoded_inst_o_imm__3_, decoded_inst_o_imm__2_, decoded_inst_o_imm__1_, decoded_inst_o_imm__0_ } :
                                                                                                              (N78)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_data_cmd_o[5:5] } :
                                                                                                              (N79)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, ack_type_r_o } :
                                                                                                              (N80)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sharers_hits_r0 } :
                                                                                                              (N81)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_req_v_i } :
                                                                                                              (N82)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_resp_v_i } :
                                                                                                              (N83)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_data_resp_v_i } :
                                                                                                              (N84)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                                                                                                              (N85)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_resp_v_i } :
                                                                                                              (N86)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_data_resp_v_i } :
                                                                                                              (N87)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N58 = N363;
  assign N59 = N369;
  assign N60 = N375;
  assign N61 = N382;
  assign N62 = N388;
  assign N63 = N395;
  assign N64 = N402;
  assign N65 = N410;
  assign N66 = N416;
  assign N67 = N423;
  assign N68 = N430;
  assign N69 = N438;
  assign N70 = N445;
  assign N71 = N453;
  assign N72 = N461;
  assign N73 = N470;
  assign N74 = N476;
  assign N75 = N483;
  assign N76 = N490;
  assign N77 = N498;
  assign N78 = N505;
  assign N79 = N513;
  assign N80 = N521;
  assign N81 = N528;
  assign N82 = N536;
  assign N83 = N544;
  assign N84 = N553;
  assign N85 = N561;
  assign N86 = N570;
  assign N87 = N577;
  assign mov_src = (N88)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                   (N595)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N88 = N594;
  assign alu_opd_b_i = (N89)? gpr_r_o[15:0] :
                       (N90)? gpr_r_o[31:16] :
                       (N91)? gpr_r_o[47:32] :
                       (N92)? gpr_r_o[63:48] :
                       (N93)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_cmd_o[29:29] } :
                       (N94)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o_1 } :
                       (N95)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o_2 } :
                       (N96)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o_3 } :
                       (N97)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_data_cmd_o[516:516] } :
                       (N98)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_data_cmd_o[515:515] } :
                       (N99)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o[6:6] } :
                       (N100)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o[7:7] } :
                       (N101)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o[8:8] } :
                       (N102)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o[9:9] } :
                       (N103)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o[10:10] } :
                       (N104)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flags_r_o[11:11] } :
                       (N105)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_cmd_o[2:2] } :
                       (N106)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                       (N107)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } :
                       (N108)? { decoded_inst_o_imm__15_, decoded_inst_o_imm__14_, decoded_inst_o_imm__13_, decoded_inst_o_imm__12_, decoded_inst_o_imm__11_, decoded_inst_o_imm__10_, decoded_inst_o_imm__9_, decoded_inst_o_imm__8_, decoded_inst_o_imm__7_, decoded_inst_o_imm__6_, decoded_inst_o_imm__5_, decoded_inst_o_imm__4_, decoded_inst_o_imm__3_, decoded_inst_o_imm__2_, decoded_inst_o_imm__1_, decoded_inst_o_imm__0_ } :
                       (N109)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_data_cmd_o[5:5] } :
                       (N110)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, ack_type_r_o } :
                       (N111)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sharers_hits_r0 } :
                       (N112)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_req_v_i } :
                       (N113)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_resp_v_i } :
                       (N114)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_data_resp_v_i } :
                       (N115)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                       (N116)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                       (N117)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } :
                       (N118)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N89 = N604;
  assign N90 = N610;
  assign N91 = N616;
  assign N92 = N623;
  assign N93 = N629;
  assign N94 = N636;
  assign N95 = N643;
  assign N96 = N651;
  assign N97 = N657;
  assign N98 = N664;
  assign N99 = N671;
  assign N100 = N679;
  assign N101 = N686;
  assign N102 = N694;
  assign N103 = N702;
  assign N104 = N711;
  assign N105 = N717;
  assign N106 = N724;
  assign N107 = N731;
  assign N108 = N739;
  assign N109 = N746;
  assign N110 = N754;
  assign N111 = N762;
  assign N112 = N769;
  assign N113 = N777;
  assign N114 = N785;
  assign N115 = N794;
  assign N116 = N802;
  assign N117 = N811;
  assign N118 = N818;
  assign alu_opd_a_i = (N89)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N90)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N91)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N92)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N93)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N94)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N95)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N96)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N97)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N98)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N99)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N100)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N101)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N102)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N103)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N104)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N105)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N106)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N107)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N108)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N109)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N110)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N111)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N112)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N113)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N114)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N115)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } :
                       (N116)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_resp_v_i } :
                       (N117)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_data_resp_v_i } :
                       (N118)? { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578 } : 1'b0;
  assign gad_v_i = decoded_inst_v_o & decoded_inst_o_gad_op_w_v_;
  assign N119 = ~decoded_inst_o_lce_cmd_lce_sel__2_;
  assign N120 = ~decoded_inst_o_lce_cmd_lce_sel__1_;
  assign N121 = ~decoded_inst_o_lce_cmd_lce_sel__0_;
  assign N124 = ~decoded_inst_o_lce_cmd_lce_sel__0_;
  assign N127 = ~N126;
  assign N128 = ~decoded_inst_o_lce_cmd_lce_sel__1_;
  assign N131 = ~N130;
  assign N132 = ~decoded_inst_o_lce_cmd_lce_sel__1_;
  assign N133 = ~decoded_inst_o_lce_cmd_lce_sel__0_;
  assign N136 = ~N135;
  assign N137 = ~decoded_inst_o_lce_cmd_lce_sel__2_;
  assign N140 = ~N139;
  assign N141 = ~decoded_inst_o_lce_cmd_lce_sel__2_;
  assign N142 = ~decoded_inst_o_lce_cmd_lce_sel__0_;
  assign N145 = ~N144;
  assign N146 = ~decoded_inst_o_lce_cmd_lce_sel__2_;
  assign N147 = ~decoded_inst_o_lce_cmd_lce_sel__1_;
  assign N150 = ~N149;
  assign N153 = ~decoded_inst_o_lce_cmd_addr_sel__2_;
  assign N154 = ~decoded_inst_o_lce_cmd_addr_sel__1_;
  assign N155 = ~decoded_inst_o_lce_cmd_addr_sel__0_;
  assign N158 = ~decoded_inst_o_lce_cmd_addr_sel__0_;
  assign N161 = ~N160;
  assign N162 = ~decoded_inst_o_lce_cmd_addr_sel__1_;
  assign N165 = ~N164;
  assign N166 = ~decoded_inst_o_lce_cmd_addr_sel__1_;
  assign N167 = ~decoded_inst_o_lce_cmd_addr_sel__0_;
  assign N170 = ~N169;
  assign N171 = ~decoded_inst_o_lce_cmd_addr_sel__2_;
  assign N174 = ~N173;
  assign N175 = ~decoded_inst_o_lce_cmd_addr_sel__2_;
  assign N176 = ~decoded_inst_o_lce_cmd_addr_sel__0_;
  assign N179 = ~N178;
  assign N180 = ~decoded_inst_o_lce_cmd_addr_sel__2_;
  assign N181 = ~decoded_inst_o_lce_cmd_addr_sel__1_;
  assign N184 = ~N183;
  assign N215 = ~decoded_inst_o_lce_cmd_way_sel__2_;
  assign N216 = ~decoded_inst_o_lce_cmd_way_sel__1_;
  assign N217 = ~decoded_inst_o_lce_cmd_way_sel__0_;
  assign N220 = ~decoded_inst_o_lce_cmd_way_sel__0_;
  assign N223 = ~N222;
  assign N224 = ~decoded_inst_o_lce_cmd_way_sel__1_;
  assign N227 = ~N226;
  assign N228 = ~decoded_inst_o_lce_cmd_way_sel__1_;
  assign N229 = ~decoded_inst_o_lce_cmd_way_sel__0_;
  assign N232 = ~N231;
  assign N233 = ~decoded_inst_o_lce_cmd_way_sel__2_;
  assign N236 = ~N235;
  assign N239 = N237 | N238;
  assign N240 = ~gpr_r_o[0];
  assign N244 = ~decoded_inst_o_mem_data_cmd_addr_sel_;
  assign N245 = decoded_inst_o_mem_data_cmd_addr_sel_;
  assign N246 = N826 | N831;
  assign N247 = ~N246;
  assign lce_data_cmd_o[4] = mem_cmd_o[2];
  assign N248 = ~lce_data_cmd_o[4];
  assign N249 = ~mem_cmd_o[2];
  assign N250 = ~decoded_inst_o_dir_way_group_sel__2_;
  assign N251 = ~decoded_inst_o_dir_way_group_sel__1_;
  assign N252 = ~decoded_inst_o_dir_way_group_sel__0_;
  assign N255 = ~decoded_inst_o_dir_way_group_sel__0_;
  assign N258 = ~N257;
  assign N259 = ~decoded_inst_o_dir_way_group_sel__1_;
  assign N262 = ~N261;
  assign N263 = ~decoded_inst_o_dir_way_group_sel__1_;
  assign N264 = ~decoded_inst_o_dir_way_group_sel__0_;
  assign N267 = ~N266;
  assign N268 = ~decoded_inst_o_dir_way_group_sel__2_;
  assign N271 = ~N270;
  assign N272 = ~decoded_inst_o_dir_way_group_sel__2_;
  assign N273 = ~decoded_inst_o_dir_way_group_sel__0_;
  assign N276 = ~N275;
  assign N278 = ~decoded_inst_o_dir_lce_sel__2_;
  assign N279 = ~decoded_inst_o_dir_lce_sel__1_;
  assign N280 = ~decoded_inst_o_dir_lce_sel__0_;
  assign N283 = ~decoded_inst_o_dir_lce_sel__0_;
  assign N286 = ~N285;
  assign N287 = ~decoded_inst_o_dir_lce_sel__1_;
  assign N290 = ~N289;
  assign N291 = ~decoded_inst_o_dir_lce_sel__1_;
  assign N292 = ~decoded_inst_o_dir_lce_sel__0_;
  assign N295 = ~N294;
  assign N296 = ~decoded_inst_o_dir_lce_sel__2_;
  assign N299 = ~N298;
  assign N300 = ~decoded_inst_o_dir_lce_sel__2_;
  assign N301 = ~decoded_inst_o_dir_lce_sel__0_;
  assign N304 = ~N303;
  assign N306 = ~decoded_inst_o_dir_way_sel__2_;
  assign N307 = ~decoded_inst_o_dir_way_sel__1_;
  assign N308 = ~decoded_inst_o_dir_way_sel__0_;
  assign N311 = ~decoded_inst_o_dir_way_sel__0_;
  assign N314 = ~N313;
  assign N315 = ~decoded_inst_o_dir_way_sel__1_;
  assign N318 = ~N317;
  assign N319 = ~decoded_inst_o_dir_way_sel__1_;
  assign N320 = ~decoded_inst_o_dir_way_sel__0_;
  assign N323 = ~N322;
  assign N324 = ~decoded_inst_o_dir_way_sel__2_;
  assign N327 = ~N326;
  assign N328 = ~decoded_inst_o_dir_way_sel__2_;
  assign N329 = ~decoded_inst_o_dir_way_sel__0_;
  assign N332 = ~N331;
  assign N333 = ~decoded_inst_o_dir_way_sel__2_;
  assign N334 = ~decoded_inst_o_dir_way_sel__1_;
  assign N337 = ~N336;
  assign N343 = ~decoded_inst_o_dir_coh_state_sel_;
  assign N344 = decoded_inst_o_dir_coh_state_sel_;
  assign N345 = ~decoded_inst_o_dir_tag_sel__1_;
  assign N346 = ~decoded_inst_o_dir_tag_sel__0_;
  assign N348 = ~decoded_inst_o_dir_tag_sel__0_;
  assign N350 = ~N349;
  assign N351 = ~decoded_inst_o_dir_tag_sel__1_;
  assign N353 = ~N352;
  assign N355 = ~decoded_inst_o_src_a__4_;
  assign N356 = ~decoded_inst_o_src_a__3_;
  assign N357 = ~decoded_inst_o_src_a__2_;
  assign N358 = ~decoded_inst_o_src_a__1_;
  assign N359 = ~decoded_inst_o_src_a__0_;
  assign N364 = ~decoded_inst_o_src_a__0_;
  assign N369 = ~N368;
  assign N370 = ~decoded_inst_o_src_a__1_;
  assign N375 = ~N374;
  assign N376 = ~decoded_inst_o_src_a__1_;
  assign N377 = ~decoded_inst_o_src_a__0_;
  assign N382 = ~N381;
  assign N383 = ~decoded_inst_o_src_a__2_;
  assign N388 = ~N387;
  assign N389 = ~decoded_inst_o_src_a__2_;
  assign N390 = ~decoded_inst_o_src_a__0_;
  assign N395 = ~N394;
  assign N396 = ~decoded_inst_o_src_a__2_;
  assign N397 = ~decoded_inst_o_src_a__1_;
  assign N402 = ~N401;
  assign N403 = ~decoded_inst_o_src_a__2_;
  assign N404 = ~decoded_inst_o_src_a__1_;
  assign N405 = ~decoded_inst_o_src_a__0_;
  assign N410 = ~N409;
  assign N411 = ~decoded_inst_o_src_a__3_;
  assign N416 = ~N415;
  assign N417 = ~decoded_inst_o_src_a__3_;
  assign N418 = ~decoded_inst_o_src_a__0_;
  assign N423 = ~N422;
  assign N424 = ~decoded_inst_o_src_a__3_;
  assign N425 = ~decoded_inst_o_src_a__1_;
  assign N430 = ~N429;
  assign N431 = ~decoded_inst_o_src_a__3_;
  assign N432 = ~decoded_inst_o_src_a__1_;
  assign N433 = ~decoded_inst_o_src_a__0_;
  assign N438 = ~N437;
  assign N439 = ~decoded_inst_o_src_a__3_;
  assign N440 = ~decoded_inst_o_src_a__2_;
  assign N445 = ~N444;
  assign N446 = ~decoded_inst_o_src_a__3_;
  assign N447 = ~decoded_inst_o_src_a__2_;
  assign N448 = ~decoded_inst_o_src_a__0_;
  assign N453 = ~N452;
  assign N454 = ~decoded_inst_o_src_a__3_;
  assign N455 = ~decoded_inst_o_src_a__2_;
  assign N456 = ~decoded_inst_o_src_a__1_;
  assign N461 = ~N460;
  assign N462 = ~decoded_inst_o_src_a__3_;
  assign N463 = ~decoded_inst_o_src_a__2_;
  assign N464 = ~decoded_inst_o_src_a__1_;
  assign N465 = ~decoded_inst_o_src_a__0_;
  assign N470 = ~N469;
  assign N471 = ~decoded_inst_o_src_a__4_;
  assign N476 = ~N475;
  assign N477 = ~decoded_inst_o_src_a__4_;
  assign N478 = ~decoded_inst_o_src_a__0_;
  assign N483 = ~N482;
  assign N484 = ~decoded_inst_o_src_a__4_;
  assign N485 = ~decoded_inst_o_src_a__1_;
  assign N490 = ~N489;
  assign N491 = ~decoded_inst_o_src_a__4_;
  assign N492 = ~decoded_inst_o_src_a__1_;
  assign N493 = ~decoded_inst_o_src_a__0_;
  assign N498 = ~N497;
  assign N499 = ~decoded_inst_o_src_a__4_;
  assign N500 = ~decoded_inst_o_src_a__2_;
  assign N505 = ~N504;
  assign N506 = ~decoded_inst_o_src_a__4_;
  assign N507 = ~decoded_inst_o_src_a__2_;
  assign N508 = ~decoded_inst_o_src_a__0_;
  assign N513 = ~N512;
  assign N514 = ~decoded_inst_o_src_a__4_;
  assign N515 = ~decoded_inst_o_src_a__2_;
  assign N516 = ~decoded_inst_o_src_a__1_;
  assign N521 = ~N520;
  assign N522 = ~decoded_inst_o_src_a__4_;
  assign N523 = ~decoded_inst_o_src_a__3_;
  assign N528 = ~N527;
  assign N529 = ~decoded_inst_o_src_a__4_;
  assign N530 = ~decoded_inst_o_src_a__3_;
  assign N531 = ~decoded_inst_o_src_a__0_;
  assign N536 = ~N535;
  assign N537 = ~decoded_inst_o_src_a__4_;
  assign N538 = ~decoded_inst_o_src_a__3_;
  assign N539 = ~decoded_inst_o_src_a__1_;
  assign N544 = ~N543;
  assign N545 = ~decoded_inst_o_src_a__4_;
  assign N546 = ~decoded_inst_o_src_a__3_;
  assign N547 = ~decoded_inst_o_src_a__1_;
  assign N548 = ~decoded_inst_o_src_a__0_;
  assign N553 = ~N552;
  assign N554 = ~decoded_inst_o_src_a__4_;
  assign N555 = ~decoded_inst_o_src_a__3_;
  assign N556 = ~decoded_inst_o_src_a__2_;
  assign N561 = ~N560;
  assign N562 = ~decoded_inst_o_src_a__4_;
  assign N563 = ~decoded_inst_o_src_a__3_;
  assign N564 = ~decoded_inst_o_src_a__2_;
  assign N565 = ~decoded_inst_o_src_a__0_;
  assign N570 = ~N569;
  assign N577 = N573 | N576;
  assign N594 = decoded_inst_o_mov_dst_w_v_;
  assign N595 = ~N594;
  assign N596 = ~decoded_inst_o_src_b__4_;
  assign N597 = ~decoded_inst_o_src_b__3_;
  assign N598 = ~decoded_inst_o_src_b__2_;
  assign N599 = ~decoded_inst_o_src_b__1_;
  assign N600 = ~decoded_inst_o_src_b__0_;
  assign N605 = ~decoded_inst_o_src_b__0_;
  assign N610 = ~N609;
  assign N611 = ~decoded_inst_o_src_b__1_;
  assign N616 = ~N615;
  assign N617 = ~decoded_inst_o_src_b__1_;
  assign N618 = ~decoded_inst_o_src_b__0_;
  assign N623 = ~N622;
  assign N624 = ~decoded_inst_o_src_b__2_;
  assign N629 = ~N628;
  assign N630 = ~decoded_inst_o_src_b__2_;
  assign N631 = ~decoded_inst_o_src_b__0_;
  assign N636 = ~N635;
  assign N637 = ~decoded_inst_o_src_b__2_;
  assign N638 = ~decoded_inst_o_src_b__1_;
  assign N643 = ~N642;
  assign N644 = ~decoded_inst_o_src_b__2_;
  assign N645 = ~decoded_inst_o_src_b__1_;
  assign N646 = ~decoded_inst_o_src_b__0_;
  assign N651 = ~N650;
  assign N652 = ~decoded_inst_o_src_b__3_;
  assign N657 = ~N656;
  assign N658 = ~decoded_inst_o_src_b__3_;
  assign N659 = ~decoded_inst_o_src_b__0_;
  assign N664 = ~N663;
  assign N665 = ~decoded_inst_o_src_b__3_;
  assign N666 = ~decoded_inst_o_src_b__1_;
  assign N671 = ~N670;
  assign N672 = ~decoded_inst_o_src_b__3_;
  assign N673 = ~decoded_inst_o_src_b__1_;
  assign N674 = ~decoded_inst_o_src_b__0_;
  assign N679 = ~N678;
  assign N680 = ~decoded_inst_o_src_b__3_;
  assign N681 = ~decoded_inst_o_src_b__2_;
  assign N686 = ~N685;
  assign N687 = ~decoded_inst_o_src_b__3_;
  assign N688 = ~decoded_inst_o_src_b__2_;
  assign N689 = ~decoded_inst_o_src_b__0_;
  assign N694 = ~N693;
  assign N695 = ~decoded_inst_o_src_b__3_;
  assign N696 = ~decoded_inst_o_src_b__2_;
  assign N697 = ~decoded_inst_o_src_b__1_;
  assign N702 = ~N701;
  assign N703 = ~decoded_inst_o_src_b__3_;
  assign N704 = ~decoded_inst_o_src_b__2_;
  assign N705 = ~decoded_inst_o_src_b__1_;
  assign N706 = ~decoded_inst_o_src_b__0_;
  assign N711 = ~N710;
  assign N712 = ~decoded_inst_o_src_b__4_;
  assign N717 = ~N716;
  assign N718 = ~decoded_inst_o_src_b__4_;
  assign N719 = ~decoded_inst_o_src_b__0_;
  assign N724 = ~N723;
  assign N725 = ~decoded_inst_o_src_b__4_;
  assign N726 = ~decoded_inst_o_src_b__1_;
  assign N731 = ~N730;
  assign N732 = ~decoded_inst_o_src_b__4_;
  assign N733 = ~decoded_inst_o_src_b__1_;
  assign N734 = ~decoded_inst_o_src_b__0_;
  assign N739 = ~N738;
  assign N740 = ~decoded_inst_o_src_b__4_;
  assign N741 = ~decoded_inst_o_src_b__2_;
  assign N746 = ~N745;
  assign N747 = ~decoded_inst_o_src_b__4_;
  assign N748 = ~decoded_inst_o_src_b__2_;
  assign N749 = ~decoded_inst_o_src_b__0_;
  assign N754 = ~N753;
  assign N755 = ~decoded_inst_o_src_b__4_;
  assign N756 = ~decoded_inst_o_src_b__2_;
  assign N757 = ~decoded_inst_o_src_b__1_;
  assign N762 = ~N761;
  assign N763 = ~decoded_inst_o_src_b__4_;
  assign N764 = ~decoded_inst_o_src_b__3_;
  assign N769 = ~N768;
  assign N770 = ~decoded_inst_o_src_b__4_;
  assign N771 = ~decoded_inst_o_src_b__3_;
  assign N772 = ~decoded_inst_o_src_b__0_;
  assign N777 = ~N776;
  assign N778 = ~decoded_inst_o_src_b__4_;
  assign N779 = ~decoded_inst_o_src_b__3_;
  assign N780 = ~decoded_inst_o_src_b__1_;
  assign N785 = ~N784;
  assign N786 = ~decoded_inst_o_src_b__4_;
  assign N787 = ~decoded_inst_o_src_b__3_;
  assign N788 = ~decoded_inst_o_src_b__1_;
  assign N789 = ~decoded_inst_o_src_b__0_;
  assign N794 = ~N793;
  assign N795 = ~decoded_inst_o_src_b__4_;
  assign N796 = ~decoded_inst_o_src_b__3_;
  assign N797 = ~decoded_inst_o_src_b__2_;
  assign N802 = ~N801;
  assign N803 = ~decoded_inst_o_src_b__4_;
  assign N804 = ~decoded_inst_o_src_b__3_;
  assign N805 = ~decoded_inst_o_src_b__2_;
  assign N806 = ~decoded_inst_o_src_b__0_;
  assign N811 = ~N810;
  assign N818 = N814 | N817;

endmodule



module bp_cce_top_num_lce_p2_num_cce_p1_paddr_width_p22_lce_assoc_p8_lce_sets_p64_block_size_in_bytes_p64_num_cce_inst_ram_els_p256_lce_req_data_width_p64
(
  clk_i,
  reset_i,
  lce_req_i,
  lce_req_v_i,
  lce_req_ready_o,
  lce_resp_i,
  lce_resp_v_i,
  lce_resp_ready_o,
  lce_data_resp_i,
  lce_data_resp_v_i,
  lce_data_resp_ready_o,
  lce_cmd_o,
  lce_cmd_v_o,
  lce_cmd_ready_i,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i,
  mem_resp_i,
  mem_resp_v_i,
  mem_resp_ready_o,
  mem_data_resp_i,
  mem_data_resp_v_i,
  mem_data_resp_ready_o,
  mem_cmd_o,
  mem_cmd_v_o,
  mem_cmd_yumi_i,
  mem_data_cmd_o,
  mem_data_cmd_v_o,
  mem_data_cmd_yumi_i,
  cce_id_i,
  boot_rom_addr_o,
  boot_rom_data_i
);

  input [96:0] lce_req_i;
  input [25:0] lce_resp_i;
  input [536:0] lce_data_resp_i;
  output [35:0] lce_cmd_o;
  output [517:0] lce_data_cmd_o;
  input [57:0] mem_resp_i;
  input [541:0] mem_data_resp_i;
  output [29:0] mem_cmd_o;
  output [569:0] mem_data_cmd_o;
  input [0:0] cce_id_i;
  output [7:0] boot_rom_addr_o;
  input [95:0] boot_rom_data_i;
  input clk_i;
  input reset_i;
  input lce_req_v_i;
  input lce_resp_v_i;
  input lce_data_resp_v_i;
  input lce_cmd_ready_i;
  input lce_data_cmd_ready_i;
  input mem_resp_v_i;
  input mem_data_resp_v_i;
  input mem_cmd_yumi_i;
  input mem_data_cmd_yumi_i;
  output lce_req_ready_o;
  output lce_resp_ready_o;
  output lce_data_resp_ready_o;
  output lce_cmd_v_o;
  output lce_data_cmd_v_o;
  output mem_resp_ready_o;
  output mem_data_resp_ready_o;
  output mem_cmd_v_o;
  output mem_data_cmd_v_o;
  wire [35:0] lce_cmd_o;
  wire [517:0] lce_data_cmd_o;
  wire [29:0] mem_cmd_o,mem_cmd_from_cce;
  wire [569:0] mem_data_cmd_o,mem_data_cmd_from_cce;
  wire [7:0] boot_rom_addr_o;
  wire lce_req_ready_o,lce_resp_ready_o,lce_data_resp_ready_o,lce_cmd_v_o,
  lce_data_cmd_v_o,mem_resp_ready_o,mem_data_resp_ready_o,mem_cmd_v_o,mem_data_cmd_v_o,
  lce_req_v_to_cce,lce_req_yumi_from_cce,lce_resp_v_to_cce,lce_resp_yumi_from_cce,
  lce_data_resp_v_to_cce,lce_data_resp_yumi_from_cce,mem_resp_v_to_cce,
  mem_resp_yumi_from_cce,mem_data_resp_v_to_cce,mem_data_resp_yumi_from_cce,mem_cmd_v_from_cce,
  mem_cmd_ready_to_cce,mem_data_cmd_v_from_cce,mem_data_cmd_ready_to_cce;
  wire [96:0] lce_req_to_cce;
  wire [25:0] lce_resp_to_cce;
  wire [536:0] lce_data_resp_to_cce;
  wire [57:0] mem_resp_to_cce;
  wire [541:0] mem_data_resp_to_cce;

  bsg_two_fifo_width_p97
  lce_cce_req_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(lce_req_ready_o),
    .data_i(lce_req_i),
    .v_i(lce_req_v_i),
    .v_o(lce_req_v_to_cce),
    .data_o(lce_req_to_cce),
    .yumi_i(lce_req_yumi_from_cce)
  );


  bsg_two_fifo_width_p26
  lce_cce_resp_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(lce_resp_ready_o),
    .data_i(lce_resp_i),
    .v_i(lce_resp_v_i),
    .v_o(lce_resp_v_to_cce),
    .data_o(lce_resp_to_cce),
    .yumi_i(lce_resp_yumi_from_cce)
  );


  bsg_two_fifo_width_p537
  lce_cce_data_resp_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(lce_data_resp_ready_o),
    .data_i(lce_data_resp_i),
    .v_i(lce_data_resp_v_i),
    .v_o(lce_data_resp_v_to_cce),
    .data_o(lce_data_resp_to_cce),
    .yumi_i(lce_data_resp_yumi_from_cce)
  );


  bsg_two_fifo_width_p58
  mem_cce_resp_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(mem_resp_ready_o),
    .data_i(mem_resp_i),
    .v_i(mem_resp_v_i),
    .v_o(mem_resp_v_to_cce),
    .data_o(mem_resp_to_cce),
    .yumi_i(mem_resp_yumi_from_cce)
  );


  bsg_two_fifo_width_p542
  mem_cce_data_resp_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(mem_data_resp_ready_o),
    .data_i(mem_data_resp_i),
    .v_i(mem_data_resp_v_i),
    .v_o(mem_data_resp_v_to_cce),
    .data_o(mem_data_resp_to_cce),
    .yumi_i(mem_data_resp_yumi_from_cce)
  );


  bsg_two_fifo_width_p30
  cce_mem_cmd_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(mem_cmd_ready_to_cce),
    .data_i(mem_cmd_from_cce),
    .v_i(mem_cmd_v_from_cce),
    .v_o(mem_cmd_v_o),
    .data_o(mem_cmd_o),
    .yumi_i(mem_cmd_yumi_i)
  );


  bsg_two_fifo_width_p570
  cce_mem_data_cmd_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(mem_data_cmd_ready_to_cce),
    .data_i(mem_data_cmd_from_cce),
    .v_i(mem_data_cmd_v_from_cce),
    .v_o(mem_data_cmd_v_o),
    .data_o(mem_data_cmd_o),
    .yumi_i(mem_data_cmd_yumi_i)
  );


  bp_cce_num_lce_p2_num_cce_p1_paddr_width_p22_lce_assoc_p8_lce_sets_p64_block_size_in_bytes_p64_num_cce_inst_ram_els_p256_lce_req_data_width_p64
  bp_cce
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .lce_req_i(lce_req_to_cce),
    .lce_req_v_i(lce_req_v_to_cce),
    .lce_req_yumi_o(lce_req_yumi_from_cce),
    .lce_resp_i(lce_resp_to_cce),
    .lce_resp_v_i(lce_resp_v_to_cce),
    .lce_resp_yumi_o(lce_resp_yumi_from_cce),
    .lce_data_resp_i(lce_data_resp_to_cce),
    .lce_data_resp_v_i(lce_data_resp_v_to_cce),
    .lce_data_resp_yumi_o(lce_data_resp_yumi_from_cce),
    .lce_cmd_o(lce_cmd_o),
    .lce_cmd_v_o(lce_cmd_v_o),
    .lce_cmd_ready_i(lce_cmd_ready_i),
    .lce_data_cmd_o(lce_data_cmd_o),
    .lce_data_cmd_v_o(lce_data_cmd_v_o),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_i),
    .mem_resp_i(mem_resp_to_cce),
    .mem_resp_v_i(mem_resp_v_to_cce),
    .mem_resp_yumi_o(mem_resp_yumi_from_cce),
    .mem_data_resp_i(mem_data_resp_to_cce),
    .mem_data_resp_v_i(mem_data_resp_v_to_cce),
    .mem_data_resp_yumi_o(mem_data_resp_yumi_from_cce),
    .mem_cmd_o(mem_cmd_from_cce),
    .mem_cmd_v_o(mem_cmd_v_from_cce),
    .mem_cmd_ready_i(mem_cmd_ready_to_cce),
    .mem_data_cmd_o(mem_data_cmd_from_cce),
    .mem_data_cmd_v_o(mem_data_cmd_v_from_cce),
    .mem_data_cmd_ready_i(mem_data_cmd_ready_to_cce),
    .cce_id_i(cce_id_i[0]),
    .boot_rom_addr_o(boot_rom_addr_o),
    .boot_rom_data_i(boot_rom_data_i)
  );


endmodule



module bp_me_top_num_lce_p2_num_cce_p1_paddr_width_p22_lce_assoc_p8_lce_sets_p64_block_size_in_bytes_p64_num_inst_ram_els_p256
(
  clk_i,
  reset_i,
  lce_req_i,
  lce_req_v_i,
  lce_req_ready_o,
  lce_resp_i,
  lce_resp_v_i,
  lce_resp_ready_o,
  lce_data_resp_i,
  lce_data_resp_v_i,
  lce_data_resp_ready_o,
  lce_cmd_o,
  lce_cmd_v_o,
  lce_cmd_ready_i,
  lce_data_cmd_o,
  lce_data_cmd_v_o,
  lce_data_cmd_ready_i,
  lce_data_cmd_i,
  lce_data_cmd_v_i,
  lce_data_cmd_ready_o,
  cce_inst_boot_rom_addr_o,
  cce_inst_boot_rom_data_i,
  mem_resp_i,
  mem_resp_v_i,
  mem_resp_ready_o,
  mem_data_resp_i,
  mem_data_resp_v_i,
  mem_data_resp_ready_o,
  mem_cmd_o,
  mem_cmd_v_o,
  mem_cmd_yumi_i,
  mem_data_cmd_o,
  mem_data_cmd_v_o,
  mem_data_cmd_yumi_i
);

  input [193:0] lce_req_i;
  input [1:0] lce_req_v_i;
  output [1:0] lce_req_ready_o;
  input [51:0] lce_resp_i;
  input [1:0] lce_resp_v_i;
  output [1:0] lce_resp_ready_o;
  input [1073:0] lce_data_resp_i;
  input [1:0] lce_data_resp_v_i;
  output [1:0] lce_data_resp_ready_o;
  output [71:0] lce_cmd_o;
  output [1:0] lce_cmd_v_o;
  input [1:0] lce_cmd_ready_i;
  output [1035:0] lce_data_cmd_o;
  output [1:0] lce_data_cmd_v_o;
  input [1:0] lce_data_cmd_ready_i;
  input [1035:0] lce_data_cmd_i;
  input [1:0] lce_data_cmd_v_i;
  output [1:0] lce_data_cmd_ready_o;
  output [7:0] cce_inst_boot_rom_addr_o;
  input [95:0] cce_inst_boot_rom_data_i;
  input [57:0] mem_resp_i;
  input [0:0] mem_resp_v_i;
  output [0:0] mem_resp_ready_o;
  input [541:0] mem_data_resp_i;
  input [0:0] mem_data_resp_v_i;
  output [0:0] mem_data_resp_ready_o;
  output [29:0] mem_cmd_o;
  output [0:0] mem_cmd_v_o;
  input [0:0] mem_cmd_yumi_i;
  output [569:0] mem_data_cmd_o;
  output [0:0] mem_data_cmd_v_o;
  input [0:0] mem_data_cmd_yumi_i;
  input clk_i;
  input reset_i;
  wire [1:0] lce_req_ready_o,lce_resp_ready_o,lce_data_resp_ready_o,lce_cmd_v_o,
  lce_data_cmd_v_o,lce_data_cmd_ready_o;
  wire [71:0] lce_cmd_o;
  wire [1035:0] lce_data_cmd_o;
  wire [7:0] cce_inst_boot_rom_addr_o;
  wire [0:0] mem_resp_ready_o,mem_data_resp_ready_o,mem_cmd_v_o,mem_data_cmd_v_o,
  lce_cmd_v_o_from_cce,lce_cmd_ready_i_to_cce,lce_data_cmd_v_o_from_cce,
  lce_data_cmd_ready_i_to_cce,lce_req_v_i_to_cce,lce_req_ready_o_from_cce,lce_resp_v_i_to_cce,
  lce_resp_ready_o_from_cce,lce_data_resp_v_i_to_cce,lce_data_resp_ready_o_from_cce;
  wire [29:0] mem_cmd_o;
  wire [569:0] mem_data_cmd_o;
  wire [35:0] lce_cmd_o_from_cce;
  wire [517:0] lce_data_cmd_o_from_cce;
  wire [96:0] lce_req_i_to_cce;
  wire [25:0] lce_resp_i_to_cce;
  wire [536:0] lce_data_resp_i_to_cce;

  bp_me_network_num_lce_p2_num_cce_p1_paddr_width_p22_lce_assoc_p8_block_size_in_bytes_p64_data_width_p64
  network
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .lce_cmd_o(lce_cmd_o),
    .lce_cmd_v_o(lce_cmd_v_o),
    .lce_cmd_ready_i(lce_cmd_ready_i),
    .lce_cmd_i(lce_cmd_o_from_cce),
    .lce_cmd_v_i(lce_cmd_v_o_from_cce[0]),
    .lce_cmd_ready_o(lce_cmd_ready_i_to_cce[0]),
    .lce_data_cmd_o(lce_data_cmd_o),
    .lce_data_cmd_v_o(lce_data_cmd_v_o),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_i),
    .cce_lce_data_cmd_i(lce_data_cmd_o_from_cce),
    .cce_lce_data_cmd_v_i(lce_data_cmd_v_o_from_cce[0]),
    .cce_lce_data_cmd_ready_o(lce_data_cmd_ready_i_to_cce[0]),
    .lce_lce_data_cmd_i(lce_data_cmd_i),
    .lce_lce_data_cmd_v_i(lce_data_cmd_v_i),
    .lce_lce_data_cmd_ready_o(lce_data_cmd_ready_o),
    .lce_req_i(lce_req_i),
    .lce_req_v_i(lce_req_v_i),
    .lce_req_ready_o(lce_req_ready_o),
    .lce_req_o(lce_req_i_to_cce),
    .lce_req_v_o(lce_req_v_i_to_cce[0]),
    .lce_req_ready_i(lce_req_ready_o_from_cce[0]),
    .lce_resp_i(lce_resp_i),
    .lce_resp_v_i(lce_resp_v_i),
    .lce_resp_ready_o(lce_resp_ready_o),
    .lce_resp_o(lce_resp_i_to_cce),
    .lce_resp_v_o(lce_resp_v_i_to_cce[0]),
    .lce_resp_ready_i(lce_resp_ready_o_from_cce[0]),
    .lce_data_resp_i(lce_data_resp_i),
    .lce_data_resp_v_i(lce_data_resp_v_i),
    .lce_data_resp_ready_o(lce_data_resp_ready_o),
    .lce_data_resp_o(lce_data_resp_i_to_cce),
    .lce_data_resp_v_o(lce_data_resp_v_i_to_cce[0]),
    .lce_data_resp_ready_i(lce_data_resp_ready_o_from_cce[0])
  );


  bp_cce_top_num_lce_p2_num_cce_p1_paddr_width_p22_lce_assoc_p8_lce_sets_p64_block_size_in_bytes_p64_num_cce_inst_ram_els_p256_lce_req_data_width_p64
  genblk1_0__bp_cce_top
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .lce_req_i(lce_req_i_to_cce),
    .lce_req_v_i(lce_req_v_i_to_cce[0]),
    .lce_req_ready_o(lce_req_ready_o_from_cce[0]),
    .lce_resp_i(lce_resp_i_to_cce),
    .lce_resp_v_i(lce_resp_v_i_to_cce[0]),
    .lce_resp_ready_o(lce_resp_ready_o_from_cce[0]),
    .lce_data_resp_i(lce_data_resp_i_to_cce),
    .lce_data_resp_v_i(lce_data_resp_v_i_to_cce[0]),
    .lce_data_resp_ready_o(lce_data_resp_ready_o_from_cce[0]),
    .lce_cmd_o(lce_cmd_o_from_cce),
    .lce_cmd_v_o(lce_cmd_v_o_from_cce[0]),
    .lce_cmd_ready_i(lce_cmd_ready_i_to_cce[0]),
    .lce_data_cmd_o(lce_data_cmd_o_from_cce),
    .lce_data_cmd_v_o(lce_data_cmd_v_o_from_cce[0]),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_i_to_cce[0]),
    .mem_resp_i(mem_resp_i),
    .mem_resp_v_i(mem_resp_v_i[0]),
    .mem_resp_ready_o(mem_resp_ready_o[0]),
    .mem_data_resp_i(mem_data_resp_i),
    .mem_data_resp_v_i(mem_data_resp_v_i[0]),
    .mem_data_resp_ready_o(mem_data_resp_ready_o[0]),
    .mem_cmd_o(mem_cmd_o),
    .mem_cmd_v_o(mem_cmd_v_o[0]),
    .mem_cmd_yumi_i(mem_cmd_yumi_i[0]),
    .mem_data_cmd_o(mem_data_cmd_o),
    .mem_data_cmd_v_o(mem_data_cmd_v_o[0]),
    .mem_data_cmd_yumi_i(mem_data_cmd_yumi_i[0]),
    .cce_id_i(1'b0),
    .boot_rom_addr_o(cce_inst_boot_rom_addr_o),
    .boot_rom_data_i(cce_inst_boot_rom_data_i)
  );


endmodule



module bp_multi_top
(
  clk_i,
  reset_i,
  cce_inst_boot_rom_addr_o,
  cce_inst_boot_rom_data_i,
  mem_resp_i,
  mem_resp_v_i,
  mem_resp_ready_o,
  mem_data_resp_i,
  mem_data_resp_v_i,
  mem_data_resp_ready_o,
  mem_cmd_o,
  mem_cmd_v_o,
  mem_cmd_yumi_i,
  mem_data_cmd_o,
  mem_data_cmd_v_o,
  mem_data_cmd_yumi_i,
  cmt_rd_w_v_o,
  cmt_rd_addr_o,
  cmt_mem_w_v_o,
  cmt_mem_addr_o,
  cmt_mem_op_o,
  cmt_data_o
);

  output [7:0] cce_inst_boot_rom_addr_o;
  input [95:0] cce_inst_boot_rom_data_i;
  input [57:0] mem_resp_i;
  input [0:0] mem_resp_v_i;
  output [0:0] mem_resp_ready_o;
  input [541:0] mem_data_resp_i;
  input [0:0] mem_data_resp_v_i;
  output [0:0] mem_data_resp_ready_o;
  output [29:0] mem_cmd_o;
  output [0:0] mem_cmd_v_o;
  input [0:0] mem_cmd_yumi_i;
  output [569:0] mem_data_cmd_o;
  output [0:0] mem_data_cmd_v_o;
  input [0:0] mem_data_cmd_yumi_i;
  output [0:0] cmt_rd_w_v_o;
  output [4:0] cmt_rd_addr_o;
  output [0:0] cmt_mem_w_v_o;
  output [63:0] cmt_mem_addr_o;
  output [3:0] cmt_mem_op_o;
  output [63:0] cmt_data_o;
  input clk_i;
  input reset_i;
  wire [7:0] cce_inst_boot_rom_addr_o;
  wire [0:0] mem_resp_ready_o,mem_data_resp_ready_o,mem_cmd_v_o,mem_data_cmd_v_o,
  cmt_rd_w_v_o,cmt_mem_w_v_o;
  wire [29:0] mem_cmd_o;
  wire [569:0] mem_data_cmd_o;
  wire [4:0] cmt_rd_addr_o;
  wire [63:0] cmt_mem_addr_o,cmt_data_o;
  wire [3:0] cmt_mem_op_o;
  wire [193:0] lce_req;
  wire [1:0] lce_req_v,lce_req_ready,lce_resp_v,lce_resp_ready,lce_data_resp_v,
  lce_data_resp_ready,lce_cmd_v,lce_cmd_ready,lce_data_cmd_v_li,lce_data_cmd_ready_lo,
  lce_data_cmd_v_lo,lce_data_cmd_ready_li;
  wire [51:0] lce_resp;
  wire [1073:0] lce_data_resp;
  wire [71:0] lce_cmd;
  wire [1035:0] lce_data_cmd_li,lce_data_cmd_lo;

  bp_core_core_els_p1_num_lce_p2_num_cce_p1_lce_assoc_p8_lce_sets_p64_cce_block_size_in_bytes_p64_data_width_p64_vaddr_width_p39_paddr_width_p22_branch_metadata_fwd_width_p36_asid_width_p10_btb_indx_width_p9_bht_indx_width_p5_ras_addr_width_p22_trace_p0
  rof1_0__core
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .proc_cfg_i({ 1'b0, 1'b0, 1'b1 }),
    .lce_req_o(lce_req),
    .lce_req_v_o(lce_req_v),
    .lce_req_ready_i(lce_req_ready),
    .lce_resp_o(lce_resp),
    .lce_resp_v_o(lce_resp_v),
    .lce_resp_ready_i(lce_resp_ready),
    .lce_data_resp_o(lce_data_resp),
    .lce_data_resp_v_o(lce_data_resp_v),
    .lce_data_resp_ready_i(lce_data_resp_ready),
    .lce_cmd_i(lce_cmd),
    .lce_cmd_v_i(lce_cmd_v),
    .lce_cmd_ready_o(lce_cmd_ready),
    .lce_data_cmd_i(lce_data_cmd_li),
    .lce_data_cmd_v_i(lce_data_cmd_v_li),
    .lce_data_cmd_ready_o(lce_data_cmd_ready_lo),
    .lce_data_cmd_o(lce_data_cmd_lo),
    .lce_data_cmd_v_o(lce_data_cmd_v_lo),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_li),
    .cmt_rd_w_v_o(cmt_rd_w_v_o[0]),
    .cmt_rd_addr_o(cmt_rd_addr_o),
    .cmt_mem_w_v_o(cmt_mem_w_v_o[0]),
    .cmt_mem_addr_o(cmt_mem_addr_o),
    .cmt_mem_op_o(cmt_mem_op_o),
    .cmt_data_o(cmt_data_o)
  );


  bp_me_top_num_lce_p2_num_cce_p1_paddr_width_p22_lce_assoc_p8_lce_sets_p64_block_size_in_bytes_p64_num_inst_ram_els_p256
  me
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .lce_req_i(lce_req),
    .lce_req_v_i(lce_req_v),
    .lce_req_ready_o(lce_req_ready),
    .lce_resp_i(lce_resp),
    .lce_resp_v_i(lce_resp_v),
    .lce_resp_ready_o(lce_resp_ready),
    .lce_data_resp_i(lce_data_resp),
    .lce_data_resp_v_i(lce_data_resp_v),
    .lce_data_resp_ready_o(lce_data_resp_ready),
    .lce_cmd_o(lce_cmd),
    .lce_cmd_v_o(lce_cmd_v),
    .lce_cmd_ready_i(lce_cmd_ready),
    .lce_data_cmd_o(lce_data_cmd_li),
    .lce_data_cmd_v_o(lce_data_cmd_v_li),
    .lce_data_cmd_ready_i(lce_data_cmd_ready_lo),
    .lce_data_cmd_i(lce_data_cmd_lo),
    .lce_data_cmd_v_i(lce_data_cmd_v_lo),
    .lce_data_cmd_ready_o(lce_data_cmd_ready_li),
    .cce_inst_boot_rom_addr_o(cce_inst_boot_rom_addr_o),
    .cce_inst_boot_rom_data_i(cce_inst_boot_rom_data_i),
    .mem_resp_i(mem_resp_i),
    .mem_resp_v_i(mem_resp_v_i[0]),
    .mem_resp_ready_o(mem_resp_ready_o[0]),
    .mem_data_resp_i(mem_data_resp_i),
    .mem_data_resp_v_i(mem_data_resp_v_i[0]),
    .mem_data_resp_ready_o(mem_data_resp_ready_o[0]),
    .mem_cmd_o(mem_cmd_o),
    .mem_cmd_v_o(mem_cmd_v_o[0]),
    .mem_cmd_yumi_i(mem_cmd_yumi_i[0]),
    .mem_data_cmd_o(mem_data_cmd_o),
    .mem_data_cmd_v_o(mem_data_cmd_v_o[0]),
    .mem_data_cmd_yumi_i(mem_data_cmd_yumi_i[0])
  );


endmodule

