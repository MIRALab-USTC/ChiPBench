VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MACRO macro_9x6
  FOREIGN macro_9x6 0 0 ;
  CLASS BLOCK ;
  SIZE 98.385 BY 146.575 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 144.115 97.28 144.285 ;
        RECT  1.14 141.315 97.28 141.485 ;
        RECT  1.14 138.515 97.28 138.685 ;
        RECT  1.14 135.715 97.28 135.885 ;
        RECT  1.14 132.915 97.28 133.085 ;
        RECT  1.14 130.115 97.28 130.285 ;
        RECT  1.14 127.315 97.28 127.485 ;
        RECT  1.14 124.515 97.28 124.685 ;
        RECT  1.14 121.715 97.28 121.885 ;
        RECT  1.14 118.915 97.28 119.085 ;
        RECT  1.14 116.115 97.28 116.285 ;
        RECT  1.14 113.315 97.28 113.485 ;
        RECT  1.14 110.515 97.28 110.685 ;
        RECT  1.14 107.715 97.28 107.885 ;
        RECT  1.14 104.915 97.28 105.085 ;
        RECT  1.14 102.115 97.28 102.285 ;
        RECT  1.14 99.315 97.28 99.485 ;
        RECT  1.14 96.515 97.28 96.685 ;
        RECT  1.14 93.715 97.28 93.885 ;
        RECT  1.14 90.915 97.28 91.085 ;
        RECT  1.14 88.115 97.28 88.285 ;
        RECT  1.14 85.315 97.28 85.485 ;
        RECT  1.14 82.515 97.28 82.685 ;
        RECT  1.14 79.715 97.28 79.885 ;
        RECT  1.14 76.915 97.28 77.085 ;
        RECT  1.14 74.115 97.28 74.285 ;
        RECT  1.14 71.315 97.28 71.485 ;
        RECT  1.14 68.515 97.28 68.685 ;
        RECT  1.14 65.715 97.28 65.885 ;
        RECT  1.14 62.915 97.28 63.085 ;
        RECT  1.14 60.115 97.28 60.285 ;
        RECT  1.14 57.315 97.28 57.485 ;
        RECT  1.14 54.515 97.28 54.685 ;
        RECT  1.14 51.715 97.28 51.885 ;
        RECT  1.14 48.915 97.28 49.085 ;
        RECT  1.14 46.115 97.28 46.285 ;
        RECT  1.14 43.315 97.28 43.485 ;
        RECT  1.14 40.515 97.28 40.685 ;
        RECT  1.14 37.715 97.28 37.885 ;
        RECT  1.14 34.915 97.28 35.085 ;
        RECT  1.14 32.115 97.28 32.285 ;
        RECT  1.14 29.315 97.28 29.485 ;
        RECT  1.14 26.515 97.28 26.685 ;
        RECT  1.14 23.715 97.28 23.885 ;
        RECT  1.14 20.915 97.28 21.085 ;
        RECT  1.14 18.115 97.28 18.285 ;
        RECT  1.14 15.315 97.28 15.485 ;
        RECT  1.14 12.515 97.28 12.685 ;
        RECT  1.14 9.715 97.28 9.885 ;
        RECT  1.14 6.915 97.28 7.085 ;
        RECT  1.14 4.115 97.28 4.285 ;
        RECT  1.14 1.315 97.28 1.485 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 142.715 97.28 142.885 ;
        RECT  1.14 139.915 97.28 140.085 ;
        RECT  1.14 137.115 97.28 137.285 ;
        RECT  1.14 134.315 97.28 134.485 ;
        RECT  1.14 131.515 97.28 131.685 ;
        RECT  1.14 128.715 97.28 128.885 ;
        RECT  1.14 125.915 97.28 126.085 ;
        RECT  1.14 123.115 97.28 123.285 ;
        RECT  1.14 120.315 97.28 120.485 ;
        RECT  1.14 117.515 97.28 117.685 ;
        RECT  1.14 114.715 97.28 114.885 ;
        RECT  1.14 111.915 97.28 112.085 ;
        RECT  1.14 109.115 97.28 109.285 ;
        RECT  1.14 106.315 97.28 106.485 ;
        RECT  1.14 103.515 97.28 103.685 ;
        RECT  1.14 100.715 97.28 100.885 ;
        RECT  1.14 97.915 97.28 98.085 ;
        RECT  1.14 95.115 97.28 95.285 ;
        RECT  1.14 92.315 97.28 92.485 ;
        RECT  1.14 89.515 97.28 89.685 ;
        RECT  1.14 86.715 97.28 86.885 ;
        RECT  1.14 83.915 97.28 84.085 ;
        RECT  1.14 81.115 97.28 81.285 ;
        RECT  1.14 78.315 97.28 78.485 ;
        RECT  1.14 75.515 97.28 75.685 ;
        RECT  1.14 72.715 97.28 72.885 ;
        RECT  1.14 69.915 97.28 70.085 ;
        RECT  1.14 67.115 97.28 67.285 ;
        RECT  1.14 64.315 97.28 64.485 ;
        RECT  1.14 61.515 97.28 61.685 ;
        RECT  1.14 58.715 97.28 58.885 ;
        RECT  1.14 55.915 97.28 56.085 ;
        RECT  1.14 53.115 97.28 53.285 ;
        RECT  1.14 50.315 97.28 50.485 ;
        RECT  1.14 47.515 97.28 47.685 ;
        RECT  1.14 44.715 97.28 44.885 ;
        RECT  1.14 41.915 97.28 42.085 ;
        RECT  1.14 39.115 97.28 39.285 ;
        RECT  1.14 36.315 97.28 36.485 ;
        RECT  1.14 33.515 97.28 33.685 ;
        RECT  1.14 30.715 97.28 30.885 ;
        RECT  1.14 27.915 97.28 28.085 ;
        RECT  1.14 25.115 97.28 25.285 ;
        RECT  1.14 22.315 97.28 22.485 ;
        RECT  1.14 19.515 97.28 19.685 ;
        RECT  1.14 16.715 97.28 16.885 ;
        RECT  1.14 13.915 97.28 14.085 ;
        RECT  1.14 11.115 97.28 11.285 ;
        RECT  1.14 8.315 97.28 8.485 ;
        RECT  1.14 5.515 97.28 5.685 ;
        RECT  1.14 2.715 97.28 2.885 ;
    END
  END VDD
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  65.545 146.435 65.685 146.575 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 33.075 0.07 33.145 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 129.955 0.07 130.025 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  98.315 129.675 98.385 129.745 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  98.315 97.475 98.385 97.545 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  98.315 64.995 98.385 65.065 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  97.465 146.435 97.605 146.575 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  98.315 16.555 98.385 16.625 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 49.035 0.07 49.105 ;
    END
  END addr[8]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 16.835 0.07 16.905 ;
    END
  END clk
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  98.315 32.795 98.385 32.865 ;
    END
  END cs
  PIN di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END di[0]
  PIN di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  32.505 0 32.645 0.14 ;
    END
  END di[1]
  PIN di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 146.435 0.725 146.575 ;
    END
  END di[2]
  PIN di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  98.315 49.035 98.385 49.105 ;
    END
  END di[3]
  PIN di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  64.985 0 65.125 0.14 ;
    END
  END di[4]
  PIN di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 113.715 0.07 113.785 ;
    END
  END di[5]
  PIN doq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  98.315 113.435 98.385 113.505 ;
    END
  END doq[0]
  PIN doq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 81.515 0.07 81.585 ;
    END
  END doq[1]
  PIN doq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  33.065 146.435 33.205 146.575 ;
    END
  END doq[2]
  PIN doq[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  97.465 0 97.605 0.14 ;
    END
  END doq[3]
  PIN doq[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 65.275 0.07 65.345 ;
    END
  END doq[4]
  PIN doq[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 97.475 0.07 97.545 ;
    END
  END doq[5]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  98.315 81.235 98.385 81.305 ;
    END
  END we
  OBS
    LAYER metal1 ;
     RECT  0 -0.085 3.23 146.575 ;
     RECT  3.23 0 98.385 146.575 ;
    LAYER metal2 ;
     RECT  0 0 98.385 146.575 ;
    LAYER metal3 ;
     RECT  0 0 98.385 146.575 ;
    LAYER metal4 ;
     RECT  0 0 98.385 146.575 ;
  END
END macro_9x6
END LIBRARY
