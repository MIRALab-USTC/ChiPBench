VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MACRO macro_11x2
  FOREIGN macro_11x2 0 0 ;
  CLASS BLOCK ;
  SIZE 81.285 BY 239.85 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 236.515 80.18 236.685 ;
        RECT  1.14 233.715 80.18 233.885 ;
        RECT  1.14 230.915 80.18 231.085 ;
        RECT  1.14 228.115 80.18 228.285 ;
        RECT  1.14 225.315 80.18 225.485 ;
        RECT  1.14 222.515 80.18 222.685 ;
        RECT  1.14 219.715 80.18 219.885 ;
        RECT  1.14 216.915 80.18 217.085 ;
        RECT  1.14 214.115 80.18 214.285 ;
        RECT  1.14 211.315 80.18 211.485 ;
        RECT  1.14 208.515 80.18 208.685 ;
        RECT  1.14 205.715 80.18 205.885 ;
        RECT  1.14 202.915 80.18 203.085 ;
        RECT  1.14 200.115 80.18 200.285 ;
        RECT  1.14 197.315 80.18 197.485 ;
        RECT  1.14 194.515 80.18 194.685 ;
        RECT  1.14 191.715 80.18 191.885 ;
        RECT  1.14 188.915 80.18 189.085 ;
        RECT  1.14 186.115 80.18 186.285 ;
        RECT  1.14 183.315 80.18 183.485 ;
        RECT  1.14 180.515 80.18 180.685 ;
        RECT  1.14 177.715 80.18 177.885 ;
        RECT  1.14 174.915 80.18 175.085 ;
        RECT  1.14 172.115 80.18 172.285 ;
        RECT  1.14 169.315 80.18 169.485 ;
        RECT  1.14 166.515 80.18 166.685 ;
        RECT  1.14 163.715 80.18 163.885 ;
        RECT  1.14 160.915 80.18 161.085 ;
        RECT  1.14 158.115 80.18 158.285 ;
        RECT  1.14 155.315 80.18 155.485 ;
        RECT  1.14 152.515 80.18 152.685 ;
        RECT  1.14 149.715 80.18 149.885 ;
        RECT  1.14 146.915 80.18 147.085 ;
        RECT  1.14 144.115 80.18 144.285 ;
        RECT  1.14 141.315 80.18 141.485 ;
        RECT  1.14 138.515 80.18 138.685 ;
        RECT  1.14 135.715 80.18 135.885 ;
        RECT  1.14 132.915 80.18 133.085 ;
        RECT  1.14 130.115 80.18 130.285 ;
        RECT  1.14 127.315 80.18 127.485 ;
        RECT  1.14 124.515 80.18 124.685 ;
        RECT  1.14 121.715 80.18 121.885 ;
        RECT  1.14 118.915 80.18 119.085 ;
        RECT  1.14 116.115 80.18 116.285 ;
        RECT  1.14 113.315 80.18 113.485 ;
        RECT  1.14 110.515 80.18 110.685 ;
        RECT  1.14 107.715 80.18 107.885 ;
        RECT  1.14 104.915 80.18 105.085 ;
        RECT  1.14 102.115 80.18 102.285 ;
        RECT  1.14 99.315 80.18 99.485 ;
        RECT  1.14 96.515 80.18 96.685 ;
        RECT  1.14 93.715 80.18 93.885 ;
        RECT  1.14 90.915 80.18 91.085 ;
        RECT  1.14 88.115 80.18 88.285 ;
        RECT  1.14 85.315 80.18 85.485 ;
        RECT  1.14 82.515 80.18 82.685 ;
        RECT  1.14 79.715 80.18 79.885 ;
        RECT  1.14 76.915 80.18 77.085 ;
        RECT  1.14 74.115 80.18 74.285 ;
        RECT  1.14 71.315 80.18 71.485 ;
        RECT  1.14 68.515 80.18 68.685 ;
        RECT  1.14 65.715 80.18 65.885 ;
        RECT  1.14 62.915 80.18 63.085 ;
        RECT  1.14 60.115 80.18 60.285 ;
        RECT  1.14 57.315 80.18 57.485 ;
        RECT  1.14 54.515 80.18 54.685 ;
        RECT  1.14 51.715 80.18 51.885 ;
        RECT  1.14 48.915 80.18 49.085 ;
        RECT  1.14 46.115 80.18 46.285 ;
        RECT  1.14 43.315 80.18 43.485 ;
        RECT  1.14 40.515 80.18 40.685 ;
        RECT  1.14 37.715 80.18 37.885 ;
        RECT  1.14 34.915 80.18 35.085 ;
        RECT  1.14 32.115 80.18 32.285 ;
        RECT  1.14 29.315 80.18 29.485 ;
        RECT  1.14 26.515 80.18 26.685 ;
        RECT  1.14 23.715 80.18 23.885 ;
        RECT  1.14 20.915 80.18 21.085 ;
        RECT  1.14 18.115 80.18 18.285 ;
        RECT  1.14 15.315 80.18 15.485 ;
        RECT  1.14 12.515 80.18 12.685 ;
        RECT  1.14 9.715 80.18 9.885 ;
        RECT  1.14 6.915 80.18 7.085 ;
        RECT  1.14 4.115 80.18 4.285 ;
        RECT  1.14 1.315 80.18 1.485 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 237.915 80.18 238.085 ;
        RECT  1.14 235.115 80.18 235.285 ;
        RECT  1.14 232.315 80.18 232.485 ;
        RECT  1.14 229.515 80.18 229.685 ;
        RECT  1.14 226.715 80.18 226.885 ;
        RECT  1.14 223.915 80.18 224.085 ;
        RECT  1.14 221.115 80.18 221.285 ;
        RECT  1.14 218.315 80.18 218.485 ;
        RECT  1.14 215.515 80.18 215.685 ;
        RECT  1.14 212.715 80.18 212.885 ;
        RECT  1.14 209.915 80.18 210.085 ;
        RECT  1.14 207.115 80.18 207.285 ;
        RECT  1.14 204.315 80.18 204.485 ;
        RECT  1.14 201.515 80.18 201.685 ;
        RECT  1.14 198.715 80.18 198.885 ;
        RECT  1.14 195.915 80.18 196.085 ;
        RECT  1.14 193.115 80.18 193.285 ;
        RECT  1.14 190.315 80.18 190.485 ;
        RECT  1.14 187.515 80.18 187.685 ;
        RECT  1.14 184.715 80.18 184.885 ;
        RECT  1.14 181.915 80.18 182.085 ;
        RECT  1.14 179.115 80.18 179.285 ;
        RECT  1.14 176.315 80.18 176.485 ;
        RECT  1.14 173.515 80.18 173.685 ;
        RECT  1.14 170.715 80.18 170.885 ;
        RECT  1.14 167.915 80.18 168.085 ;
        RECT  1.14 165.115 80.18 165.285 ;
        RECT  1.14 162.315 80.18 162.485 ;
        RECT  1.14 159.515 80.18 159.685 ;
        RECT  1.14 156.715 80.18 156.885 ;
        RECT  1.14 153.915 80.18 154.085 ;
        RECT  1.14 151.115 80.18 151.285 ;
        RECT  1.14 148.315 80.18 148.485 ;
        RECT  1.14 145.515 80.18 145.685 ;
        RECT  1.14 142.715 80.18 142.885 ;
        RECT  1.14 139.915 80.18 140.085 ;
        RECT  1.14 137.115 80.18 137.285 ;
        RECT  1.14 134.315 80.18 134.485 ;
        RECT  1.14 131.515 80.18 131.685 ;
        RECT  1.14 128.715 80.18 128.885 ;
        RECT  1.14 125.915 80.18 126.085 ;
        RECT  1.14 123.115 80.18 123.285 ;
        RECT  1.14 120.315 80.18 120.485 ;
        RECT  1.14 117.515 80.18 117.685 ;
        RECT  1.14 114.715 80.18 114.885 ;
        RECT  1.14 111.915 80.18 112.085 ;
        RECT  1.14 109.115 80.18 109.285 ;
        RECT  1.14 106.315 80.18 106.485 ;
        RECT  1.14 103.515 80.18 103.685 ;
        RECT  1.14 100.715 80.18 100.885 ;
        RECT  1.14 97.915 80.18 98.085 ;
        RECT  1.14 95.115 80.18 95.285 ;
        RECT  1.14 92.315 80.18 92.485 ;
        RECT  1.14 89.515 80.18 89.685 ;
        RECT  1.14 86.715 80.18 86.885 ;
        RECT  1.14 83.915 80.18 84.085 ;
        RECT  1.14 81.115 80.18 81.285 ;
        RECT  1.14 78.315 80.18 78.485 ;
        RECT  1.14 75.515 80.18 75.685 ;
        RECT  1.14 72.715 80.18 72.885 ;
        RECT  1.14 69.915 80.18 70.085 ;
        RECT  1.14 67.115 80.18 67.285 ;
        RECT  1.14 64.315 80.18 64.485 ;
        RECT  1.14 61.515 80.18 61.685 ;
        RECT  1.14 58.715 80.18 58.885 ;
        RECT  1.14 55.915 80.18 56.085 ;
        RECT  1.14 53.115 80.18 53.285 ;
        RECT  1.14 50.315 80.18 50.485 ;
        RECT  1.14 47.515 80.18 47.685 ;
        RECT  1.14 44.715 80.18 44.885 ;
        RECT  1.14 41.915 80.18 42.085 ;
        RECT  1.14 39.115 80.18 39.285 ;
        RECT  1.14 36.315 80.18 36.485 ;
        RECT  1.14 33.515 80.18 33.685 ;
        RECT  1.14 30.715 80.18 30.885 ;
        RECT  1.14 27.915 80.18 28.085 ;
        RECT  1.14 25.115 80.18 25.285 ;
        RECT  1.14 22.315 80.18 22.485 ;
        RECT  1.14 19.515 80.18 19.685 ;
        RECT  1.14 16.715 80.18 16.885 ;
        RECT  1.14 13.915 80.18 14.085 ;
        RECT  1.14 11.115 80.18 11.285 ;
        RECT  1.14 8.315 80.18 8.485 ;
        RECT  1.14 5.515 80.18 5.685 ;
        RECT  1.14 2.715 80.18 2.885 ;
    END
  END VDD
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  81.215 115.395 81.285 115.465 ;
    END
  END addr[0]
  PIN addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  81.215 208.075 81.285 208.145 ;
    END
  END addr[10]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 217.315 0.07 217.385 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  81.215 53.515 81.285 53.585 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 124.355 0.07 124.425 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 186.235 0.07 186.305 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  80.105 239.71 80.245 239.85 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  81.215 84.315 81.285 84.385 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  62.185 0 62.325 0.14 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.675 0.07 31.745 ;
    END
  END addr[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  81.215 177.275 81.285 177.345 ;
    END
  END clk
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 62.475 0.07 62.545 ;
    END
  END cs
  PIN di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  18.505 239.71 18.645 239.85 ;
    END
  END di[0]
  PIN di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  81.215 22.435 81.285 22.505 ;
    END
  END di[1]
  PIN doq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 93.555 0.07 93.625 ;
    END
  END doq[0]
  PIN doq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 155.435 0.07 155.505 ;
    END
  END doq[1]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  81.215 146.195 81.285 146.265 ;
    END
  END we
  OBS
    LAYER metal1 ;
     RECT  0 -0.085 3.23 239.85 ;
     RECT  3.23 0 81.285 239.85 ;
    LAYER metal2 ;
     RECT  0 0 81.285 239.85 ;
    LAYER metal3 ;
     RECT  0 0 81.285 239.85 ;
    LAYER metal4 ;
     RECT  0 0 81.285 239.85 ;
  END
END macro_11x2
END LIBRARY
