VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MACRO memMod_dist_1
  FOREIGN memMod_dist_1 0 0 ;
  CLASS BLOCK ;
  SIZE 54.285 BY 106.565 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 104.915 53.2 105.085 ;
        RECT  1.14 102.115 53.2 102.285 ;
        RECT  1.14 99.315 53.2 99.485 ;
        RECT  1.14 96.515 53.2 96.685 ;
        RECT  1.14 93.715 53.2 93.885 ;
        RECT  1.14 90.915 53.2 91.085 ;
        RECT  1.14 88.115 53.2 88.285 ;
        RECT  1.14 85.315 53.2 85.485 ;
        RECT  1.14 82.515 53.2 82.685 ;
        RECT  1.14 79.715 53.2 79.885 ;
        RECT  1.14 76.915 53.2 77.085 ;
        RECT  1.14 74.115 53.2 74.285 ;
        RECT  1.14 71.315 53.2 71.485 ;
        RECT  1.14 68.515 53.2 68.685 ;
        RECT  1.14 65.715 53.2 65.885 ;
        RECT  1.14 62.915 53.2 63.085 ;
        RECT  1.14 60.115 53.2 60.285 ;
        RECT  1.14 57.315 53.2 57.485 ;
        RECT  1.14 54.515 53.2 54.685 ;
        RECT  1.14 51.715 53.2 51.885 ;
        RECT  1.14 48.915 53.2 49.085 ;
        RECT  1.14 46.115 53.2 46.285 ;
        RECT  1.14 43.315 53.2 43.485 ;
        RECT  1.14 40.515 53.2 40.685 ;
        RECT  1.14 37.715 53.2 37.885 ;
        RECT  1.14 34.915 53.2 35.085 ;
        RECT  1.14 32.115 53.2 32.285 ;
        RECT  1.14 29.315 53.2 29.485 ;
        RECT  1.14 26.515 53.2 26.685 ;
        RECT  1.14 23.715 53.2 23.885 ;
        RECT  1.14 20.915 53.2 21.085 ;
        RECT  1.14 18.115 53.2 18.285 ;
        RECT  1.14 15.315 53.2 15.485 ;
        RECT  1.14 12.515 53.2 12.685 ;
        RECT  1.14 9.715 53.2 9.885 ;
        RECT  1.14 6.915 53.2 7.085 ;
        RECT  1.14 4.115 53.2 4.285 ;
        RECT  1.14 1.315 53.2 1.485 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 103.515 53.2 103.685 ;
        RECT  1.14 100.715 53.2 100.885 ;
        RECT  1.14 97.915 53.2 98.085 ;
        RECT  1.14 95.115 53.2 95.285 ;
        RECT  1.14 92.315 53.2 92.485 ;
        RECT  1.14 89.515 53.2 89.685 ;
        RECT  1.14 86.715 53.2 86.885 ;
        RECT  1.14 83.915 53.2 84.085 ;
        RECT  1.14 81.115 53.2 81.285 ;
        RECT  1.14 78.315 53.2 78.485 ;
        RECT  1.14 75.515 53.2 75.685 ;
        RECT  1.14 72.715 53.2 72.885 ;
        RECT  1.14 69.915 53.2 70.085 ;
        RECT  1.14 67.115 53.2 67.285 ;
        RECT  1.14 64.315 53.2 64.485 ;
        RECT  1.14 61.515 53.2 61.685 ;
        RECT  1.14 58.715 53.2 58.885 ;
        RECT  1.14 55.915 53.2 56.085 ;
        RECT  1.14 53.115 53.2 53.285 ;
        RECT  1.14 50.315 53.2 50.485 ;
        RECT  1.14 47.515 53.2 47.685 ;
        RECT  1.14 44.715 53.2 44.885 ;
        RECT  1.14 41.915 53.2 42.085 ;
        RECT  1.14 39.115 53.2 39.285 ;
        RECT  1.14 36.315 53.2 36.485 ;
        RECT  1.14 33.515 53.2 33.685 ;
        RECT  1.14 30.715 53.2 30.885 ;
        RECT  1.14 27.915 53.2 28.085 ;
        RECT  1.14 25.115 53.2 25.285 ;
        RECT  1.14 22.315 53.2 22.485 ;
        RECT  1.14 19.515 53.2 19.685 ;
        RECT  1.14 16.715 53.2 16.885 ;
        RECT  1.14 13.915 53.2 14.085 ;
        RECT  1.14 11.115 53.2 11.285 ;
        RECT  1.14 8.315 53.2 8.485 ;
        RECT  1.14 5.515 53.2 5.685 ;
        RECT  1.14 2.715 53.2 2.885 ;
    END
  END VDD
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 34.475 54.285 34.545 ;
    END
  END clk
  PIN inAddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 52.395 54.285 52.465 ;
    END
  END inAddr[0]
  PIN inAddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 80.955 54.285 81.025 ;
    END
  END inAddr[1]
  PIN inAddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 47.075 0.07 47.145 ;
    END
  END inAddr[2]
  PIN inAddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 25.515 0.07 25.585 ;
    END
  END inAddr[3]
  PIN in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  35.865 0 36.005 0.14 ;
    END
  END in[0]
  PIN in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.945 106.425 18.085 106.565 ;
    END
  END in[10]
  PIN in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  53.225 106.425 53.365 106.565 ;
    END
  END in[11]
  PIN in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 39.795 0.07 39.865 ;
    END
  END in[12]
  PIN in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 27.475 54.285 27.545 ;
    END
  END in[13]
  PIN in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 48.755 54.285 48.825 ;
    END
  END in[14]
  PIN in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 59.395 54.285 59.465 ;
    END
  END in[15]
  PIN in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 87.955 54.285 88.025 ;
    END
  END in[16]
  PIN in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 91.595 54.285 91.665 ;
    END
  END in[17]
  PIN in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 89.635 0.07 89.705 ;
    END
  END in[18]
  PIN in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 54.075 0.07 54.145 ;
    END
  END in[19]
  PIN in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  49.865 0 50.005 0.14 ;
    END
  END in[1]
  PIN in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.875 0.07 7.945 ;
    END
  END in[20]
  PIN in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 56.035 54.285 56.105 ;
    END
  END in[21]
  PIN in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 4.235 0.07 4.305 ;
    END
  END in[22]
  PIN in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 77.315 54.285 77.385 ;
    END
  END in[23]
  PIN in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 84.315 54.285 84.385 ;
    END
  END in[24]
  PIN in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 23.835 54.285 23.905 ;
    END
  END in[25]
  PIN in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 61.075 0.07 61.145 ;
    END
  END in[26]
  PIN in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 78.995 0.07 79.065 ;
    END
  END in[27]
  PIN in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 13.195 54.285 13.265 ;
    END
  END in[28]
  PIN in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 43.435 0.07 43.505 ;
    END
  END in[29]
  PIN in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 71.995 0.07 72.065 ;
    END
  END in[2]
  PIN in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 50.435 0.07 50.505 ;
    END
  END in[30]
  PIN in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.665 106.425 10.805 106.565 ;
    END
  END in[31]
  PIN in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 11.515 0.07 11.585 ;
    END
  END in[3]
  PIN in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  28.585 0 28.725 0.14 ;
    END
  END in[4]
  PIN in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 14.875 0.07 14.945 ;
    END
  END in[5]
  PIN in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 68.355 0.07 68.425 ;
    END
  END in[6]
  PIN in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 38.115 54.285 38.185 ;
    END
  END in[7]
  PIN in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 96.635 0.07 96.705 ;
    END
  END in[8]
  PIN in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  46.505 106.425 46.645 106.565 ;
    END
  END in[9]
  PIN outAddr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 31.115 54.285 31.185 ;
    END
  END outAddr[0]
  PIN outAddr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 100.275 0.07 100.345 ;
    END
  END outAddr[1]
  PIN outAddr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 45.395 54.285 45.465 ;
    END
  END outAddr[2]
  PIN outAddr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 63.035 54.285 63.105 ;
    END
  END outAddr[3]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 16.835 54.285 16.905 ;
    END
  END out[0]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 66.675 54.285 66.745 ;
    END
  END out[10]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 93.275 0.07 93.345 ;
    END
  END out[11]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  3.945 106.425 4.085 106.565 ;
    END
  END out[12]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 64.715 0.07 64.785 ;
    END
  END out[13]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END out[14]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 32.795 0.07 32.865 ;
    END
  END out[15]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 103.915 0.07 103.985 ;
    END
  END out[16]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  25.225 106.425 25.365 106.565 ;
    END
  END out[17]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 102.235 54.285 102.305 ;
    END
  END out[18]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 85.995 0.07 86.065 ;
    END
  END out[19]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.585 0 14.725 0.14 ;
    END
  END out[1]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.305 0 7.445 0.14 ;
    END
  END out[20]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 98.595 54.285 98.665 ;
    END
  END out[21]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 29.155 0.07 29.225 ;
    END
  END out[22]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 2.555 54.285 2.625 ;
    END
  END out[23]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 94.955 54.285 95.025 ;
    END
  END out[24]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 41.755 54.285 41.825 ;
    END
  END out[25]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 18.515 0.07 18.585 ;
    END
  END out[26]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 36.435 0.07 36.505 ;
    END
  END out[27]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  21.865 0 22.005 0.14 ;
    END
  END out[28]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  43.145 0 43.285 0.14 ;
    END
  END out[29]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 6.195 54.285 6.265 ;
    END
  END out[2]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 73.675 54.285 73.745 ;
    END
  END out[30]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 9.835 54.285 9.905 ;
    END
  END out[31]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  39.225 106.425 39.365 106.565 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.945 106.425 32.085 106.565 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 75.355 0.07 75.425 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 82.635 0.07 82.705 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 20.475 54.285 20.545 ;
    END
  END out[7]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 22.155 0.07 22.225 ;
    END
  END out[8]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 57.715 0.07 57.785 ;
    END
  END out[9]
  PIN writeSel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  54.215 70.035 54.285 70.105 ;
    END
  END writeSel
  OBS
    LAYER metal1 ;
     RECT  0 -0.085 3.23 106.565 ;
     RECT  3.23 0 54.285 106.565 ;
    LAYER metal2 ;
     RECT  0 0 54.285 106.565 ;
    LAYER metal3 ;
     RECT  0 0 54.285 106.565 ;
    LAYER metal4 ;
     RECT  0 0 54.285 106.565 ;
  END
END memMod_dist_1
END LIBRARY
