# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2010, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *     NGLibraryCreator, v2010.08-HR32-SP3-2010-08-05 - build 1009061800      *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on brazil06.nangate.com.br for user Giancarlo Franciscatto (gfr).
# Local time is now Fri, 3 Dec 2010, 19:32:18.
# Main process id is 27821.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.0050 ;

LAYER poly
  TYPE MASTERSLICE ;
END poly

LAYER active
  TYPE MASTERSLICE ;
END active

LAYER metal1
  TYPE ROUTING ;
  SPACING 0.065 ;
  WIDTH 0.07 ;
  PITCH 0.14 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.38 ;
  THICKNESS 0.13 ;
  HEIGHT 0.37 ;
  CAPACITANCE CPERSQDIST 7.7161e-05 ;
  EDGECAPACITANCE 2.7365e-05 ;
END metal1

LAYER via1
  TYPE CUT ;
  SPACING 0.08 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via1

LAYER metal2
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.3000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.0700     0.0700     0.0700     0.0700     0.0700     0.0700     
      WIDTH 0.0900       0.0700     0.0900     0.0900     0.0900     0.0900     0.0900     
      WIDTH 0.2700       0.0700     0.0900     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.0700     0.0900     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.0700     0.0900     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.0700     0.0900     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.07 ;
  PITCH 0.19 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.25 ;
  THICKNESS 0.14 ;
  HEIGHT 0.62 ;
  CAPACITANCE CPERSQDIST 4.0896e-05 ;
  EDGECAPACITANCE 2.5157e-05 ;
END metal2

LAYER via2
  TYPE CUT ;
  SPACING 0.09 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via2

LAYER metal3
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.3000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.0700     0.0700     0.0700     0.0700     0.0700     0.0700     
      WIDTH 0.0900       0.0700     0.0900     0.0900     0.0900     0.0900     0.0900     
      WIDTH 0.2700       0.0700     0.0900     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.0700     0.0900     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.0700     0.0900     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.0700     0.0900     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.07 ;
  PITCH 0.14 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.25 ;
  THICKNESS 0.14 ;
  HEIGHT 0.88 ;
  CAPACITANCE CPERSQDIST 2.7745e-05 ;
  EDGECAPACITANCE 2.5157e-05 ;
END metal3

LAYER via3
  TYPE CUT ;
  SPACING 0.09 ;
  WIDTH 0.07 ;
  RESISTANCE 5 ;
END via3

LAYER metal4
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.1400     0.1400     0.1400     0.1400     0.1400     
      WIDTH 0.2700       0.1400     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.1400     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.1400     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.1400     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.14 ;
  PITCH 0.28 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  HEIGHT 1.14 ;
  CAPACITANCE CPERSQDIST 2.0743e-05 ;
  EDGECAPACITANCE 3.0908e-05 ;
END metal4

LAYER via4
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  RESISTANCE 3 ;
END via4

LAYER metal5
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.1400     0.1400     0.1400     0.1400     0.1400     
      WIDTH 0.2700       0.1400     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.1400     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.1400     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.1400     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.14 ;
  PITCH 0.28 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  HEIGHT 1.71 ;
  CAPACITANCE CPERSQDIST 1.3527e-05 ;
  EDGECAPACITANCE 2.3863e-06 ;
END metal5

LAYER via5
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  RESISTANCE 3 ;
END via5

LAYER metal6
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     0.9000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.1400     0.1400     0.1400     0.1400     0.1400     
      WIDTH 0.2700       0.1400     0.2700     0.2700     0.2700     0.2700     
      WIDTH 0.5000       0.1400     0.2700     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.1400     0.2700     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.1400     0.2700     0.5000     0.9000     1.5000      ;
  WIDTH 0.14 ;
  PITCH 0.28 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.21 ;
  THICKNESS 0.28 ;
  HEIGHT 2.28 ;
  CAPACITANCE CPERSQDIST 1.0036e-05 ;
  EDGECAPACITANCE 2.3863e-05 ;
END metal6

LAYER via6
  TYPE CUT ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
  RESISTANCE 3 ;
END via6

LAYER metal7
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.4000     0.4000     0.4000     0.4000     
      WIDTH 0.5000       0.4000     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.4000     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.4000     0.5000     0.9000     1.5000      ;
  WIDTH 0.4 ;
  PITCH 0.8 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.075 ;
  THICKNESS 0.8 ;
  HEIGHT 2.85 ;
  CAPACITANCE CPERSQDIST 7.9771e-06 ;
  EDGECAPACITANCE 3.2577e-05 ;
END metal7

LAYER via7
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  RESISTANCE 1 ;
END via7

LAYER metal8
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     1.8000     2.7000     4.0000     
      WIDTH 0.0000       0.4000     0.4000     0.4000     0.4000     
      WIDTH 0.5000       0.4000     0.5000     0.5000     0.5000     
      WIDTH 0.9000       0.4000     0.5000     0.9000     0.9000     
      WIDTH 1.5000       0.4000     0.5000     0.9000     1.5000      ;
  WIDTH 0.4 ;
  PITCH 0.8 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.075 ;
  THICKNESS 0.8 ;
  HEIGHT 4.47 ;
  CAPACITANCE CPERSQDIST 5.0391e-06 ;
  EDGECAPACITANCE 2.3932e-05 ;
END metal8

LAYER via8
  TYPE CUT ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
  RESISTANCE 1 ;
END via8

LAYER metal9
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     2.7000     4.0000     
      WIDTH 0.0000       0.8000     0.8000     0.8000     
      WIDTH 0.9000       0.8000     0.9000     0.9000     
      WIDTH 1.5000       0.8000     0.9000     1.5000      ;
  WIDTH 0.8 ;
  PITCH 1.6 ;
  DIRECTION HORIZONTAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.03 ;
  THICKNESS 2 ;
  HEIGHT 6.09 ;
  CAPACITANCE CPERSQDIST 3.6827e-06 ;
  EDGECAPACITANCE 3.0803e-05 ;
END metal9

LAYER via9
  TYPE CUT ;
  SPACING 0.88 ;
  WIDTH 0.8 ;
  RESISTANCE 0.5 ;
END via9

LAYER metal10
  TYPE ROUTING ;
  SPACINGTABLE 
    PARALLELRUNLENGTH    0.0000     2.7000     4.0000     
      WIDTH 0.0000       0.8000     0.8000     0.8000     
      WIDTH 0.9000       0.8000     0.9000     0.9000     
      WIDTH 1.5000       0.8000     0.9000     1.5000      ;
  WIDTH 0.8 ;
  PITCH 1.6 ;
  DIRECTION VERTICAL ;
  OFFSET 0.095 0.07 ;
  RESISTANCE RPERSQ 0.03 ;
  THICKNESS 2 ;
  HEIGHT 10.09 ;
  CAPACITANCE CPERSQDIST 2.2124e-06 ;
  EDGECAPACITANCE 2.3667e-05 ;
END metal10

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA via1_4 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via1_4

VIA via1_0 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via1_0

VIA via1_1 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via1_1

VIA via1_2 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via1_2

VIA via1_3 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via1_3

VIA via1_5 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via1_5

VIA via1_6 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via1_6

VIA via1_7 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via1_7

VIA via1_8 DEFAULT
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal1 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via1_8

VIA via2_8 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via2_8

VIA via2_4 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via2_4

VIA via2_5 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via2_5

VIA via2_7 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via2_7

VIA via2_6 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2_6

VIA via2_0 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2_0

VIA via2_1 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
END via2_1

VIA via2_2 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
END via2_2

VIA via2_3 DEFAULT
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal2 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2_3

VIA via3_2 DEFAULT
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.035 0.07 0.035 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3_2

VIA via3_0 DEFAULT
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3_0

VIA via3_1 DEFAULT
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER metal3 ;
    RECT -0.035 -0.07 0.035 0.07 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3_1

VIA via4_0 DEFAULT
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via4_0

VIA via5_0 DEFAULT
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via5_0

VIA via6_0 DEFAULT
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END via6_0

VIA via7_0 DEFAULT
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END via7_0

VIA via8_0 DEFAULT
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END via8_0

VIA via9_0 DEFAULT
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER metal9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER metal10 ;
    RECT -0.4 -0.4 0.4 0.4 ;
END via9_0

VIARULE Via1Array-0 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER metal2 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-0

VIARULE Via1Array-1 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-1

VIARULE Via1Array-2 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0.035 0 ;
  LAYER metal2 ;
    ENCLOSURE 0.035 0 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-2

VIARULE Via1Array-3 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal2 ;
    ENCLOSURE 0.035 0 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-3

VIARULE Via1Array-4 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0.035 0 ;
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER via1 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.15 BY 0.15 ;
END Via1Array-4

VIARULE Via2Array-0 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER metal3 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-0

VIARULE Via2Array-1 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-1

VIARULE Via2Array-2 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0.035 0 ;
  LAYER metal3 ;
    ENCLOSURE 0.035 0 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-2

VIARULE Via2Array-3 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal3 ;
    ENCLOSURE 0.035 0 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-3

VIARULE Via2Array-4 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0.035 0 ;
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER via2 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via2Array-4

VIARULE Via3Array-0 GENERATE
  LAYER metal3 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER metal4 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via3Array-0

VIARULE Via3Array-1 GENERATE
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal4 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via3Array-1

VIARULE Via3Array-2 GENERATE
  LAYER metal3 ;
    ENCLOSURE 0.035 0 ;
  LAYER metal4 ;
    ENCLOSURE 0.035 0.035 ;
  LAYER via3 ;
    RECT -0.035 -0.035 0.035 0.035 ;
    SPACING 0.16 BY 0.16 ;
END Via3Array-2

VIARULE Via4Array-0 GENERATE
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via4Array-0

VIARULE Via5Array-0 GENERATE
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via5Array-0

VIARULE Via6Array-0 GENERATE
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER metal7 ;
    ENCLOSURE 0.13 0.13 ;
  LAYER via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.3 BY 0.3 ;
END Via6Array-0

VIARULE Via7Array-0 GENERATE
  LAYER metal7 ;
    ENCLOSURE 0 0 ;
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER via7 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via7Array-0

VIARULE Via8Array-0 GENERATE
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER metal9 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER via8 ;
    RECT -0.2 -0.2 0.2 0.2 ;
    SPACING 0.84 BY 0.84 ;
END Via8Array-0

VIARULE Via9Array-0 GENERATE
  LAYER metal10 ;
    ENCLOSURE 0 0 ;
  LAYER metal9 ;
    ENCLOSURE 0 0 ;
  LAYER via9 ;
    RECT -0.4 -0.4 0.4 0.4 ;
    SPACING 1.68 BY 1.68 ;
END Via9Array-0

SPACING
  SAMENET metal1 metal1 0.065 ;
  SAMENET metal2 metal2 0.07 ;
  SAMENET metal3 metal3 0.07 ;
  SAMENET metal4 metal4 0.14 ;
  SAMENET metal5 metal5 0.14 ;
  SAMENET metal6 metal6 0.14 ;
  SAMENET metal7 metal7 0.4 ;
  SAMENET metal8 metal8 0.4 ;
  SAMENET metal9 metal9 0.8 ;
  SAMENET metal10 metal10 0.8 ;
  SAMENET via1 via1 0.08 ;
  SAMENET via2 via2 0.09 ;
  SAMENET via3 via3 0.09 ;
  SAMENET via4 via4 0.16 ;
  SAMENET via5 via5 0.16 ;
  SAMENET via6 via6 0.16 ;
  SAMENET via7 via7 0.44 ;
  SAMENET via8 via8 0.44 ;
  SAMENET via9 via9 0.88 ;
  SAMENET via1 via2 0.0 STACK ;
  SAMENET via2 via3 0.0 STACK ;
  SAMENET via3 via4 0.0 STACK ;
  SAMENET via4 via5 0.0 STACK ;
  SAMENET via5 via6 0.0 STACK ;
  SAMENET via6 via7 0.0 STACK ;
  SAMENET via7 via8 0.0 STACK ;
  SAMENET via8 via9 0.0 STACK ;
END SPACING

SITE FreePDK45_38x28_10R_NP_162NW_34O
  SYMMETRY y ;
  CLASS core ;
  SIZE 0.19 BY 1.4 ;
END FreePDK45_38x28_10R_NP_162NW_34O

# END LIBRARY
#
# End of file
#




#VERSION 5.6 ;
#BUSBITCHARS "[]" ;
#DIVIDERCHAR "/" ;

MACRO AND2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_X1 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.38 0.7 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.61 0.19 0.7 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
        RECT 0.415 0.975 0.485 1.485 ;
        RECT 0.04 0.975 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
        RECT 0.415 -0.085 0.485 0.325 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.235 0.84 0.305 1.25 ;
      RECT 0.235 0.84 0.54 0.91 ;
      RECT 0.47 0.39 0.54 0.91 ;
      RECT 0.045 0.39 0.54 0.46 ;
      RECT 0.045 0.19 0.115 0.46 ;
  END
END AND2_X1

MACRO AND2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_X2 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.38 0.7 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.615 0.15 0.7 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.95 1.485 ;
        RECT 0.795 0.975 0.865 1.485 ;
        RECT 0.415 0.975 0.485 1.485 ;
        RECT 0.04 0.975 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.95 0.085 ;
        RECT 0.795 -0.085 0.865 0.425 ;
        RECT 0.415 -0.085 0.485 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.235 0.84 0.305 1.25 ;
      RECT 0.235 0.84 0.545 0.91 ;
      RECT 0.475 0.39 0.545 0.91 ;
      RECT 0.045 0.39 0.545 0.46 ;
      RECT 0.045 0.15 0.115 0.46 ;
  END
END AND2_X2

MACRO AND2_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_X4 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.42 0.38 0.66 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.725 0.76 0.795 ;
        RECT 0.69 0.525 0.76 0.795 ;
        RECT 0.06 0.42 0.185 0.795 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.365 0.15 1.435 1.25 ;
        RECT 0.995 0.68 1.435 0.75 ;
        RECT 0.995 0.15 1.08 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.71 1.485 ;
        RECT 1.555 0.995 1.625 1.485 ;
        RECT 1.175 0.995 1.245 1.485 ;
        RECT 0.795 0.995 0.865 1.485 ;
        RECT 0.415 0.995 0.485 1.485 ;
        RECT 0.04 0.995 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.71 0.085 ;
        RECT 1.555 -0.085 1.625 0.355 ;
        RECT 1.175 -0.085 1.245 0.355 ;
        RECT 0.795 -0.085 0.865 0.215 ;
        RECT 0.04 -0.085 0.11 0.355 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.605 0.86 0.675 1.25 ;
      RECT 0.235 0.86 0.305 1.25 ;
      RECT 0.235 0.86 0.92 0.93 ;
      RECT 0.85 0.285 0.92 0.93 ;
      RECT 0.425 0.285 0.92 0.355 ;
      RECT 0.425 0.22 0.495 0.355 ;
  END
END AND2_X4

MACRO AND3_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3_X1 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.375 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.57 0.7 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.8 0.975 0.89 1.25 ;
        RECT 0.82 0.15 0.89 1.25 ;
        RECT 0.8 0.15 0.89 0.425 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.95 1.485 ;
        RECT 0.605 1 0.675 1.485 ;
        RECT 0.225 1.04 0.295 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.95 0.085 ;
        RECT 0.605 -0.085 0.675 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.415 0.865 0.485 1.25 ;
      RECT 0.045 0.865 0.115 1.25 ;
      RECT 0.045 0.865 0.705 0.935 ;
      RECT 0.635 0.35 0.705 0.935 ;
      RECT 0.635 0.525 0.755 0.66 ;
      RECT 0.045 0.35 0.705 0.42 ;
      RECT 0.045 0.15 0.115 0.42 ;
  END
END AND3_X1

MACRO AND3_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3_X2 0 0 ;
  SIZE 1.14 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.375 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.57 0.7 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.805 0.15 0.89 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.14 1.485 ;
        RECT 0.99 0.975 1.06 1.485 ;
        RECT 0.605 0.975 0.675 1.485 ;
        RECT 0.225 0.975 0.295 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.14 0.085 ;
        RECT 0.99 -0.085 1.06 0.425 ;
        RECT 0.605 -0.085 0.675 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.415 0.8 0.485 1.25 ;
      RECT 0.045 0.8 0.115 1.25 ;
      RECT 0.045 0.8 0.735 0.87 ;
      RECT 0.665 0.355 0.735 0.87 ;
      RECT 0.045 0.355 0.735 0.425 ;
      RECT 0.045 0.15 0.115 0.425 ;
  END
END AND3_X2

MACRO AND3_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3_X4 0 0 ;
  SIZE 2.09 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.595 0.555 0.73 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.82 0.42 0.95 0.7 ;
        RECT 0.34 0.42 0.95 0.49 ;
        RECT 0.34 0.42 0.41 0.66 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.12 0.765 1.14 0.835 ;
        RECT 1.07 0.525 1.14 0.835 ;
        RECT 0.12 0.525 0.19 0.835 ;
        RECT 0.06 0.525 0.19 0.7 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.745 0.15 1.815 1.25 ;
        RECT 1.375 0.56 1.815 0.7 ;
        RECT 1.375 0.15 1.445 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.09 1.485 ;
        RECT 1.935 1.035 2.005 1.485 ;
        RECT 1.555 1.035 1.625 1.485 ;
        RECT 1.175 1.035 1.245 1.485 ;
        RECT 0.795 1.035 0.865 1.485 ;
        RECT 0.415 1.035 0.485 1.485 ;
        RECT 0.04 1.035 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.09 0.085 ;
        RECT 1.935 -0.085 2.005 0.425 ;
        RECT 1.555 -0.085 1.625 0.425 ;
        RECT 1.175 -0.085 1.245 0.195 ;
        RECT 0.04 -0.085 0.11 0.425 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.985 0.9 1.055 1.25 ;
      RECT 0.605 0.9 0.675 1.25 ;
      RECT 0.235 0.9 0.305 1.25 ;
      RECT 0.235 0.9 1.305 0.97 ;
      RECT 1.235 0.26 1.305 0.97 ;
      RECT 0.615 0.26 1.305 0.33 ;
      RECT 0.615 0.15 0.685 0.33 ;
  END
END AND3_X4

MACRO AND4_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4_X1 0 0 ;
  SIZE 1.14 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.375 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.565 0.7 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.525 0.76 0.7 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.99 0.15 1.08 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.14 1.485 ;
        RECT 0.795 0.975 0.865 1.485 ;
        RECT 0.415 0.975 0.485 1.485 ;
        RECT 0.04 0.975 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.14 0.085 ;
        RECT 0.795 -0.085 0.865 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.605 0.84 0.675 1.25 ;
      RECT 0.235 0.84 0.305 1.25 ;
      RECT 0.235 0.84 0.925 0.91 ;
      RECT 0.855 0.35 0.925 0.91 ;
      RECT 0.045 0.35 0.925 0.42 ;
      RECT 0.045 0.15 0.115 0.42 ;
  END
END AND4_X1

MACRO AND4_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4_X2 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.375 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.565 0.7 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.525 0.76 0.7 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.995 0.15 1.08 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.33 1.485 ;
        RECT 1.18 0.975 1.25 1.485 ;
        RECT 0.795 0.975 0.865 1.485 ;
        RECT 0.415 0.975 0.485 1.485 ;
        RECT 0.04 0.975 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.33 0.085 ;
        RECT 1.18 -0.085 1.25 0.425 ;
        RECT 0.795 -0.085 0.865 0.27 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.605 0.8 0.675 1.25 ;
      RECT 0.235 0.8 0.305 1.25 ;
      RECT 0.235 0.8 0.925 0.87 ;
      RECT 0.855 0.355 0.925 0.87 ;
      RECT 0.045 0.355 0.925 0.425 ;
      RECT 0.045 0.15 0.115 0.425 ;
  END
END AND4_X2

MACRO AND4_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4_X4 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.8 0.56 0.935 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.065 0.425 1.135 0.66 ;
        RECT 0.565 0.425 1.135 0.495 ;
        RECT 0.565 0.425 0.7 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.355 0.77 1.345 0.84 ;
        RECT 1.2 0.525 1.345 0.84 ;
        RECT 0.355 0.525 0.425 0.84 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.135 0.905 1.535 0.975 ;
        RECT 1.465 0.525 1.535 0.975 ;
        RECT 0.135 0.525 0.205 0.975 ;
        RECT 0.06 0.525 0.205 0.7 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.14 0.15 2.21 0.925 ;
        RECT 1.77 0.56 2.21 0.7 ;
        RECT 1.77 0.15 1.84 0.925 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.47 1.485 ;
        RECT 2.33 1.065 2.4 1.485 ;
        RECT 1.95 1.065 2.02 1.485 ;
        RECT 1.57 1.175 1.64 1.485 ;
        RECT 1.19 1.175 1.26 1.485 ;
        RECT 0.81 1.175 0.88 1.485 ;
        RECT 0.43 1.175 0.5 1.485 ;
        RECT 0.055 1.065 0.125 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.47 0.085 ;
        RECT 2.33 -0.085 2.4 0.425 ;
        RECT 1.95 -0.085 2.02 0.425 ;
        RECT 1.57 -0.085 1.64 0.195 ;
        RECT 0.055 -0.085 0.125 0.425 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.215 1.04 1.705 1.11 ;
      RECT 1.635 0.29 1.705 1.11 ;
      RECT 0.785 0.29 1.705 0.36 ;
  END
END AND4_X4

MACRO ANTENNA_X1
  CLASS CORE ANTENNACELL ;
  ORIGIN 0 0 ;
  FOREIGN ANTENNA_X1 0 0 ;
  SIZE 0.19 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    # unknown
    ANTENNADIFFAREA  0.0 ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.42 0.13 0.75 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.19 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.19 0.085 ;
    END
  END VSS
END ANTENNA_X1

MACRO AOI211_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211_X1 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765 0.525 0.89 0.7 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.575 0.525 0.7 0.7 ;
    END
  END B
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.41 0.525 0.51 0.7 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.21 0.7 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.275 0.355 0.905 0.425 ;
        RECT 0.835 0.15 0.905 0.425 ;
        RECT 0.44 0.15 0.525 0.425 ;
        RECT 0.275 0.355 0.345 1.115 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.95 1.485 ;
        RECT 0.835 0.905 0.905 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.95 0.085 ;
        RECT 0.645 -0.085 0.715 0.285 ;
        RECT 0.08 -0.085 0.15 0.425 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.085 1.18 0.525 1.25 ;
      RECT 0.455 0.905 0.525 1.25 ;
      RECT 0.085 0.905 0.155 1.25 ;
  END
END AOI211_X1

MACRO AOI211_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211_X2 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.39 0.56 0.525 0.7 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.765 0.75 0.835 ;
        RECT 0.68 0.525 0.75 0.835 ;
        RECT 0.06 0.525 0.185 0.835 ;
    END
  END B
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.19 0.56 1.325 0.7 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.54 0.425 1.65 0.7 ;
        RECT 0.965 0.425 1.65 0.495 ;
        RECT 0.965 0.425 1.035 0.66 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.405 0.765 1.475 1.055 ;
        RECT 0.82 0.765 1.475 0.835 ;
        RECT 0.2 0.285 1.32 0.355 ;
        RECT 1.185 0.15 1.32 0.355 ;
        RECT 1.025 0.765 1.095 1.055 ;
        RECT 0.82 0.285 0.89 0.835 ;
        RECT 0.2 0.15 0.335 0.355 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.71 1.485 ;
        RECT 0.42 1.035 0.49 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.71 0.085 ;
        RECT 1.595 -0.085 1.665 0.355 ;
        RECT 0.825 -0.085 0.895 0.215 ;
        RECT 0.43 -0.085 0.5 0.215 ;
        RECT 0.045 -0.085 0.115 0.355 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.815 1.18 1.665 1.25 ;
      RECT 1.595 0.975 1.665 1.25 ;
      RECT 0.05 0.9 0.12 1.25 ;
      RECT 1.22 0.975 1.29 1.25 ;
      RECT 0.815 0.9 0.885 1.25 ;
      RECT 0.05 0.9 0.885 0.97 ;
  END
END AOI211_X2

MACRO AOI211_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211_X4 0 0 ;
  SIZE 2.09 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.525 0.76 0.7 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.565 0.7 ;
    END
  END B
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.375 0.7 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.75 0.15 1.82 1.175 ;
        RECT 1.375 0.56 1.82 0.7 ;
        RECT 1.375 0.15 1.445 1.175 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.09 1.485 ;
        RECT 1.935 0.9 2.005 1.485 ;
        RECT 1.555 0.9 1.625 1.485 ;
        RECT 1.175 0.9 1.245 1.485 ;
        RECT 0.795 0.9 0.865 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.09 0.085 ;
        RECT 1.935 -0.085 2.005 0.425 ;
        RECT 1.555 -0.085 1.625 0.425 ;
        RECT 1.175 -0.085 1.245 0.425 ;
        RECT 0.795 -0.085 0.865 0.285 ;
        RECT 0.415 -0.085 0.485 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.995 0.15 1.065 1.175 ;
      RECT 0.995 0.525 1.31 0.66 ;
      RECT 0.235 0.765 0.305 1.115 ;
      RECT 0.235 0.765 0.93 0.835 ;
      RECT 0.86 0.39 0.93 0.835 ;
      RECT 0.045 0.39 0.93 0.46 ;
      RECT 0.605 0.15 0.675 0.46 ;
      RECT 0.045 0.15 0.115 0.46 ;
      RECT 0.045 1.18 0.485 1.25 ;
      RECT 0.415 0.9 0.485 1.25 ;
      RECT 0.045 0.9 0.115 1.25 ;
  END
END AOI211_X4

MACRO AOI21_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21_X1 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.575 0.525 0.7 0.7 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.4 0.525 0.51 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.2 0.7 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.265 0.355 0.525 0.425 ;
        RECT 0.44 0.15 0.525 0.425 ;
        RECT 0.265 0.355 0.335 1.115 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
        RECT 0.645 0.905 0.715 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
        RECT 0.645 -0.085 0.715 0.355 ;
        RECT 0.08 -0.085 0.15 0.425 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.085 1.18 0.525 1.25 ;
      RECT 0.455 0.905 0.525 1.25 ;
      RECT 0.085 0.905 0.155 1.25 ;
  END
END AOI21_X1

MACRO AOI21_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21_X2 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.215 0.56 0.35 0.7 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765 0.56 0.9 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.77 1.18 0.84 ;
        RECT 1.11 0.525 1.18 0.84 ;
        RECT 0.63 0.525 0.7 0.84 ;
        RECT 0.57 0.525 0.7 0.7 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.435 0.905 1.13 0.975 ;
        RECT 0.25 0.355 0.905 0.425 ;
        RECT 0.835 0.15 0.905 0.425 ;
        RECT 0.435 0.355 0.505 0.975 ;
        RECT 0.25 0.15 0.335 0.425 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.33 1.485 ;
        RECT 0.265 1.205 0.335 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.33 0.085 ;
        RECT 1.215 -0.085 1.285 0.425 ;
        RECT 0.455 -0.085 0.525 0.285 ;
        RECT 0.08 -0.085 0.15 0.425 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.215 0.975 1.285 1.25 ;
      RECT 0.085 0.975 0.155 1.25 ;
      RECT 0.085 1.07 1.285 1.14 ;
  END
END AOI21_X2

MACRO AOI21_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21_X4 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.4 0.525 0.535 0.7 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.165 0.69 2.06 0.76 ;
        RECT 1.925 0.56 2.06 0.76 ;
        RECT 1.165 0.56 1.3 0.76 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.25 0.42 2.32 0.66 ;
        RECT 0.925 0.42 2.32 0.49 ;
        RECT 1.525 0.42 1.66 0.625 ;
        RECT 0.925 0.42 0.995 0.66 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.14 0.825 2.21 1.115 ;
        RECT 0.63 0.825 2.21 0.895 ;
        RECT 0.63 0.26 2.055 0.33 ;
        RECT 1.76 0.825 1.83 1.115 ;
        RECT 1.38 0.825 1.45 1.115 ;
        RECT 1 0.825 1.07 1.115 ;
        RECT 0.63 0.15 0.7 0.895 ;
        RECT 0.25 0.355 0.7 0.425 ;
        RECT 0.25 0.15 0.32 0.425 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.47 1.485 ;
        RECT 0.62 1.205 0.69 1.485 ;
        RECT 0.24 1.205 0.31 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.47 0.085 ;
        RECT 2.33 -0.085 2.4 0.35 ;
        RECT 1.57 -0.085 1.64 0.195 ;
        RECT 0.81 -0.085 0.88 0.195 ;
        RECT 0.43 -0.085 0.5 0.195 ;
        RECT 0.055 -0.085 0.125 0.425 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.81 1.18 2.4 1.25 ;
      RECT 2.33 0.84 2.4 1.25 ;
      RECT 0.43 0.965 0.5 1.24 ;
      RECT 0.06 0.965 0.13 1.24 ;
      RECT 1.95 0.96 2.02 1.25 ;
      RECT 1.57 0.96 1.64 1.25 ;
      RECT 1.19 0.96 1.26 1.25 ;
      RECT 0.81 0.965 0.88 1.25 ;
      RECT 0.06 0.965 0.88 1.035 ;
  END
END AOI21_X4

MACRO AOI221_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221_X1 0 0 ;
  SIZE 1.14 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.565 0.7 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.375 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.955 0.525 1.08 0.7 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.525 0.74 0.7 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425 0.355 1.055 0.425 ;
        RECT 0.985 0.15 1.055 0.425 ;
        RECT 0.805 0.355 0.89 1.115 ;
        RECT 0.425 0.15 0.495 0.425 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.14 1.485 ;
        RECT 0.225 0.905 0.295 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.14 0.085 ;
        RECT 0.605 -0.085 0.675 0.215 ;
        RECT 0.04 -0.085 0.11 0.355 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.615 1.18 1.055 1.25 ;
      RECT 0.985 0.905 1.055 1.25 ;
      RECT 0.615 0.905 0.685 1.25 ;
      RECT 0.415 0.77 0.485 1.18 ;
      RECT 0.045 0.77 0.115 1.18 ;
      RECT 0.045 0.77 0.485 0.84 ;
  END
END AOI221_X1

MACRO AOI221_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221_X2 0 0 ;
  SIZE 2.09 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.18 0.79 1.13 0.86 ;
        RECT 1.06 0.525 1.13 0.86 ;
        RECT 0.18 0.56 0.25 0.86 ;
        RECT 0.06 0.56 0.25 0.7 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.82 0.42 0.945 0.7 ;
        RECT 0.34 0.42 0.945 0.49 ;
        RECT 0.34 0.42 0.41 0.66 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.585 0.56 0.725 0.7 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.57 0.525 1.66 0.7 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.77 0.525 1.91 0.7 ;
        RECT 1.34 0.765 1.84 0.835 ;
        RECT 1.77 0.525 1.84 0.835 ;
        RECT 1.34 0.525 1.41 0.835 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.195 0.9 1.86 0.97 ;
        RECT 0.2 0.28 1.675 0.35 ;
        RECT 1.195 0.28 1.275 0.97 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.09 1.485 ;
        RECT 0.795 1.205 0.865 1.485 ;
        RECT 0.415 1.205 0.485 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.09 0.085 ;
        RECT 1.945 -0.085 2.015 0.425 ;
        RECT 1.175 -0.085 1.245 0.195 ;
        RECT 0.605 -0.085 0.675 0.195 ;
        RECT 0.04 -0.085 0.11 0.425 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 1.07 2.015 1.14 ;
      RECT 1.945 0.865 2.015 1.14 ;
      RECT 0.045 0.865 0.115 1.14 ;
      RECT 0.2 0.93 1.09 1 ;
  END
END AOI221_X2

MACRO AOI221_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221_X4 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.61 0.525 0.7 0.7 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.8 0.525 0.89 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.01 0.525 1.18 0.7 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.27 0.7 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.42 0.525 0.51 0.7 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.17 0.15 2.24 1.25 ;
        RECT 1.795 0.56 2.24 0.7 ;
        RECT 1.795 0.15 1.885 0.7 ;
        RECT 1.795 0.15 1.865 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.47 1.485 ;
        RECT 2.355 0.975 2.425 1.485 ;
        RECT 1.975 0.975 2.045 1.485 ;
        RECT 1.6 1.005 1.67 1.485 ;
        RECT 1.215 0.975 1.285 1.485 ;
        RECT 0.875 1.035 0.945 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.47 0.085 ;
        RECT 2.355 -0.085 2.425 0.425 ;
        RECT 1.975 -0.085 2.045 0.425 ;
        RECT 1.605 -0.085 1.675 0.425 ;
        RECT 1.215 -0.085 1.285 0.285 ;
        RECT 0.495 -0.085 0.565 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.415 0.15 1.485 1.25 ;
      RECT 1.415 0.525 1.73 0.66 ;
      RECT 0.315 0.765 0.385 1.04 ;
      RECT 0.315 0.765 1.35 0.835 ;
      RECT 1.28 0.355 1.35 0.835 ;
      RECT 0.125 0.355 1.35 0.425 ;
      RECT 0.71 0.15 0.78 0.425 ;
      RECT 0.125 0.15 0.195 0.425 ;
      RECT 1.03 0.9 1.1 1.25 ;
      RECT 0.695 0.9 0.765 1.25 ;
      RECT 0.695 0.9 1.1 0.97 ;
      RECT 0.495 0.975 0.565 1.25 ;
      RECT 0.125 0.975 0.195 1.25 ;
      RECT 0.125 1.105 0.565 1.175 ;
  END
END AOI221_X4

MACRO AOI222_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222_X1 0 0 ;
  SIZE 1.52 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.315 0.525 1.46 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.995 0.525 1.08 0.7 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.62 0.525 0.72 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.82 0.525 0.91 0.7 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.385 0.525 0.51 0.7 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.215 0.7 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.5 0.375 1.46 0.45 ;
        RECT 1.325 0.175 1.46 0.45 ;
        RECT 1.145 0.375 1.215 1.115 ;
        RECT 0.5 0.175 0.57 0.45 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.52 1.485 ;
        RECT 0.415 0.905 0.485 1.485 ;
        RECT 0.04 0.905 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.52 0.085 ;
        RECT 0.945 -0.085 1.015 0.31 ;
        RECT 0.04 -0.085 0.11 0.45 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.575 1.18 1.395 1.25 ;
      RECT 1.325 0.905 1.395 1.25 ;
      RECT 0.945 0.905 1.015 1.25 ;
      RECT 0.575 0.905 0.645 1.25 ;
      RECT 0.235 0.77 0.305 1.18 ;
      RECT 0.755 0.77 0.825 1.115 ;
      RECT 0.235 0.77 0.825 0.84 ;
  END
END AOI222_X1

MACRO AOI222_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222_X2 0 0 ;
  SIZE 2.66 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.91 0.56 2.045 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.285 0.56 2.42 0.7 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.145 0.56 1.28 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.475 0.42 1.545 0.66 ;
        RECT 0.91 0.42 1.545 0.49 ;
        RECT 0.91 0.42 1.08 0.66 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.385 0.56 0.52 0.7 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.69 0.425 0.76 0.66 ;
        RECT 0.06 0.425 0.76 0.495 ;
        RECT 0.06 0.425 0.19 0.7 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.31 0.77 2.38 1.115 ;
        RECT 1.77 0.77 2.38 0.84 ;
        RECT 0.39 0.285 2.035 0.355 ;
        RECT 1.94 0.77 2.01 1.115 ;
        RECT 1.77 0.285 1.84 0.84 ;
        RECT 1.145 0.15 1.28 0.355 ;
        RECT 0.39 0.15 0.525 0.355 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.66 1.485 ;
        RECT 0.605 0.905 0.675 1.485 ;
        RECT 0.225 0.905 0.295 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.66 0.085 ;
        RECT 2.31 -0.085 2.38 0.25 ;
        RECT 1.555 -0.085 1.625 0.195 ;
        RECT 0.765 -0.085 0.9 0.215 ;
        RECT 0.04 -0.085 0.11 0.25 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 2.1 0.355 2.57 0.425 ;
      RECT 2.5 0.15 2.57 0.425 ;
      RECT 2.1 0.15 2.17 0.425 ;
      RECT 1.715 0.15 2.17 0.22 ;
      RECT 0.995 1.18 2.57 1.25 ;
      RECT 2.5 0.905 2.57 1.25 ;
      RECT 2.12 0.905 2.19 1.25 ;
      RECT 1.745 0.905 1.815 1.25 ;
      RECT 1.365 0.905 1.435 1.25 ;
      RECT 0.995 0.905 1.065 1.25 ;
      RECT 0.795 0.77 0.865 1.18 ;
      RECT 0.415 0.77 0.485 1.18 ;
      RECT 0.045 0.77 0.115 1.18 ;
      RECT 1.555 0.77 1.625 1.115 ;
      RECT 1.175 0.77 1.245 1.115 ;
      RECT 0.045 0.77 1.625 0.84 ;
  END
END AOI222_X2

MACRO AOI222_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222_X4 0 0 ;
  SIZE 2.66 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.235 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.385 0.525 0.51 0.7 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765 0.525 0.89 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.575 0.525 0.7 0.7 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.01 0.525 1.135 0.7 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.2 0.525 1.335 0.7 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.33 0.15 2.41 1.205 ;
        RECT 1.95 0.56 2.41 0.7 ;
        RECT 2.325 0.15 2.41 0.7 ;
        RECT 1.95 0.15 2.02 1.205 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.66 1.485 ;
        RECT 2.51 0.93 2.58 1.485 ;
        RECT 2.13 0.93 2.2 1.485 ;
        RECT 1.75 0.93 1.82 1.485 ;
        RECT 1.37 0.93 1.44 1.485 ;
        RECT 0.995 1.065 1.065 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.66 0.085 ;
        RECT 2.51 -0.085 2.58 0.425 ;
        RECT 2.14 -0.085 2.21 0.425 ;
        RECT 1.75 -0.085 1.82 0.425 ;
        RECT 1.37 -0.085 1.44 0.285 ;
        RECT 0.46 -0.085 0.53 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.57 0.15 1.64 1.205 ;
      RECT 1.57 0.525 1.885 0.66 ;
      RECT 0.28 0.765 0.35 1.04 ;
      RECT 0.28 0.765 1.505 0.835 ;
      RECT 1.435 0.355 1.505 0.835 ;
      RECT 0.09 0.355 1.505 0.425 ;
      RECT 0.84 0.15 0.91 0.425 ;
      RECT 0.09 0.15 0.16 0.425 ;
      RECT 1.18 0.93 1.25 1.205 ;
      RECT 0.66 0.93 0.73 1.065 ;
      RECT 0.66 0.93 1.25 1 ;
      RECT 0.09 1.135 0.91 1.205 ;
      RECT 0.84 1.07 0.91 1.205 ;
      RECT 0.46 0.93 0.53 1.205 ;
      RECT 0.09 0.93 0.16 1.205 ;
  END
END AOI222_X4

MACRO AOI22_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22_X1 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.575 0.42 0.7 0.66 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765 0.42 0.89 0.66 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.375 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.62 0.725 0.69 1.005 ;
        RECT 0.44 0.725 0.69 0.795 ;
        RECT 0.44 0.15 0.51 0.795 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.95 1.485 ;
        RECT 0.24 1.205 0.31 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.95 0.085 ;
        RECT 0.81 -0.085 0.88 0.355 ;
        RECT 0.055 -0.085 0.125 0.355 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.06 1.07 0.88 1.14 ;
      RECT 0.81 0.865 0.88 1.14 ;
      RECT 0.435 0.865 0.505 1.14 ;
      RECT 0.06 0.865 0.13 1.14 ;
  END
END AOI22_X1

MACRO AOI22_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22_X2 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.155 0.56 1.29 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.48 0.425 1.55 0.66 ;
        RECT 0.955 0.425 1.55 0.495 ;
        RECT 0.955 0.425 1.08 0.7 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.395 0.56 0.53 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.765 0.755 0.835 ;
        RECT 0.685 0.525 0.755 0.835 ;
        RECT 0.06 0.525 0.195 0.835 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.375 0.765 1.445 1.065 ;
        RECT 0.82 0.765 1.445 0.835 ;
        RECT 0.395 0.28 1.285 0.355 ;
        RECT 1.15 0.15 1.285 0.355 ;
        RECT 0.99 0.765 1.06 1.065 ;
        RECT 0.82 0.28 0.89 0.835 ;
        RECT 0.395 0.15 0.53 0.355 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.71 1.485 ;
        RECT 0.61 1.035 0.68 1.485 ;
        RECT 0.23 1.035 0.3 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.71 0.085 ;
        RECT 1.56 -0.085 1.63 0.36 ;
        RECT 0.77 -0.085 0.905 0.205 ;
        RECT 0.045 -0.085 0.115 0.39 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.8 1.18 1.63 1.25 ;
      RECT 1.56 0.975 1.63 1.25 ;
      RECT 0.42 0.9 0.49 1.25 ;
      RECT 0.05 0.9 0.12 1.25 ;
      RECT 1.18 0.975 1.25 1.25 ;
      RECT 0.8 0.9 0.87 1.25 ;
      RECT 0.05 0.9 0.87 0.97 ;
  END
END AOI22_X2

MACRO AOI22_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22_X4 0 0 ;
  SIZE 3.23 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.915 0.69 2.79 0.76 ;
        RECT 2.655 0.56 2.79 0.76 ;
        RECT 1.915 0.56 2.05 0.76 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.91 0.42 3.045 0.66 ;
        RECT 1.715 0.42 3.045 0.49 ;
        RECT 2.295 0.42 2.43 0.625 ;
        RECT 1.715 0.42 1.785 0.66 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.395 0.69 1.29 0.76 ;
        RECT 1.155 0.56 1.29 0.76 ;
        RECT 0.395 0.56 0.53 0.76 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.445 0.42 1.515 0.66 ;
        RECT 0.125 0.42 1.515 0.49 ;
        RECT 0.755 0.42 0.89 0.625 ;
        RECT 0.125 0.42 0.195 0.66 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.89 0.825 2.96 1.115 ;
        RECT 1.75 0.825 2.96 0.895 ;
        RECT 0.395 0.26 2.805 0.33 ;
        RECT 2.51 0.825 2.58 1.115 ;
        RECT 2.13 0.825 2.2 1.115 ;
        RECT 1.75 0.725 1.82 1.115 ;
        RECT 1.58 0.725 1.82 0.795 ;
        RECT 1.58 0.26 1.65 0.795 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 3.23 1.485 ;
        RECT 1.37 1.065 1.44 1.485 ;
        RECT 0.99 1.065 1.06 1.485 ;
        RECT 0.61 1.065 0.68 1.485 ;
        RECT 0.23 1.065 0.3 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 3.23 0.085 ;
        RECT 3.08 -0.085 3.15 0.335 ;
        RECT 2.29 -0.085 2.425 0.16 ;
        RECT 1.53 -0.085 1.665 0.16 ;
        RECT 0.77 -0.085 0.905 0.16 ;
        RECT 0.045 -0.085 0.115 0.335 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.56 1.18 3.15 1.25 ;
      RECT 3.08 0.84 3.15 1.25 ;
      RECT 2.7 0.96 2.77 1.25 ;
      RECT 2.32 0.96 2.39 1.25 ;
      RECT 1.94 0.96 2.01 1.25 ;
      RECT 1.56 0.87 1.63 1.25 ;
      RECT 1.18 0.87 1.25 1.16 ;
      RECT 0.8 0.87 0.87 1.16 ;
      RECT 0.42 0.87 0.49 1.16 ;
      RECT 0.05 0.87 0.12 1.16 ;
      RECT 0.05 0.87 1.63 0.94 ;
  END
END AOI22_X4

MACRO BUF_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X1 0 0 ;
  SIZE 0.57 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.19 0.7 ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.42 0.19 0.51 1.24 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.57 1.485 ;
        RECT 0.225 0.965 0.295 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.57 0.085 ;
        RECT 0.225 -0.085 0.295 0.325 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.83 0.115 1.24 ;
      RECT 0.045 0.83 0.355 0.9 ;
      RECT 0.285 0.39 0.355 0.9 ;
      RECT 0.045 0.39 0.355 0.46 ;
      RECT 0.045 0.19 0.115 0.46 ;
  END
END BUF_X1

MACRO BUF_X16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X16 0 0 ;
  SIZE 4.75 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.715 ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.42 0.15 4.49 0.925 ;
        RECT 1.77 0.28 4.49 0.42 ;
        RECT 4.05 0.28 4.12 0.925 ;
        RECT 4.04 0.15 4.11 0.42 ;
        RECT 3.66 0.15 3.73 0.925 ;
        RECT 3.28 0.15 3.35 0.925 ;
        RECT 2.9 0.15 2.97 0.925 ;
        RECT 2.52 0.15 2.59 0.925 ;
        RECT 2.14 0.15 2.21 0.925 ;
        RECT 1.77 0.15 1.84 0.925 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 4.75 1.485 ;
        RECT 4.61 1.205 4.68 1.485 ;
        RECT 4.23 1.205 4.3 1.485 ;
        RECT 3.85 1.205 3.92 1.485 ;
        RECT 3.47 1.205 3.54 1.485 ;
        RECT 3.09 1.205 3.16 1.485 ;
        RECT 2.71 1.205 2.78 1.485 ;
        RECT 2.33 1.205 2.4 1.485 ;
        RECT 1.95 1.205 2.02 1.485 ;
        RECT 1.57 1.205 1.64 1.485 ;
        RECT 1.19 0.975 1.26 1.485 ;
        RECT 0.81 0.975 0.88 1.485 ;
        RECT 0.43 0.975 0.5 1.485 ;
        RECT 0.055 0.975 0.125 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 4.75 0.085 ;
        RECT 4.61 -0.085 4.68 0.2 ;
        RECT 4.23 -0.085 4.3 0.2 ;
        RECT 3.85 -0.085 3.92 0.2 ;
        RECT 3.47 -0.085 3.54 0.2 ;
        RECT 3.09 -0.085 3.16 0.2 ;
        RECT 2.71 -0.085 2.78 0.2 ;
        RECT 2.33 -0.085 2.4 0.2 ;
        RECT 1.95 -0.085 2.02 0.2 ;
        RECT 1.57 -0.085 1.64 0.34 ;
        RECT 1.19 -0.085 1.26 0.34 ;
        RECT 0.81 -0.085 0.88 0.34 ;
        RECT 0.43 -0.085 0.5 0.34 ;
        RECT 0.055 -0.085 0.125 0.34 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.38 0.15 1.45 1.25 ;
      RECT 1 0.15 1.07 1.25 ;
      RECT 0.62 0.15 0.69 1.25 ;
      RECT 0.25 0.15 0.32 1.25 ;
      RECT 1.635 1.05 4.63 1.12 ;
      RECT 4.56 0.525 4.63 1.12 ;
      RECT 3.45 0.525 3.52 1.12 ;
      RECT 2.69 0.525 2.76 1.12 ;
      RECT 1.635 0.525 1.705 1.12 ;
      RECT 0.25 0.525 1.705 0.66 ;
  END
END BUF_X16

MACRO BUF_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X2 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.23 0.7 ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.465 0.56 0.7 0.7 ;
        RECT 0.465 0.15 0.535 1.25 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
        RECT 0.645 0.975 0.715 1.485 ;
        RECT 0.265 1.04 0.335 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
        RECT 0.645 -0.085 0.715 0.425 ;
        RECT 0.265 -0.085 0.335 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.085 0.82 0.155 1.25 ;
      RECT 0.085 0.82 0.395 0.89 ;
      RECT 0.325 0.39 0.395 0.89 ;
      RECT 0.085 0.39 0.395 0.46 ;
      RECT 0.085 0.15 0.155 0.46 ;
  END
END BUF_X2

MACRO BUF_X32
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X32 0 0 ;
  SIZE 9.31 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.1 0.93 2.8 1 ;
        RECT 2.665 0.56 2.8 1 ;
        RECT 1.905 0.56 2.04 1 ;
        RECT 1.12 0.56 1.255 1 ;
        RECT 0.1 0.525 0.17 1 ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 8.99 0.15 9.06 1.25 ;
        RECT 3.3 0.28 9.06 0.42 ;
        RECT 8.61 0.15 8.68 0.785 ;
        RECT 8.23 0.15 8.3 0.785 ;
        RECT 7.85 0.15 7.92 0.785 ;
        RECT 7.47 0.15 7.54 0.785 ;
        RECT 7.09 0.15 7.16 0.785 ;
        RECT 6.71 0.15 6.78 0.785 ;
        RECT 6.33 0.15 6.4 0.785 ;
        RECT 5.95 0.15 6.02 0.785 ;
        RECT 5.57 0.15 5.64 0.785 ;
        RECT 5.19 0.15 5.26 0.785 ;
        RECT 4.81 0.15 4.88 0.785 ;
        RECT 4.43 0.15 4.5 0.785 ;
        RECT 4.05 0.15 4.12 0.785 ;
        RECT 3.67 0.15 3.74 0.785 ;
        RECT 3.3 0.15 3.37 0.785 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 9.31 1.485 ;
        RECT 9.18 1.065 9.25 1.485 ;
        RECT 8.8 1.065 8.87 1.485 ;
        RECT 8.42 1.065 8.49 1.485 ;
        RECT 8.04 1.065 8.11 1.485 ;
        RECT 7.66 1.065 7.73 1.485 ;
        RECT 7.28 1.065 7.35 1.485 ;
        RECT 6.9 1.065 6.97 1.485 ;
        RECT 6.52 1.065 6.59 1.485 ;
        RECT 6.14 1.065 6.21 1.485 ;
        RECT 5.76 1.065 5.83 1.485 ;
        RECT 5.38 1.065 5.45 1.485 ;
        RECT 5 1.065 5.07 1.485 ;
        RECT 4.62 1.065 4.69 1.485 ;
        RECT 4.24 1.065 4.31 1.485 ;
        RECT 3.86 1.065 3.93 1.485 ;
        RECT 3.48 1.065 3.55 1.485 ;
        RECT 3.08 1.065 3.15 1.485 ;
        RECT 2.695 1.065 2.765 1.485 ;
        RECT 2.315 1.065 2.385 1.485 ;
        RECT 1.935 1.065 2.005 1.485 ;
        RECT 1.555 1.065 1.625 1.485 ;
        RECT 1.175 1.065 1.245 1.485 ;
        RECT 0.795 1.065 0.865 1.485 ;
        RECT 0.415 1.065 0.485 1.485 ;
        RECT 0.04 1.065 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 9.31 0.085 ;
        RECT 9.18 -0.085 9.25 0.2 ;
        RECT 8.8 -0.085 8.87 0.2 ;
        RECT 8.42 -0.085 8.49 0.2 ;
        RECT 8.04 -0.085 8.11 0.2 ;
        RECT 7.66 -0.085 7.73 0.2 ;
        RECT 7.28 -0.085 7.35 0.2 ;
        RECT 6.9 -0.085 6.97 0.2 ;
        RECT 6.52 -0.085 6.59 0.2 ;
        RECT 6.14 -0.085 6.21 0.2 ;
        RECT 5.76 -0.085 5.83 0.2 ;
        RECT 5.38 -0.085 5.45 0.2 ;
        RECT 5 -0.085 5.07 0.2 ;
        RECT 4.62 -0.085 4.69 0.2 ;
        RECT 4.24 -0.085 4.31 0.2 ;
        RECT 3.86 -0.085 3.93 0.2 ;
        RECT 3.48 -0.085 3.55 0.2 ;
        RECT 3.08 -0.085 3.15 0.22 ;
        RECT 2.695 -0.085 2.765 0.34 ;
        RECT 2.315 -0.085 2.385 0.34 ;
        RECT 1.935 -0.085 2.005 0.34 ;
        RECT 1.555 -0.085 1.625 0.34 ;
        RECT 1.175 -0.085 1.245 0.34 ;
        RECT 0.795 -0.085 0.865 0.34 ;
        RECT 0.415 -0.085 0.485 0.34 ;
        RECT 0.04 -0.085 0.11 0.36 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 3.165 0.85 8.88 0.92 ;
      RECT 8.745 0.56 8.88 0.92 ;
      RECT 2.885 0.405 2.955 0.865 ;
      RECT 2.505 0.15 2.575 0.865 ;
      RECT 2.13 0.15 2.2 0.865 ;
      RECT 1.745 0.405 1.815 0.865 ;
      RECT 1.365 0.15 1.435 0.865 ;
      RECT 0.985 0.15 1.055 0.865 ;
      RECT 0.615 0.405 0.685 0.865 ;
      RECT 0.235 0.15 0.305 0.865 ;
      RECT 7.605 0.56 7.74 0.92 ;
      RECT 6.465 0.56 6.6 0.92 ;
      RECT 5.325 0.56 5.46 0.92 ;
      RECT 4.185 0.56 4.32 0.92 ;
      RECT 3.165 0.405 3.235 0.92 ;
      RECT 0.235 0.405 3.235 0.495 ;
      RECT 2.89 0.15 2.96 0.495 ;
      RECT 1.75 0.15 1.82 0.495 ;
      RECT 0.605 0.15 0.675 0.495 ;
  END
END BUF_X32

MACRO BUF_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X4 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.17 0.7 ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.995 0.15 1.065 1.25 ;
        RECT 0.615 0.56 1.065 0.7 ;
        RECT 0.615 0.15 0.685 1.25 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.33 1.485 ;
        RECT 1.175 0.975 1.245 1.485 ;
        RECT 0.795 0.975 0.865 1.485 ;
        RECT 0.415 0.975 0.485 1.485 ;
        RECT 0.04 0.975 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.33 0.085 ;
        RECT 1.175 -0.085 1.245 0.37 ;
        RECT 0.795 -0.085 0.865 0.37 ;
        RECT 0.415 -0.085 0.485 0.37 ;
        RECT 0.04 -0.085 0.11 0.37 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.235 0.15 0.305 1.25 ;
      RECT 0.235 0.525 0.55 0.66 ;
  END
END BUF_X4

MACRO BUF_X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X8 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.17 0.7 ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.125 0.15 2.195 1.25 ;
        RECT 0.995 0.56 2.195 0.7 ;
        RECT 1.755 0.56 1.825 1.25 ;
        RECT 1.745 0.15 1.815 0.7 ;
        RECT 1.365 0.15 1.435 1.25 ;
        RECT 0.995 0.15 1.065 1.25 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.47 1.485 ;
        RECT 2.315 0.975 2.385 1.485 ;
        RECT 1.935 0.975 2.005 1.485 ;
        RECT 1.555 0.975 1.625 1.485 ;
        RECT 1.175 0.975 1.245 1.485 ;
        RECT 0.795 0.975 0.865 1.485 ;
        RECT 0.415 0.975 0.485 1.485 ;
        RECT 0.04 0.975 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.47 0.085 ;
        RECT 2.315 -0.085 2.385 0.425 ;
        RECT 1.935 -0.085 2.005 0.425 ;
        RECT 1.555 -0.085 1.625 0.425 ;
        RECT 1.185 -0.085 1.255 0.425 ;
        RECT 0.795 -0.085 0.865 0.425 ;
        RECT 0.415 -0.085 0.485 0.425 ;
        RECT 0.04 -0.085 0.11 0.425 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.605 0.15 0.675 1.25 ;
      RECT 0.235 0.15 0.305 1.25 ;
      RECT 0.235 0.525 0.925 0.66 ;
  END
END BUF_X8

MACRO CLKBUF_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUF_X1 0 0 ;
  SIZE 0.57 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.21 0.7 ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.15 0.51 1.24 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.57 1.485 ;
        RECT 0.245 0.965 0.315 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.57 0.085 ;
        RECT 0.245 -0.085 0.315 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.065 0.83 0.135 1.24 ;
      RECT 0.065 0.83 0.37 0.9 ;
      RECT 0.3 0.35 0.37 0.9 ;
      RECT 0.065 0.35 0.37 0.42 ;
      RECT 0.065 0.15 0.135 0.42 ;
  END
END CLKBUF_X1

MACRO CLKBUF_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUF_X2 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.19 0.7 ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425 0.15 0.51 1.25 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
        RECT 0.605 0.975 0.675 1.485 ;
        RECT 0.225 1.04 0.295 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
        RECT 0.605 -0.085 0.675 0.285 ;
        RECT 0.225 -0.085 0.295 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.905 0.115 1.25 ;
      RECT 0.045 0.905 0.36 0.975 ;
      RECT 0.29 0.35 0.36 0.975 ;
      RECT 0.045 0.35 0.36 0.42 ;
      RECT 0.045 0.15 0.115 0.42 ;
  END
END CLKBUF_X2

MACRO CLKBUF_X3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUF_X3 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.19 0.7 ;
    END
  END A
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.795 0.18 0.865 1.175 ;
        RECT 0.425 0.42 0.865 0.56 ;
        RECT 0.425 0.18 0.495 1.175 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.95 1.485 ;
        RECT 0.605 0.9 0.675 1.485 ;
        RECT 0.225 0.9 0.295 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.95 0.085 ;
        RECT 0.605 -0.085 0.675 0.235 ;
        RECT 0.225 -0.085 0.295 0.235 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.765 0.115 1.175 ;
      RECT 0.045 0.765 0.355 0.835 ;
      RECT 0.285 0.38 0.355 0.835 ;
      RECT 0.045 0.38 0.355 0.45 ;
      RECT 0.045 0.18 0.115 0.45 ;
  END
END CLKBUF_X3

MACRO CLKGATETST_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKGATETST_X1 0 0 ;
  SIZE 2.85 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.075 0.7 2.22 0.84 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.7 0.38 0.84 ;
    END
  END E
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.7 0.185 0.84 ;
    END
  END SE
  PIN GCK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.705 0.35 2.79 1.235 ;
    END
  END GCK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.85 1.485 ;
        RECT 2.48 1.045 2.615 1.485 ;
        RECT 2.135 0.94 2.205 1.485 ;
        RECT 1.755 0.94 1.825 1.485 ;
        RECT 1.185 1.01 1.32 1.485 ;
        RECT 0.385 1.04 0.52 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.85 0.085 ;
        RECT 2.485 -0.085 2.62 0.385 ;
        RECT 1.75 -0.085 1.82 0.42 ;
        RECT 1.185 -0.085 1.32 0.38 ;
        RECT 0.385 -0.085 0.52 0.385 ;
        RECT 0.04 -0.085 0.11 0.42 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 2.33 0.525 2.4 1.005 ;
      RECT 2.33 0.525 2.64 0.66 ;
      RECT 2.14 0.525 2.64 0.595 ;
      RECT 2.14 0.285 2.21 0.595 ;
      RECT 1.935 0.15 2.005 1.21 ;
      RECT 1.935 0.15 2.07 0.22 ;
      RECT 1.565 0.93 1.69 1.205 ;
      RECT 1.62 0.585 1.69 1.205 ;
      RECT 1.105 0.585 1.69 0.655 ;
      RECT 1.565 0.285 1.635 0.655 ;
      RECT 0.805 0.285 0.875 1.095 ;
      RECT 0.805 0.735 1.555 0.805 ;
      RECT 1.405 0.875 1.475 1.235 ;
      RECT 0.67 1.16 1.12 1.23 ;
      RECT 1.05 0.875 1.12 1.23 ;
      RECT 0.67 0.15 0.74 1.23 ;
      RECT 1.05 0.875 1.475 0.945 ;
      RECT 0.945 0.445 1.475 0.515 ;
      RECT 1.405 0.285 1.475 0.515 ;
      RECT 0.945 0.15 1.015 0.515 ;
      RECT 0.67 0.15 1.015 0.22 ;
      RECT 0.045 0.905 0.115 1.235 ;
      RECT 0.045 0.905 0.57 0.975 ;
      RECT 0.5 0.45 0.57 0.975 ;
      RECT 0.235 0.45 0.57 0.52 ;
      RECT 0.235 0.285 0.305 0.52 ;
  END
END CLKGATETST_X1

MACRO CLKGATETST_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKGATETST_X2 0 0 ;
  SIZE 3.04 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.18 0.85 2.825 0.92 ;
        RECT 2.72 0.525 2.825 0.92 ;
        RECT 2.18 0.525 2.25 0.92 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.56 0.375 0.725 ;
    END
  END E
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.56 0.545 0.725 ;
    END
  END SE
  PIN GCK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.52 0.15 2.6 0.785 ;
    END
  END GCK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 3.04 1.485 ;
        RECT 2.675 1.24 2.81 1.485 ;
        RECT 2.275 1.24 2.41 1.485 ;
        RECT 1.83 1.24 1.965 1.485 ;
        RECT 1.515 0.91 1.585 1.485 ;
        RECT 0.73 1.115 0.865 1.485 ;
        RECT 0.225 0.94 0.295 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 3.04 0.085 ;
        RECT 2.7 -0.085 2.77 0.195 ;
        RECT 2.325 -0.085 2.395 0.195 ;
        RECT 1.765 -0.085 1.9 0.185 ;
        RECT 1.45 -0.085 1.52 0.405 ;
        RECT 0.605 -0.085 0.675 0.285 ;
        RECT 0.225 -0.085 0.295 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.68 1.08 1.75 1.245 ;
      RECT 2.895 0.15 2.965 1.24 ;
      RECT 1.68 1.08 2.965 1.15 ;
      RECT 2.045 0.39 2.115 0.925 ;
      RECT 2.045 0.39 2.45 0.46 ;
      RECT 2.17 0.325 2.45 0.46 ;
      RECT 2.17 0.15 2.24 0.46 ;
      RECT 1.38 0.76 1.775 0.83 ;
      RECT 1.705 0.28 1.775 0.83 ;
      RECT 1.61 0.28 1.775 0.35 ;
      RECT 1.145 0.285 1.215 1.03 ;
      RECT 1.145 0.525 1.63 0.66 ;
      RECT 1.08 0.285 1.215 0.42 ;
      RECT 0.045 0.15 0.115 1.125 ;
      RECT 0.41 0.95 1.015 1.02 ;
      RECT 0.945 0.15 1.015 1.02 ;
      RECT 0.41 0.805 0.48 1.02 ;
      RECT 0.045 0.805 0.48 0.875 ;
      RECT 0.945 0.61 1.08 0.745 ;
      RECT 0.945 0.15 1.285 0.22 ;
      RECT 0.61 0.41 0.68 0.885 ;
      RECT 0.61 0.41 0.87 0.545 ;
      RECT 0.425 0.41 0.87 0.48 ;
      RECT 0.425 0.15 0.495 0.48 ;
  END
END CLKGATETST_X2

MACRO CLKGATETST_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKGATETST_X4 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.21 0.77 2.85 0.85 ;
        RECT 2.72 0.525 2.85 0.85 ;
        RECT 2.21 0.525 2.28 0.85 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.56 0.38 0.775 ;
    END
  END E
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.56 0.185 0.775 ;
    END
  END SE
  PIN GCK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.455 0.18 3.525 0.925 ;
        RECT 3.085 0.42 3.525 0.56 ;
        RECT 3.085 0.18 3.155 0.925 ;
    END
  END GCK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 3.8 1.485 ;
        RECT 3.645 0.975 3.715 1.485 ;
        RECT 3.265 0.975 3.335 1.485 ;
        RECT 2.885 1.2 2.955 1.485 ;
        RECT 2.505 1.2 2.575 1.485 ;
        RECT 2.13 1.205 2.2 1.485 ;
        RECT 1.49 1.165 1.625 1.485 ;
        RECT 0.755 1.13 0.825 1.485 ;
        RECT 0.415 0.975 0.485 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 3.8 0.085 ;
        RECT 3.645 -0.085 3.715 0.2 ;
        RECT 3.265 -0.085 3.335 0.2 ;
        RECT 2.885 -0.085 2.955 0.2 ;
        RECT 2.125 -0.085 2.195 0.285 ;
        RECT 1.53 -0.085 1.6 0.285 ;
        RECT 0.755 -0.085 0.825 0.195 ;
        RECT 0.415 -0.085 0.485 0.285 ;
        RECT 0.04 -0.085 0.11 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 2.29 0.93 3.015 1 ;
      RECT 2.945 0.35 3.015 1 ;
      RECT 2.655 0.35 3.015 0.42 ;
      RECT 2.655 0.185 2.725 0.42 ;
      RECT 2.48 0.185 2.725 0.255 ;
      RECT 1.13 1.03 1.205 1.25 ;
      RECT 1.13 1.03 2.125 1.1 ;
      RECT 2.055 0.39 2.125 1.1 ;
      RECT 1.13 0.525 1.2 1.25 ;
      RECT 2.425 0.39 2.495 0.66 ;
      RECT 1.13 0.525 1.645 0.66 ;
      RECT 1.39 0.185 1.46 0.66 ;
      RECT 2.055 0.39 2.495 0.46 ;
      RECT 1.11 0.185 1.46 0.255 ;
      RECT 1.265 0.865 1.99 0.935 ;
      RECT 1.92 0.15 1.99 0.935 ;
      RECT 1.265 0.795 1.335 0.935 ;
      RECT 1.405 0.725 1.78 0.795 ;
      RECT 1.71 0.15 1.78 0.795 ;
      RECT 0.575 0.975 0.645 1.25 ;
      RECT 0.575 0.975 1.065 1.045 ;
      RECT 0.975 0.39 1.065 1.045 ;
      RECT 0.975 0.39 1.325 0.46 ;
      RECT 0.975 0.26 1.045 1.045 ;
      RECT 0.575 0.26 1.045 0.33 ;
      RECT 0.575 0.15 0.645 0.33 ;
      RECT 0.045 0.84 0.115 1.25 ;
      RECT 0.045 0.84 0.91 0.91 ;
      RECT 0.84 0.415 0.91 0.91 ;
      RECT 0.235 0.415 0.91 0.485 ;
      RECT 0.235 0.15 0.335 0.485 ;
  END
END CLKGATETST_X4

MACRO CLKGATETST_X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKGATETST_X8 0 0 ;
  SIZE 5.51 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.385 0.845 3.925 0.915 ;
        RECT 3.855 0.56 3.925 0.915 ;
        RECT 3.765 0.56 3.925 0.63 ;
        RECT 3.1 0.56 3.17 0.915 ;
        RECT 3.035 0.56 3.17 0.63 ;
        RECT 2.385 0.525 2.455 0.915 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.33 0.7 0.51 0.84 ;
    END
  END E
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.7 0.25 0.84 ;
    END
  END SE
  PIN GCK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 5.205 0.15 5.275 1.25 ;
        RECT 4.12 0.56 5.275 0.7 ;
        RECT 4.825 0.15 4.895 1.25 ;
        RECT 4.445 0.15 4.515 1.25 ;
        RECT 4.075 0.975 4.19 1.25 ;
        RECT 4.12 0.15 4.19 1.25 ;
        RECT 4.075 0.15 4.19 0.285 ;
    END
  END GCK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 5.51 1.485 ;
        RECT 5.395 0.975 5.465 1.485 ;
        RECT 5.015 0.975 5.085 1.485 ;
        RECT 4.635 0.975 4.705 1.485 ;
        RECT 4.26 0.975 4.33 1.485 ;
        RECT 3.845 1.01 3.98 1.485 ;
        RECT 3.465 1.01 3.6 1.485 ;
        RECT 3.085 1.01 3.22 1.485 ;
        RECT 2.705 1.01 2.84 1.485 ;
        RECT 2.365 1.06 2.435 1.485 ;
        RECT 1.915 1.1 2.05 1.485 ;
        RECT 1.535 1.1 1.67 1.485 ;
        RECT 0.75 1.24 0.885 1.485 ;
        RECT 0.41 1.215 0.545 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 5.51 0.085 ;
        RECT 5.395 -0.085 5.465 0.285 ;
        RECT 5.015 -0.085 5.085 0.285 ;
        RECT 4.635 -0.085 4.705 0.285 ;
        RECT 4.255 -0.085 4.325 0.285 ;
        RECT 3.845 -0.085 3.98 0.25 ;
        RECT 3.085 -0.085 3.22 0.16 ;
        RECT 2.33 -0.085 2.465 0.16 ;
        RECT 1.95 -0.085 2.02 0.425 ;
        RECT 1.575 -0.085 1.645 0.265 ;
        RECT 0.75 -0.085 0.885 0.175 ;
        RECT 0.44 -0.085 0.51 0.285 ;
        RECT 0.065 -0.085 0.135 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 3.235 0.71 3.79 0.78 ;
      RECT 2.52 0.71 3.03 0.78 ;
      RECT 3.235 0.705 3.7 0.78 ;
      RECT 3.63 0.16 3.7 0.78 ;
      RECT 2.9 0.425 2.97 0.78 ;
      RECT 3.235 0.425 3.305 0.78 ;
      RECT 2.71 0.425 3.305 0.495 ;
      RECT 3.63 0.35 4.055 0.485 ;
      RECT 3.47 0.16 3.7 0.23 ;
      RECT 1.16 0.56 1.23 1.185 ;
      RECT 1.16 0.965 2.305 1.035 ;
      RECT 2.235 0.29 2.305 1.035 ;
      RECT 2.575 0.56 2.735 0.63 ;
      RECT 1.16 0.56 1.75 0.63 ;
      RECT 3.37 0.555 3.52 0.625 ;
      RECT 2.575 0.29 2.645 0.63 ;
      RECT 1.435 0.18 1.505 0.63 ;
      RECT 3.37 0.29 3.44 0.625 ;
      RECT 2.235 0.29 3.44 0.36 ;
      RECT 1.155 0.18 1.505 0.25 ;
      RECT 1.315 0.83 2.17 0.9 ;
      RECT 2.1 0.195 2.17 0.9 ;
      RECT 1.315 0.715 1.385 0.9 ;
      RECT 1.45 0.695 1.885 0.765 ;
      RECT 1.815 0.185 1.885 0.765 ;
      RECT 1.73 0.185 1.885 0.39 ;
      RECT 0.565 1.065 1.085 1.135 ;
      RECT 1.015 0.25 1.085 1.135 ;
      RECT 1.015 0.425 1.37 0.495 ;
      RECT 0.6 0.25 1.085 0.32 ;
      RECT 0.6 0.15 0.67 0.32 ;
      RECT 0.07 0.905 0.14 1.25 ;
      RECT 0.07 0.905 0.95 0.975 ;
      RECT 0.87 0.42 0.95 0.975 ;
      RECT 0.26 0.42 0.95 0.49 ;
      RECT 0.26 0.15 0.33 0.49 ;
  END
END CLKGATETST_X8

MACRO CLKGATE_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKGATE_X1 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.54 0.42 1.895 0.56 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.91 0.525 1.08 0.7 ;
    END
  END E
  PIN GCK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.31 0.175 2.41 1.09 ;
    END
  END GCK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.47 1.485 ;
        RECT 2.03 0.915 2.1 1.485 ;
        RECT 1.585 0.89 1.655 1.485 ;
        RECT 0.955 0.9 1.09 1.485 ;
        RECT 0.225 0.955 0.295 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.47 0.085 ;
        RECT 2.12 -0.085 2.19 0.225 ;
        RECT 1.585 -0.085 1.655 0.195 ;
        RECT 0.985 -0.085 1.055 0.32 ;
        RECT 0.225 -0.085 0.295 0.32 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.785 0.765 1.855 1.09 ;
      RECT 1.785 0.765 2.245 0.835 ;
      RECT 2.175 0.35 2.245 0.835 ;
      RECT 1.97 0.35 2.245 0.42 ;
      RECT 1.97 0.185 2.04 0.42 ;
      RECT 1.405 0.195 1.475 1.09 ;
      RECT 1.145 0.525 1.475 0.66 ;
      RECT 1.175 0.765 1.245 1.05 ;
      RECT 0.695 0.765 1.245 0.835 ;
      RECT 0.695 0.39 0.765 0.835 ;
      RECT 0.695 0.39 1.245 0.46 ;
      RECT 1.175 0.27 1.245 0.46 ;
      RECT 0.51 0.98 0.715 1.05 ;
      RECT 0.51 0.22 0.58 1.05 ;
      RECT 0.175 0.59 0.58 0.725 ;
      RECT 0.51 0.22 0.71 0.29 ;
      RECT 0.04 0.265 0.11 1.04 ;
      RECT 0.04 0.45 0.44 0.52 ;
  END
END CLKGATE_X1

MACRO CLKGATE_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKGATE_X2 0 0 ;
  SIZE 2.66 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.58 0.42 1.65 0.66 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.34 0.42 0.51 0.59 ;
    END
  END E
  PIN GCK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.32 0.185 2.41 1.215 ;
    END
  END GCK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.66 1.485 ;
        RECT 2.505 0.94 2.575 1.485 ;
        RECT 2.095 0.94 2.165 1.485 ;
        RECT 1.725 0.89 1.795 1.485 ;
        RECT 0.985 0.98 1.055 1.485 ;
        RECT 0.225 0.94 0.295 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.66 0.085 ;
        RECT 2.505 -0.085 2.575 0.22 ;
        RECT 2.095 -0.085 2.165 0.22 ;
        RECT 1.565 -0.085 1.635 0.235 ;
        RECT 0.955 -0.085 1.09 0.285 ;
        RECT 0.225 -0.085 0.295 0.32 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.915 0.805 1.985 1.215 ;
      RECT 1.915 0.805 2.255 0.875 ;
      RECT 2.185 0.39 2.255 0.875 ;
      RECT 1.725 0.39 2.255 0.46 ;
      RECT 1.725 0.185 1.795 0.46 ;
      RECT 1.12 1.18 1.64 1.25 ;
      RECT 1.57 0.755 1.64 1.25 ;
      RECT 0.36 1.18 0.92 1.25 ;
      RECT 0.85 0.79 0.92 1.25 ;
      RECT 1.12 0.79 1.19 1.25 ;
      RECT 0.36 0.805 0.43 1.25 ;
      RECT 0.04 0.295 0.11 1.17 ;
      RECT 0.04 0.805 0.43 0.875 ;
      RECT 0.85 0.79 1.19 0.86 ;
      RECT 1.57 0.755 1.785 0.825 ;
      RECT 1.715 0.56 1.785 0.825 ;
      RECT 1.715 0.56 2.095 0.63 ;
      RECT 1.42 0.49 1.49 0.975 ;
      RECT 1.065 0.49 1.49 0.56 ;
      RECT 1.385 0.185 1.455 0.56 ;
      RECT 1.255 0.65 1.325 1.115 ;
      RECT 0.74 0.65 1.325 0.72 ;
      RECT 0.74 0.585 0.99 0.72 ;
      RECT 0.92 0.35 0.99 0.72 ;
      RECT 0.92 0.35 1.28 0.42 ;
      RECT 0.605 0.2 0.675 1.115 ;
      RECT 0.175 0.655 0.675 0.725 ;
      RECT 0.175 0.525 0.245 0.725 ;
  END
END CLKGATE_X2

MACRO CLKGATE_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKGATE_X4 0 0 ;
  SIZE 3.23 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.895 0.39 1.965 0.66 ;
        RECT 1.535 0.39 1.965 0.46 ;
        RECT 1.535 0.39 1.65 0.7 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.35 0.42 0.51 0.63 ;
    END
  END E
  PIN GCK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.925 0.15 2.995 1.24 ;
        RECT 2.555 0.42 2.995 0.56 ;
        RECT 2.555 0.15 2.625 1.24 ;
    END
  END GCK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 3.23 1.485 ;
        RECT 3.115 0.965 3.185 1.485 ;
        RECT 2.735 0.965 2.805 1.485 ;
        RECT 2.355 1.065 2.425 1.485 ;
        RECT 1.975 1.065 2.045 1.485 ;
        RECT 1.57 1.24 1.705 1.485 ;
        RECT 0.995 0.965 1.065 1.485 ;
        RECT 0.235 0.965 0.305 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 3.23 0.085 ;
        RECT 3.115 -0.085 3.185 0.215 ;
        RECT 2.735 -0.085 2.805 0.215 ;
        RECT 2.325 -0.085 2.46 0.185 ;
        RECT 1.58 -0.085 1.65 0.285 ;
        RECT 0.995 -0.085 1.065 0.32 ;
        RECT 0.235 -0.085 0.305 0.32 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 2.165 0.905 2.235 1.24 ;
      RECT 1.79 0.905 1.86 1.24 ;
      RECT 1.79 0.905 2.49 0.975 ;
      RECT 2.42 0.255 2.49 0.975 ;
      RECT 1.95 0.255 2.49 0.325 ;
      RECT 0.05 0.15 0.12 1.24 ;
      RECT 0.37 1.165 0.885 1.235 ;
      RECT 0.815 0.83 0.885 1.235 ;
      RECT 1.13 1.105 1.64 1.175 ;
      RECT 1.57 0.765 1.64 1.175 ;
      RECT 0.37 0.83 0.44 1.235 ;
      RECT 1.13 0.83 1.2 1.175 ;
      RECT 0.815 0.83 1.2 0.9 ;
      RECT 0.05 0.83 0.44 0.9 ;
      RECT 1.57 0.765 2.32 0.835 ;
      RECT 2.25 0.525 2.32 0.835 ;
      RECT 0.92 0.56 0.99 0.9 ;
      RECT 1.715 0.525 1.785 0.835 ;
      RECT 1.4 0.15 1.47 1.04 ;
      RECT 1.19 0.56 1.47 0.63 ;
      RECT 1.265 0.695 1.335 0.87 ;
      RECT 1.055 0.695 1.335 0.765 ;
      RECT 1.055 0.39 1.125 0.765 ;
      RECT 0.75 0.39 0.82 0.66 ;
      RECT 0.75 0.39 1.255 0.46 ;
      RECT 1.185 0.3 1.255 0.46 ;
      RECT 0.615 0.2 0.685 1.095 ;
      RECT 0.185 0.695 0.685 0.765 ;
      RECT 0.185 0.525 0.255 0.765 ;
  END
END CLKGATE_X4

MACRO CLKGATE_X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKGATE_X8 0 0 ;
  SIZE 4.94 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.625 0.86 2.935 0.93 ;
        RECT 2.865 0.525 2.935 0.93 ;
        RECT 2.13 0.525 2.22 0.93 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.345 0.56 0.51 0.7 ;
    END
  END E
  PIN GCK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.615 0.15 4.685 1.235 ;
        RECT 3.485 0.42 4.685 0.56 ;
        RECT 4.235 0.15 4.305 1.235 ;
        RECT 3.855 0.15 3.925 1.235 ;
        RECT 3.485 0.15 3.555 1.235 ;
    END
  END GCK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 4.94 1.485 ;
        RECT 4.805 0.96 4.875 1.485 ;
        RECT 4.425 0.96 4.495 1.485 ;
        RECT 4.045 0.96 4.115 1.485 ;
        RECT 3.665 0.96 3.735 1.485 ;
        RECT 3.275 0.96 3.345 1.485 ;
        RECT 2.88 1.205 2.95 1.485 ;
        RECT 2.5 1.205 2.57 1.485 ;
        RECT 2.12 1.205 2.19 1.485 ;
        RECT 1.725 1.065 1.795 1.485 ;
        RECT 1.355 1.175 1.49 1.485 ;
        RECT 1.005 0.995 1.075 1.485 ;
        RECT 0.23 0.96 0.3 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 4.94 0.085 ;
        RECT 4.805 -0.085 4.875 0.285 ;
        RECT 4.425 -0.085 4.495 0.285 ;
        RECT 4.045 -0.085 4.115 0.285 ;
        RECT 3.67 -0.085 3.74 0.285 ;
        RECT 3.245 -0.085 3.38 0.16 ;
        RECT 2.47 -0.085 2.605 0.16 ;
        RECT 1.715 -0.085 1.85 0.16 ;
        RECT 1.355 -0.085 1.49 0.16 ;
        RECT 1.005 -0.085 1.075 0.285 ;
        RECT 0.2 -0.085 0.335 0.25 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 3.07 0.725 3.14 1.235 ;
      RECT 2.66 0.995 2.795 1.2 ;
      RECT 2.28 0.995 2.415 1.2 ;
      RECT 1.905 0.995 2.04 1.2 ;
      RECT 1.905 0.995 3.14 1.065 ;
      RECT 3.005 0.725 3.42 0.795 ;
      RECT 3.35 0.525 3.42 0.795 ;
      RECT 2.31 0.725 2.74 0.795 ;
      RECT 2.67 0.39 2.74 0.795 ;
      RECT 3.005 0.39 3.075 0.795 ;
      RECT 2.31 0.39 2.38 0.795 ;
      RECT 2.67 0.39 3.075 0.46 ;
      RECT 2.095 0.39 2.38 0.46 ;
      RECT 0.87 0.725 1.275 0.795 ;
      RECT 1.205 0.15 1.275 0.795 ;
      RECT 3.155 0.255 3.225 0.66 ;
      RECT 2.5 0.255 2.57 0.66 ;
      RECT 1.825 0.255 1.895 0.66 ;
      RECT 1.205 0.255 3.225 0.325 ;
      RECT 0.44 1.15 0.94 1.22 ;
      RECT 0.87 0.86 0.94 1.22 ;
      RECT 0.44 0.765 0.51 1.22 ;
      RECT 1.49 1.005 1.645 1.075 ;
      RECT 1.49 0.43 1.56 1.075 ;
      RECT 0.87 0.86 1.56 0.93 ;
      RECT 0.18 0.765 0.51 0.835 ;
      RECT 0.18 0.605 0.25 0.835 ;
      RECT 1.49 0.43 1.645 0.5 ;
      RECT 0.585 1.01 0.805 1.08 ;
      RECT 0.735 0.525 0.805 1.08 ;
      RECT 0.735 0.525 1.14 0.66 ;
      RECT 0.865 0.18 0.935 0.66 ;
      RECT 0.585 0.18 0.935 0.25 ;
      RECT 0.045 0.15 0.115 1.235 ;
      RECT 0.575 0.39 0.645 0.87 ;
      RECT 0.045 0.39 0.8 0.46 ;
  END
END CLKGATE_X8

MACRO DFFRS_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRS_X1 0 0 ;
  SIZE 4.56 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.12 0.585 4.31 0.84 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.2 0.7 1.345 0.84 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.8 0.7 0.89 0.84 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.24 0.28 4.385 0.495 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.4 0.51 0.875 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.185 0.13 1.075 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 4.56 1.485 ;
        RECT 4.255 0.915 4.325 1.485 ;
        RECT 3.325 1.03 3.46 1.485 ;
        RECT 2.795 0.835 2.93 1.485 ;
        RECT 2.415 0.89 2.55 1.485 ;
        RECT 1.655 0.99 1.79 1.485 ;
        RECT 1.345 0.925 1.415 1.485 ;
        RECT 0.965 1.065 1.035 1.485 ;
        RECT 0.56 1.095 0.695 1.485 ;
        RECT 0.215 1.1 0.35 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 4.56 0.085 ;
        RECT 4.225 -0.085 4.36 0.16 ;
        RECT 3.135 -0.085 3.27 0.285 ;
        RECT 2.415 -0.085 2.55 0.285 ;
        RECT 1.47 -0.085 1.605 0.285 ;
        RECT 0.935 -0.085 1.07 0.285 ;
        RECT 0.215 -0.085 0.35 0.2 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 3.68 1.18 4.055 1.25 ;
      RECT 3.985 0.15 4.055 1.25 ;
      RECT 1.955 1.165 2.275 1.235 ;
      RECT 2.205 0.35 2.275 1.235 ;
      RECT 3.68 0.76 3.75 1.25 ;
      RECT 3.02 0.76 3.09 1.07 ;
      RECT 3.02 0.76 3.75 0.83 ;
      RECT 3.62 0.15 3.69 0.46 ;
      RECT 2.98 0.35 3.69 0.42 ;
      RECT 2.205 0.35 2.76 0.42 ;
      RECT 2.69 0.165 2.76 0.42 ;
      RECT 2.98 0.165 3.05 0.42 ;
      RECT 2.69 0.165 3.05 0.235 ;
      RECT 3.62 0.15 4.055 0.22 ;
      RECT 3.85 0.62 3.92 1.115 ;
      RECT 2.5 0.62 3.92 0.69 ;
      RECT 3.76 0.285 3.83 0.69 ;
      RECT 3.545 0.895 3.615 1.115 ;
      RECT 3.175 0.895 3.245 1.115 ;
      RECT 3.175 0.895 3.615 0.965 ;
      RECT 2.635 0.755 2.705 1.07 ;
      RECT 2.345 0.755 2.705 0.825 ;
      RECT 2.345 0.485 2.415 0.825 ;
      RECT 2.345 0.485 3.545 0.555 ;
      RECT 2.825 0.3 2.895 0.555 ;
      RECT 2.065 0.185 2.135 1.085 ;
      RECT 1.09 0.495 2.135 0.63 ;
      RECT 1.875 0.855 1.945 1.075 ;
      RECT 1.505 0.855 1.575 1.075 ;
      RECT 1.505 0.855 1.945 0.925 ;
      RECT 0.955 0.925 1.26 0.995 ;
      RECT 0.955 0.35 1.025 0.995 ;
      RECT 0.595 0.555 1.025 0.625 ;
      RECT 0.95 0.35 1.025 0.625 ;
      RECT 0.95 0.35 1.9 0.425 ;
      RECT 0.2 0.96 0.88 1.03 ;
      RECT 0.2 0.265 0.27 1.03 ;
      RECT 0.2 0.265 0.695 0.335 ;
      RECT 4.45 0.185 4.52 1.25 ;
  END
END DFFRS_X1

MACRO DFFRS_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRS_X2 0 0 ;
  SIZE 4.94 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.485 0.28 4.69 0.46 ;
        RECT 4.485 0.28 4.555 0.575 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.39 0.545 1.46 0.7 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.2 0.545 1.27 0.7 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.62 0.54 4.72 0.7 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.625 0.4 0.7 0.965 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.24 0.2 0.32 0.965 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 4.94 1.485 ;
        RECT 4.59 0.765 4.66 1.485 ;
        RECT 3.695 1.03 3.83 1.485 ;
        RECT 3.195 0.765 3.265 1.485 ;
        RECT 2.815 0.955 2.885 1.485 ;
        RECT 2.055 0.955 2.125 1.485 ;
        RECT 1.715 0.895 1.785 1.485 ;
        RECT 1.335 1.08 1.405 1.485 ;
        RECT 0.875 1.205 0.945 1.485 ;
        RECT 0.425 1.205 0.495 1.485 ;
        RECT 0.05 0.925 0.12 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 4.94 0.085 ;
        RECT 4.56 -0.085 4.695 0.215 ;
        RECT 3.505 -0.085 3.64 0.285 ;
        RECT 2.785 -0.085 2.92 0.285 ;
        RECT 1.87 -0.085 1.94 0.32 ;
        RECT 1.335 -0.085 1.405 0.32 ;
        RECT 0.805 -0.085 0.875 0.2 ;
        RECT 0.425 -0.085 0.495 0.2 ;
        RECT 0.05 -0.085 0.12 0.415 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 4.05 1.18 4.39 1.25 ;
      RECT 4.32 0.15 4.39 1.25 ;
      RECT 2.325 1.14 2.64 1.21 ;
      RECT 2.57 0.35 2.64 1.21 ;
      RECT 4.05 0.76 4.12 1.25 ;
      RECT 3.39 0.76 3.46 1.04 ;
      RECT 3.39 0.76 4.12 0.83 ;
      RECT 3.985 0.15 4.055 0.46 ;
      RECT 3.35 0.35 4.055 0.42 ;
      RECT 2.57 0.35 3.13 0.42 ;
      RECT 3.06 0.185 3.13 0.42 ;
      RECT 3.35 0.185 3.42 0.42 ;
      RECT 3.06 0.185 3.42 0.255 ;
      RECT 3.985 0.15 4.39 0.22 ;
      RECT 4.185 0.62 4.255 1.115 ;
      RECT 2.895 0.62 4.255 0.69 ;
      RECT 4.13 0.285 4.2 0.69 ;
      RECT 3.915 0.895 3.985 1.115 ;
      RECT 3.545 0.895 3.615 1.115 ;
      RECT 3.545 0.895 3.985 0.965 ;
      RECT 3.005 0.755 3.075 1.04 ;
      RECT 2.76 0.755 3.075 0.825 ;
      RECT 2.76 0.485 2.83 0.825 ;
      RECT 2.76 0.485 3.915 0.555 ;
      RECT 3.195 0.32 3.265 0.555 ;
      RECT 2.425 0.2 2.505 1.075 ;
      RECT 1.58 0.58 2.505 0.65 ;
      RECT 2.245 0.82 2.315 1.075 ;
      RECT 1.875 0.82 1.945 1.075 ;
      RECT 1.875 0.82 2.315 0.89 ;
      RECT 1.065 0.845 1.63 0.915 ;
      RECT 1.065 0.41 1.135 0.915 ;
      RECT 0.84 0.525 1.135 0.66 ;
      RECT 1.065 0.41 2.27 0.48 ;
      RECT 1.715 0.205 1.785 0.48 ;
      RECT 0.49 1.035 1.225 1.105 ;
      RECT 0.49 0.265 0.56 1.105 ;
      RECT 0.385 0.525 0.56 0.66 ;
      RECT 0.49 0.265 1.065 0.335 ;
      RECT 4.785 0.25 4.855 1.24 ;
  END
END DFFRS_X2

MACRO DFFR_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFR_X1 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6 0.56 0.72 0.745 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.455 0.64 2.89 0.71 ;
        RECT 2.455 0.56 2.6 0.71 ;
        RECT 2.105 1.18 2.525 1.25 ;
        RECT 2.455 0.56 2.525 1.25 ;
        RECT 2.105 0.93 2.175 1.25 ;
        RECT 1.815 0.93 2.175 1 ;
        RECT 1.495 1.165 1.885 1.235 ;
        RECT 1.815 0.93 1.885 1.235 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.175 0.42 0.32 0.56 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.66 0.185 3.74 1.25 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.285 0.4 3.36 1.25 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 3.8 1.485 ;
        RECT 3.465 0.975 3.535 1.485 ;
        RECT 3.08 1.065 3.15 1.485 ;
        RECT 2.7 0.98 2.77 1.485 ;
        RECT 1.95 1.065 2.02 1.485 ;
        RECT 1.295 1.03 1.43 1.485 ;
        RECT 0.575 1.015 0.645 1.485 ;
        RECT 0.23 1.065 0.3 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 3.8 0.085 ;
        RECT 3.465 -0.085 3.535 0.195 ;
        RECT 2.7 -0.085 2.77 0.32 ;
        RECT 1.895 -0.085 2.03 0.285 ;
        RECT 1.515 -0.085 1.585 0.41 ;
        RECT 0.575 -0.085 0.645 0.32 ;
        RECT 0.23 -0.085 0.3 0.32 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 2.89 0.81 2.96 1.25 ;
      RECT 2.59 0.81 3.185 0.88 ;
      RECT 3.115 0.265 3.185 0.88 ;
      RECT 3.525 0.265 3.595 0.66 ;
      RECT 3.05 0.265 3.595 0.335 ;
      RECT 2.32 0.185 2.39 1.115 ;
      RECT 2.98 0.425 3.05 0.66 ;
      RECT 2.32 0.425 3.05 0.495 ;
      RECT 1.68 0.76 1.75 0.96 ;
      RECT 1.19 0.76 2.255 0.83 ;
      RECT 2.185 0.35 2.255 0.83 ;
      RECT 1.69 0.35 2.255 0.42 ;
      RECT 1.69 0.185 1.76 0.42 ;
      RECT 0.42 0.185 0.49 1.25 ;
      RECT 0.82 0.15 0.89 0.785 ;
      RECT 1.985 0.485 2.12 0.67 ;
      RECT 1.09 0.485 2.12 0.555 ;
      RECT 0.42 0.425 0.89 0.495 ;
      RECT 1.09 0.15 1.16 0.555 ;
      RECT 0.82 0.15 1.16 0.22 ;
      RECT 0.955 0.29 1.025 1.125 ;
      RECT 0.955 0.625 1.895 0.695 ;
      RECT 1.135 0.895 1.205 1.125 ;
      RECT 1.495 1.025 1.63 1.095 ;
      RECT 1.495 0.895 1.565 1.095 ;
      RECT 1.135 0.895 1.565 0.965 ;
      RECT 0.04 0.185 0.11 1.25 ;
      RECT 0.04 0.7 0.355 0.835 ;
  END
END DFFR_X1

MACRO DFFR_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFR_X2 0 0 ;
  SIZE 4.18 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.52 0.74 0.7 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.52 0.56 2.905 0.7 ;
        RECT 2.17 1.15 2.59 1.22 ;
        RECT 2.52 0.56 2.59 1.22 ;
        RECT 2.17 0.965 2.24 1.22 ;
        RECT 1.835 0.965 2.24 1.035 ;
        RECT 1.515 1.165 1.905 1.235 ;
        RECT 1.835 0.965 1.905 1.235 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.195 0.42 0.32 0.56 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.86 0.185 3.935 1.08 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.41 0.645 3.55 0.785 ;
        RECT 3.48 0.185 3.55 0.785 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 4.18 1.485 ;
        RECT 4.05 1.065 4.12 1.485 ;
        RECT 3.67 1.065 3.74 1.485 ;
        RECT 3.19 1.065 3.26 1.485 ;
        RECT 2.725 1 2.86 1.485 ;
        RECT 1.97 1.1 2.105 1.485 ;
        RECT 1.315 1.03 1.45 1.485 ;
        RECT 0.59 1.015 0.66 1.485 ;
        RECT 0.245 0.945 0.315 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 4.18 0.085 ;
        RECT 4.05 -0.085 4.12 0.335 ;
        RECT 3.67 -0.085 3.74 0.335 ;
        RECT 3.295 -0.085 3.365 0.195 ;
        RECT 2.69 -0.085 2.76 0.32 ;
        RECT 1.9 -0.085 2.035 0.285 ;
        RECT 1.535 -0.085 1.605 0.41 ;
        RECT 0.59 -0.085 0.66 0.32 ;
        RECT 0.245 -0.085 0.315 0.32 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 2.97 0.85 3.04 1.22 ;
      RECT 2.655 0.85 3.79 0.92 ;
      RECT 3.72 0.525 3.79 0.92 ;
      RECT 3.07 0.4 3.14 0.92 ;
      RECT 2.655 0.765 2.725 0.92 ;
      RECT 2.375 0.215 2.445 1.085 ;
      RECT 3.24 0.265 3.31 0.66 ;
      RECT 2.375 0.385 2.95 0.455 ;
      RECT 2.88 0.265 2.95 0.455 ;
      RECT 2.88 0.265 3.31 0.335 ;
      RECT 2.285 0.215 2.445 0.285 ;
      RECT 1.7 0.76 1.77 0.96 ;
      RECT 1.7 0.83 2.26 0.9 ;
      RECT 2.19 0.35 2.26 0.9 ;
      RECT 1.235 0.76 1.77 0.83 ;
      RECT 1.75 0.35 2.26 0.42 ;
      RECT 1.75 0.185 1.82 0.42 ;
      RECT 0.44 0.185 0.51 0.98 ;
      RECT 0.83 0.15 0.9 0.82 ;
      RECT 2.055 0.485 2.125 0.705 ;
      RECT 1.105 0.485 2.125 0.555 ;
      RECT 1.105 0.15 1.175 0.555 ;
      RECT 0.44 0.385 0.9 0.455 ;
      RECT 0.83 0.15 1.175 0.22 ;
      RECT 0.97 0.29 1.04 1.125 ;
      RECT 1.85 0.625 1.925 0.765 ;
      RECT 0.97 0.625 1.925 0.695 ;
      RECT 1.155 0.895 1.225 1.125 ;
      RECT 1.515 1.025 1.65 1.095 ;
      RECT 1.515 0.895 1.585 1.095 ;
      RECT 1.155 0.895 1.585 0.965 ;
      RECT 0.06 0.185 0.13 1.22 ;
      RECT 0.06 0.655 0.375 0.79 ;
  END
END DFFR_X2

MACRO DFFS_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFS_X1 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.34 0.56 0.51 0.7 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.625 0.7 2.79 0.84 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.77 0.59 1.84 0.84 ;
        RECT 1.705 0.59 1.84 0.725 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.575 0.56 3.74 0.7 ;
        RECT 3.575 0.185 3.645 1.16 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.195 0.56 3.36 0.7 ;
        RECT 3.195 0.185 3.265 0.925 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 3.8 1.485 ;
        RECT 3.38 1.205 3.45 1.485 ;
        RECT 2.855 1.005 2.925 1.485 ;
        RECT 2.48 1.065 2.615 1.485 ;
        RECT 1.755 0.905 1.825 1.485 ;
        RECT 1.41 0.885 1.48 1.485 ;
        RECT 1.015 0.94 1.085 1.485 ;
        RECT 0.225 0.9 0.295 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 3.8 0.085 ;
        RECT 3.385 -0.085 3.455 0.46 ;
        RECT 2.67 -0.085 2.805 0.34 ;
        RECT 1.75 -0.085 1.82 0.375 ;
        RECT 1.04 -0.085 1.11 0.32 ;
        RECT 0.225 -0.085 0.295 0.32 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 3.01 0.995 3.505 1.065 ;
      RECT 3.435 0.525 3.505 1.065 ;
      RECT 3.01 0.42 3.08 1.065 ;
      RECT 2.375 0.42 3.08 0.49 ;
      RECT 2.905 0.185 2.975 0.49 ;
      RECT 2.105 1.045 2.24 1.115 ;
      RECT 2.17 0.29 2.24 1.115 ;
      RECT 2.17 0.56 2.925 0.63 ;
      RECT 2.105 0.29 2.24 0.36 ;
      RECT 2.7 0.93 2.77 1.15 ;
      RECT 2.33 0.93 2.4 1.15 ;
      RECT 2.33 0.93 2.77 1 ;
      RECT 1.57 0.815 1.67 1.09 ;
      RECT 0.635 0.72 0.73 0.855 ;
      RECT 1.57 0.15 1.64 1.09 ;
      RECT 1.97 0.665 2.095 0.8 ;
      RECT 0.635 0.42 0.705 0.855 ;
      RECT 0.175 0.42 0.245 0.685 ;
      RECT 1.97 0.15 2.04 0.8 ;
      RECT 1.57 0.44 2.04 0.51 ;
      RECT 0.175 0.42 0.705 0.49 ;
      RECT 0.905 0.385 1.35 0.455 ;
      RECT 1.28 0.15 1.35 0.455 ;
      RECT 0.445 0.15 0.515 0.49 ;
      RECT 0.905 0.15 0.975 0.455 ;
      RECT 1.97 0.15 2.32 0.22 ;
      RECT 1.28 0.15 1.64 0.22 ;
      RECT 0.445 0.15 0.975 0.22 ;
      RECT 1.22 0.75 1.29 1.09 ;
      RECT 0.94 0.75 1.485 0.82 ;
      RECT 1.415 0.285 1.485 0.82 ;
      RECT 0.94 0.685 1.01 0.82 ;
      RECT 0.59 0.975 0.865 1.045 ;
      RECT 0.795 0.545 0.865 1.045 ;
      RECT 1.28 0.545 1.35 0.685 ;
      RECT 0.77 0.545 1.35 0.615 ;
      RECT 0.77 0.285 0.84 0.615 ;
      RECT 0.59 0.285 0.84 0.355 ;
      RECT 0.04 0.185 0.11 1.16 ;
      RECT 0.04 0.765 0.57 0.835 ;
  END
END DFFS_X1

MACRO DFFS_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFS_X2 0 0 ;
  SIZE 3.99 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.35 0.56 0.51 0.7 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.675 0.56 2.79 0.7 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.75 0.59 1.84 0.84 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.1 0.4 3.17 0.925 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.48 0.4 3.55 0.925 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 3.99 1.485 ;
        RECT 3.66 1.205 3.73 1.485 ;
        RECT 3.285 1.205 3.355 1.485 ;
        RECT 2.91 1.205 2.98 1.485 ;
        RECT 2.53 1.065 2.665 1.485 ;
        RECT 1.805 0.94 1.875 1.485 ;
        RECT 1.46 0.94 1.53 1.485 ;
        RECT 1.08 0.94 1.15 1.485 ;
        RECT 0.235 0.94 0.305 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 3.99 0.085 ;
        RECT 3.66 -0.085 3.73 0.195 ;
        RECT 3.28 -0.085 3.35 0.195 ;
        RECT 2.72 -0.085 2.855 0.34 ;
        RECT 1.8 -0.085 1.87 0.32 ;
        RECT 1.09 -0.085 1.16 0.37 ;
        RECT 0.235 -0.085 0.305 0.32 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 3.85 0.26 3.92 1.215 ;
      RECT 2.92 0.99 3.92 1.06 ;
      RECT 3.235 0.525 3.305 1.06 ;
      RECT 2.92 0.795 2.99 1.06 ;
      RECT 2.45 0.795 2.99 0.865 ;
      RECT 2.155 1.045 2.29 1.115 ;
      RECT 2.22 0.29 2.29 1.115 ;
      RECT 3.615 0.265 3.685 0.66 ;
      RECT 2.22 0.405 3.035 0.475 ;
      RECT 2.965 0.265 3.035 0.475 ;
      RECT 2.155 0.29 2.29 0.36 ;
      RECT 2.965 0.265 3.685 0.335 ;
      RECT 2.75 0.93 2.82 1.15 ;
      RECT 2.38 0.93 2.45 1.15 ;
      RECT 2.38 0.93 2.82 1 ;
      RECT 1.615 0.94 1.72 1.075 ;
      RECT 1.615 0.15 1.685 1.075 ;
      RECT 0.65 0.735 0.755 0.87 ;
      RECT 2.02 0.665 2.145 0.8 ;
      RECT 0.65 0.425 0.72 0.87 ;
      RECT 0.19 0.425 0.26 0.695 ;
      RECT 2.02 0.15 2.09 0.8 ;
      RECT 1.615 0.455 2.09 0.525 ;
      RECT 0.955 0.435 1.295 0.505 ;
      RECT 1.225 0.15 1.295 0.505 ;
      RECT 0.19 0.425 0.72 0.495 ;
      RECT 0.955 0.15 1.025 0.505 ;
      RECT 0.455 0.15 0.525 0.495 ;
      RECT 2.02 0.15 2.395 0.22 ;
      RECT 1.225 0.15 1.685 0.22 ;
      RECT 0.455 0.15 1.025 0.22 ;
      RECT 0.965 0.77 1.535 0.84 ;
      RECT 1.465 0.285 1.535 0.84 ;
      RECT 0.585 0.975 0.89 1.045 ;
      RECT 0.82 0.285 0.89 1.045 ;
      RECT 0.82 0.57 1.4 0.705 ;
      RECT 0.59 0.285 0.89 0.355 ;
      RECT 0.05 0.185 0.12 1.215 ;
      RECT 0.05 0.765 0.585 0.835 ;
  END
END DFFS_X2

MACRO DFF_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFF_X1 0 0 ;
  SIZE 3.23 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.81 0.53 0.97 0.7 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.56 0.53 1.67 0.7 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.1 0.26 3.17 1.13 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.72 0.26 2.79 0.785 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 3.23 1.485 ;
        RECT 2.905 0.985 2.975 1.485 ;
        RECT 2.345 1.1 2.48 1.485 ;
        RECT 1.61 0.9 1.68 1.485 ;
        RECT 1.005 1.08 1.075 1.485 ;
        RECT 0.24 0.98 0.31 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 3.23 0.085 ;
        RECT 2.905 -0.085 2.975 0.46 ;
        RECT 2.345 -0.085 2.48 0.37 ;
        RECT 1.61 -0.085 1.68 0.36 ;
        RECT 0.975 -0.085 1.11 0.3 ;
        RECT 0.24 -0.085 0.31 0.405 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 2.57 0.225 2.64 1.115 ;
      RECT 2.57 0.85 3.035 0.92 ;
      RECT 2.965 0.525 3.035 0.92 ;
      RECT 2.265 0.73 2.64 0.8 ;
      RECT 2 0.285 2.07 1.2 ;
      RECT 2 0.525 2.505 0.66 ;
      RECT 1.14 1.18 1.495 1.25 ;
      RECT 1.425 0.225 1.495 1.25 ;
      RECT 0.485 1.18 0.94 1.25 ;
      RECT 0.87 0.945 0.94 1.25 ;
      RECT 1.14 0.945 1.21 1.25 ;
      RECT 0.87 0.945 1.21 1.015 ;
      RECT 1.425 0.765 1.925 0.835 ;
      RECT 1.855 0.15 1.925 0.835 ;
      RECT 1.855 0.15 2.205 0.22 ;
      RECT 1.275 0.37 1.345 0.995 ;
      RECT 0.38 0.15 0.45 0.545 ;
      RECT 0.785 0.37 1.345 0.44 ;
      RECT 1.2 0.27 1.27 0.44 ;
      RECT 0.785 0.15 0.855 0.44 ;
      RECT 0.38 0.15 0.855 0.22 ;
      RECT 0.635 0.285 0.705 1.115 ;
      RECT 0.635 0.765 1.19 0.835 ;
      RECT 1.12 0.53 1.19 0.835 ;
      RECT 0.06 0.27 0.13 1.13 ;
      RECT 0.06 0.61 0.57 0.745 ;
  END
END DFF_X1

MACRO DFF_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFF_X2 0 0 ;
  SIZE 3.61 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.94 0.56 1.08 0.7 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.57 0.56 1.65 0.7 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.29 0.25 3.36 1.115 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.91 0.25 2.98 0.925 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 3.61 1.485 ;
        RECT 3.485 0.84 3.555 1.485 ;
        RECT 3.105 1.205 3.175 1.485 ;
        RECT 2.73 1.205 2.8 1.485 ;
        RECT 2.35 0.875 2.485 1.485 ;
        RECT 1.62 0.9 1.69 1.485 ;
        RECT 1.015 1.08 1.085 1.485 ;
        RECT 0.255 0.965 0.325 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 3.61 0.085 ;
        RECT 3.485 -0.085 3.555 0.46 ;
        RECT 3.105 -0.085 3.175 0.46 ;
        RECT 2.73 -0.085 2.8 0.46 ;
        RECT 2.35 -0.085 2.485 0.45 ;
        RECT 1.62 -0.085 1.69 0.385 ;
        RECT 0.985 -0.085 1.12 0.215 ;
        RECT 0.255 -0.085 0.325 0.385 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 2.575 1.045 3.215 1.115 ;
      RECT 3.145 0.525 3.215 1.115 ;
      RECT 2.575 0.2 2.645 1.115 ;
      RECT 2.245 0.735 2.645 0.805 ;
      RECT 2.01 0.35 2.08 0.975 ;
      RECT 2.01 0.525 2.51 0.66 ;
      RECT 1.15 1.18 1.505 1.25 ;
      RECT 1.435 0.25 1.505 1.25 ;
      RECT 0.5 1.18 0.935 1.25 ;
      RECT 0.865 0.945 0.935 1.25 ;
      RECT 1.15 0.945 1.22 1.25 ;
      RECT 0.865 0.945 1.22 1.015 ;
      RECT 1.435 0.765 1.945 0.835 ;
      RECT 1.875 0.215 1.945 0.835 ;
      RECT 1.875 0.215 2.215 0.285 ;
      RECT 1.285 0.285 1.355 1.115 ;
      RECT 0.39 0.15 0.46 0.7 ;
      RECT 0.825 0.285 1.355 0.355 ;
      RECT 0.825 0.15 0.895 0.355 ;
      RECT 0.39 0.15 0.895 0.22 ;
      RECT 0.61 1 0.76 1.07 ;
      RECT 0.69 0.285 0.76 1.07 ;
      RECT 0.69 0.765 1.215 0.835 ;
      RECT 1.145 0.565 1.215 0.835 ;
      RECT 0.61 0.285 0.76 0.355 ;
      RECT 0.075 0.325 0.145 1.055 ;
      RECT 0.075 0.765 0.625 0.835 ;
      RECT 0.555 0.565 0.625 0.835 ;
  END
END DFF_X2

MACRO DLH_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLH_X1 0 0 ;
  SIZE 1.9 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.95 0.525 1.08 0.7 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 0.525 0.32 0.7 ;
    END
  END G
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.185 0.51 0.785 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.9 1.485 ;
        RECT 1.595 1.025 1.665 1.485 ;
        RECT 0.845 0.965 0.915 1.485 ;
        RECT 0.25 0.985 0.32 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.9 0.085 ;
        RECT 1.595 -0.085 1.665 0.445 ;
        RECT 0.805 -0.085 0.94 0.285 ;
        RECT 0.25 -0.085 0.32 0.32 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.79 0.32 1.86 1.16 ;
      RECT 1.485 0.525 1.86 0.595 ;
      RECT 1.19 1.045 1.415 1.115 ;
      RECT 1.345 0.35 1.415 1.115 ;
      RECT 1.345 0.66 1.725 0.795 ;
      RECT 0.785 0.35 0.855 0.66 ;
      RECT 0.785 0.35 1.415 0.42 ;
      RECT 1.025 1.18 1.43 1.25 ;
      RECT 1.025 0.765 1.095 1.25 ;
      RECT 0.65 0.185 0.72 1.115 ;
      RECT 0.65 0.765 1.215 0.835 ;
      RECT 1.145 0.49 1.215 0.835 ;
      RECT 1.145 0.49 1.28 0.56 ;
      RECT 0.505 1.18 0.78 1.25 ;
      RECT 0.065 0.185 0.135 1.24 ;
      RECT 0.505 0.85 0.575 1.25 ;
      RECT 0.065 0.85 0.575 0.92 ;
  END
END DLH_X1

MACRO DLH_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLH_X2 0 0 ;
  SIZE 2.09 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.135 0.525 1.27 0.7 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.18 0.525 0.32 0.7 ;
    END
  END G
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.185 0.51 0.785 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.09 1.485 ;
        RECT 1.78 1.08 1.85 1.485 ;
        RECT 1.03 1.04 1.1 1.485 ;
        RECT 0.62 1 0.69 1.485 ;
        RECT 0.24 1.055 0.31 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.09 0.085 ;
        RECT 1.78 -0.085 1.85 0.32 ;
        RECT 1.03 -0.085 1.1 0.32 ;
        RECT 0.62 -0.085 0.69 0.255 ;
        RECT 0.24 -0.085 0.31 0.255 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.975 0.185 2.045 1.215 ;
      RECT 1.705 0.495 2.045 0.63 ;
      RECT 1.4 0.78 1.47 1.2 ;
      RECT 1.4 0.78 1.91 0.875 ;
      RECT 1.545 0.74 1.91 0.875 ;
      RECT 0.985 0.78 1.91 0.85 ;
      RECT 0.985 0.525 1.055 0.85 ;
      RECT 1.545 0.185 1.615 0.875 ;
      RECT 1.41 0.185 1.615 0.32 ;
      RECT 0.82 0.975 0.92 1.25 ;
      RECT 0.85 0.175 0.92 1.25 ;
      RECT 1.405 0.39 1.475 0.67 ;
      RECT 0.85 0.39 1.475 0.46 ;
      RECT 0.82 0.175 0.92 0.31 ;
      RECT 0.045 0.185 0.115 1.24 ;
      RECT 0.045 0.85 0.78 0.92 ;
      RECT 0.71 0.375 0.78 0.92 ;
  END
END DLH_X2

MACRO DLL_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLL_X1 0 0 ;
  SIZE 1.9 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.56 0.43 0.7 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.58 0.525 1.705 0.7 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.39 0.26 1.46 0.84 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.9 1.485 ;
        RECT 1.575 1.04 1.645 1.485 ;
        RECT 1.035 0.95 1.105 1.485 ;
        RECT 0.275 0.915 0.345 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.9 0.085 ;
        RECT 1.575 -0.085 1.645 0.235 ;
        RECT 1.035 -0.085 1.105 0.42 ;
        RECT 0.275 -0.085 0.345 0.415 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.235 1.18 1.51 1.25 ;
      RECT 1.44 0.905 1.51 1.25 ;
      RECT 1.77 0.195 1.84 1.24 ;
      RECT 1.44 0.905 1.84 0.975 ;
      RECT 1.23 0.285 1.3 1.085 ;
      RECT 0.9 0.775 1.3 0.845 ;
      RECT 0.665 0.285 0.735 1.085 ;
      RECT 0.665 0.525 1.165 0.66 ;
      RECT 0.53 0.15 0.6 1.25 ;
      RECT 0.095 0.28 0.165 1.085 ;
      RECT 0.095 0.78 0.6 0.85 ;
      RECT 0.53 0.15 0.845 0.22 ;
  END
END DLL_X1

MACRO DLL_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLL_X2 0 0 ;
  SIZE 2.09 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.51 0.38 0.7 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.77 0.525 1.89 0.7 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.58 0.26 1.65 1.005 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.09 1.485 ;
        RECT 1.76 1.205 1.83 1.485 ;
        RECT 1.385 1.205 1.455 1.485 ;
        RECT 0.985 0.875 1.055 1.485 ;
        RECT 0.225 0.9 0.295 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.09 0.085 ;
        RECT 1.76 -0.085 1.83 0.195 ;
        RECT 1.385 -0.085 1.455 0.395 ;
        RECT 0.985 -0.085 1.055 0.46 ;
        RECT 0.225 -0.085 0.295 0.37 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.185 1.07 1.32 1.25 ;
      RECT 1.955 0.195 2.025 1.24 ;
      RECT 1.185 1.07 2.025 1.14 ;
      RECT 1.19 0.325 1.26 1.005 ;
      RECT 0.85 0.73 1.26 0.8 ;
      RECT 0.615 0.335 0.685 1.015 ;
      RECT 0.615 0.525 1.125 0.66 ;
      RECT 0.045 0.3 0.115 1.145 ;
      RECT 0.045 0.765 0.55 0.835 ;
      RECT 0.48 0.195 0.55 0.835 ;
      RECT 0.48 0.195 0.82 0.265 ;
  END
END DLL_X2

MACRO FA_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FA_X1 0 0 ;
  SIZE 3.04 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.905 0.825 2.66 0.895 ;
        RECT 2.53 0.7 2.66 0.895 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.34 0.42 2.47 0.56 ;
        RECT 1.41 0.42 2.47 0.49 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.555 2.275 0.625 ;
        RECT 0.63 0.42 0.7 0.625 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.195 0.135 1.215 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.89 0.195 2.98 1.215 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 3.04 1.485 ;
        RECT 2.695 1.205 2.765 1.485 ;
        RECT 1.705 1.095 1.84 1.485 ;
        RECT 1.36 0.965 1.43 1.485 ;
        RECT 1.015 1.095 1.085 1.485 ;
        RECT 0.25 0.94 0.32 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 3.04 0.085 ;
        RECT 2.665 -0.085 2.8 0.16 ;
        RECT 1.705 -0.085 1.84 0.16 ;
        RECT 1.36 -0.085 1.43 0.195 ;
        RECT 1.025 -0.085 1.095 0.33 ;
        RECT 0.25 -0.085 0.32 0.33 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 2.13 0.96 2.2 1.24 ;
      RECT 2.13 0.96 2.82 1.03 ;
      RECT 2.75 0.225 2.82 1.03 ;
      RECT 2.1 0.225 2.82 0.295 ;
      RECT 0.63 0.69 0.7 1.215 ;
      RECT 0.495 0.69 2.115 0.76 ;
      RECT 0.495 0.23 0.565 0.76 ;
      RECT 0.205 0.525 0.565 0.66 ;
      RECT 0.495 0.23 0.735 0.3 ;
      RECT 1.93 0.96 2 1.24 ;
      RECT 1.555 0.96 1.625 1.24 ;
      RECT 1.555 0.96 2 1.03 ;
      RECT 0.835 0.395 1.275 0.465 ;
      RECT 1.205 0.195 1.275 0.465 ;
      RECT 0.835 0.195 0.905 0.465 ;
      RECT 1.205 0.96 1.275 1.235 ;
      RECT 0.8 0.96 0.935 1.215 ;
      RECT 0.8 0.96 1.275 1.03 ;
      RECT 1.52 0.225 2.03 0.295 ;
  END
END FA_X1

MACRO TAPCELL_X1
  #CLASS CORE ;
  CLASS CORE WELLTAP ;
  ORIGIN 0 0 ;
  FOREIGN TAPCELL_X1 0 0 ;
  SIZE 0.19 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.19 1.485 ;
        RECT 0.06 0.975 0.13 1.315 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.19 0.085 ;
        RECT 0.06 0.085 0.13 0.425 ;
    END
  END VSS
END TAPCELL_X1

MACRO FILLCELL_X1
  #CLASS CORE ;
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN FILLCELL_X1 0 0 ;
  SIZE 0.19 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.19 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.19 0.085 ;
    END
  END VSS
END FILLCELL_X1

MACRO FILLCELL_X16
  #CLASS CORE ;
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN FILLCELL_X16 0 0 ;
  SIZE 3.04 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 3.04 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 3.04 0.085 ;
    END
  END VSS
END FILLCELL_X16

MACRO FILLCELL_X2
  #CLASS CORE ;
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN FILLCELL_X2 0 0 ;
  SIZE 0.38 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.19 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.19 0.085 ;
    END
  END VSS
END FILLCELL_X2

MACRO FILLCELL_X32
  #CLASS CORE ;
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN FILLCELL_X32 0 0 ;
  SIZE 6.08 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 6.08 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 6.08 0.085 ;
    END
  END VSS
END FILLCELL_X32

MACRO FILLCELL_X4
  #CLASS CORE ;
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN FILLCELL_X4 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
    END
  END VSS
END FILLCELL_X4

MACRO FILLCELL_X8
  #CLASS CORE ;
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN FILLCELL_X8 0 0 ;
  SIZE 1.52 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.52 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.52 0.085 ;
    END
  END VSS
END FILLCELL_X8

MACRO HA_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HA_X1 0 0 ;
  SIZE 1.9 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.01 0.56 1.08 0.7 ;
        RECT 0.67 0.56 1.08 0.63 ;
        RECT 0.355 0.725 0.74 0.795 ;
        RECT 0.67 0.56 0.74 0.795 ;
        RECT 0.355 0.525 0.425 0.795 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.195 0.86 0.89 0.93 ;
        RECT 0.805 0.7 0.89 0.93 ;
        RECT 0.195 0.525 0.265 0.93 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.77 0.15 1.85 1.25 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.29 0.525 0.36 ;
        RECT 0.455 0.15 0.525 0.36 ;
        RECT 0.06 0.995 0.37 1.065 ;
        RECT 0.06 0.29 0.13 1.065 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.9 1.485 ;
        RECT 1.59 1.08 1.66 1.485 ;
        RECT 1.22 0.94 1.29 1.485 ;
        RECT 0.645 1.08 0.715 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.9 0.085 ;
        RECT 1.59 -0.085 1.66 0.285 ;
        RECT 1.03 -0.085 1.1 0.285 ;
        RECT 0.645 -0.085 0.715 0.285 ;
        RECT 0.08 -0.085 0.15 0.225 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.4 0.15 1.47 1.115 ;
      RECT 1.4 0.525 1.705 0.66 ;
      RECT 1.22 0.15 1.47 0.285 ;
      RECT 1.035 0.765 1.105 1.115 ;
      RECT 1.035 0.765 1.25 0.835 ;
      RECT 1.18 0.425 1.25 0.835 ;
      RECT 0.535 0.425 0.605 0.66 ;
      RECT 0.535 0.425 1.25 0.495 ;
      RECT 0.84 0.15 0.91 0.495 ;
      RECT 0.05 1.13 0.56 1.2 ;
  END
END HA_X1

MACRO INV_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X1 0 0 ;
  SIZE 0.38 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.165 0.7 ;
    END
  END A
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.23 0.15 0.325 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.38 1.485 ;
        RECT 0.04 0.975 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.38 0.085 ;
        RECT 0.04 -0.085 0.11 0.425 ;
    END
  END VSS
END INV_X1

MACRO INV_X16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X16 0 0 ;
  SIZE 3.23 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.095 1.05 3.095 1.12 ;
        RECT 3.025 0.525 3.095 1.12 ;
        RECT 2 0.525 2.07 1.12 ;
        RECT 1.2 0.525 1.27 1.12 ;
        RECT 0.095 0.525 0.165 1.12 ;
    END
  END A
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.885 0.15 2.955 0.985 ;
        RECT 0.235 0.28 2.955 0.42 ;
        RECT 2.505 0.15 2.575 0.985 ;
        RECT 2.135 0.28 2.205 0.985 ;
        RECT 2.125 0.15 2.195 0.42 ;
        RECT 1.745 0.15 1.815 0.985 ;
        RECT 1.365 0.15 1.435 0.985 ;
        RECT 0.985 0.15 1.055 0.985 ;
        RECT 0.605 0.16 0.675 0.985 ;
        RECT 0.235 0.18 0.305 0.985 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 3.23 1.485 ;
        RECT 3.075 1.205 3.145 1.485 ;
        RECT 2.695 1.205 2.765 1.485 ;
        RECT 2.315 1.205 2.385 1.485 ;
        RECT 1.935 1.205 2.005 1.485 ;
        RECT 1.555 1.205 1.625 1.485 ;
        RECT 1.175 1.205 1.245 1.485 ;
        RECT 0.795 1.205 0.865 1.485 ;
        RECT 0.415 1.205 0.485 1.485 ;
        RECT 0.04 1.205 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 3.23 0.085 ;
        RECT 3.075 -0.085 3.145 0.365 ;
        RECT 2.695 -0.085 2.765 0.21 ;
        RECT 2.315 -0.085 2.385 0.21 ;
        RECT 1.935 -0.085 2.005 0.21 ;
        RECT 1.555 -0.085 1.625 0.21 ;
        RECT 1.175 -0.085 1.245 0.21 ;
        RECT 0.795 -0.085 0.865 0.21 ;
        RECT 0.415 -0.085 0.485 0.21 ;
        RECT 0.04 -0.085 0.11 0.365 ;
    END
  END VSS
END INV_X16

MACRO INV_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X2 0 0 ;
  SIZE 0.57 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.15 0.32 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.57 1.485 ;
        RECT 0.43 0.975 0.5 1.485 ;
        RECT 0.055 0.975 0.125 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.57 0.085 ;
        RECT 0.43 -0.085 0.5 0.425 ;
        RECT 0.055 -0.085 0.125 0.425 ;
    END
  END VSS
END INV_X2

MACRO INV_X32
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X32 0 0 ;
  SIZE 6.27 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.115 0.93 5.85 1 ;
        RECT 5.78 0.525 5.85 1 ;
        RECT 4.62 0.525 4.69 1 ;
        RECT 3.48 0.525 3.55 1 ;
        RECT 2.34 0.525 2.41 1 ;
        RECT 1.2 0.525 1.27 1 ;
        RECT 0.115 0.525 0.185 1 ;
    END
  END A
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 5.945 0.16 6.015 1.005 ;
        RECT 0.25 0.28 6.015 0.42 ;
        RECT 5.56 0.16 5.63 0.865 ;
        RECT 5.18 0.16 5.25 0.865 ;
        RECT 4.81 0.28 4.88 0.865 ;
        RECT 4.8 0.16 4.87 0.42 ;
        RECT 4.42 0.16 4.49 0.865 ;
        RECT 4.04 0.16 4.11 0.865 ;
        RECT 3.665 0.16 3.735 0.865 ;
        RECT 3.28 0.16 3.35 0.865 ;
        RECT 2.9 0.16 2.97 0.865 ;
        RECT 2.525 0.16 2.595 0.865 ;
        RECT 2.14 0.16 2.21 0.865 ;
        RECT 1.76 0.16 1.83 0.865 ;
        RECT 1.39 0.16 1.46 0.865 ;
        RECT 1 0.16 1.07 0.865 ;
        RECT 0.62 0.16 0.69 0.865 ;
        RECT 0.25 0.16 0.32 0.865 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 6.27 1.485 ;
        RECT 6.13 1.065 6.2 1.485 ;
        RECT 5.75 1.065 5.82 1.485 ;
        RECT 5.37 1.065 5.44 1.485 ;
        RECT 4.99 1.065 5.06 1.485 ;
        RECT 4.61 1.065 4.68 1.485 ;
        RECT 4.23 1.065 4.3 1.485 ;
        RECT 3.85 1.065 3.92 1.485 ;
        RECT 3.47 1.065 3.54 1.485 ;
        RECT 3.09 1.065 3.16 1.485 ;
        RECT 2.71 1.065 2.78 1.485 ;
        RECT 2.33 1.065 2.4 1.485 ;
        RECT 1.95 1.065 2.02 1.485 ;
        RECT 1.57 1.065 1.64 1.485 ;
        RECT 1.19 1.065 1.26 1.485 ;
        RECT 0.81 1.065 0.88 1.485 ;
        RECT 0.43 1.065 0.5 1.485 ;
        RECT 0.055 1.065 0.125 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 6.27 0.085 ;
        RECT 6.13 -0.085 6.2 0.335 ;
        RECT 5.75 -0.085 5.82 0.195 ;
        RECT 5.37 -0.085 5.44 0.195 ;
        RECT 4.99 -0.085 5.06 0.195 ;
        RECT 4.61 -0.085 4.68 0.195 ;
        RECT 4.23 -0.085 4.3 0.195 ;
        RECT 3.85 -0.085 3.92 0.195 ;
        RECT 3.47 -0.085 3.54 0.195 ;
        RECT 3.09 -0.085 3.16 0.195 ;
        RECT 2.71 -0.085 2.78 0.195 ;
        RECT 2.33 -0.085 2.4 0.195 ;
        RECT 1.95 -0.085 2.02 0.195 ;
        RECT 1.57 -0.085 1.64 0.195 ;
        RECT 1.19 -0.085 1.26 0.195 ;
        RECT 0.81 -0.085 0.88 0.195 ;
        RECT 0.43 -0.085 0.5 0.195 ;
        RECT 0.055 -0.085 0.125 0.335 ;
    END
  END VSS
END INV_X32

MACRO INV_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X4 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.17 0.7 ;
    END
  END A
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.615 0.15 0.685 1.04 ;
        RECT 0.235 0.56 0.685 0.7 ;
        RECT 0.61 0.15 0.685 0.7 ;
        RECT 0.235 0.15 0.305 1.04 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.95 1.485 ;
        RECT 0.795 0.98 0.865 1.485 ;
        RECT 0.415 0.98 0.485 1.485 ;
        RECT 0.04 0.98 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.95 0.085 ;
        RECT 0.795 -0.085 0.865 0.425 ;
        RECT 0.415 -0.085 0.485 0.425 ;
        RECT 0.04 -0.085 0.11 0.425 ;
    END
  END VSS
END INV_X4

MACRO INV_X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X8 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.17 0.7 ;
    END
  END A
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.375 0.15 1.445 1.04 ;
        RECT 0.235 0.56 1.445 0.7 ;
        RECT 0.985 0.15 1.055 1.04 ;
        RECT 0.605 0.15 0.675 1.04 ;
        RECT 0.235 0.15 0.305 1.04 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.71 1.485 ;
        RECT 1.555 0.97 1.625 1.485 ;
        RECT 1.175 0.97 1.245 1.485 ;
        RECT 0.795 0.97 0.865 1.485 ;
        RECT 0.415 0.97 0.485 1.485 ;
        RECT 0.04 0.97 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.71 0.085 ;
        RECT 1.555 -0.085 1.625 0.36 ;
        RECT 1.175 -0.085 1.245 0.36 ;
        RECT 0.795 -0.085 0.865 0.36 ;
        RECT 0.415 -0.085 0.485 0.36 ;
        RECT 0.04 -0.085 0.11 0.36 ;
    END
  END VSS
END INV_X8

MACRO LOGIC0_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LOGIC0_X1 0 0 ;
  SIZE 0.38 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.15 0.13 0.84 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.38 1.485 ;
        RECT 0.245 1.115 0.315 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.38 0.085 ;
        RECT 0.24 -0.085 0.31 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.06 0.975 0.18 1.25 ;
  END
END LOGIC0_X1

MACRO LOGIC1_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LOGIC1_X1 0 0 ;
  SIZE 0.38 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.56 0.13 1.25 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.38 1.485 ;
        RECT 0.24 1.115 0.31 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.38 0.085 ;
        RECT 0.245 -0.085 0.315 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.06 0.15 0.18 0.425 ;
  END
END LOGIC1_X1

MACRO MUX2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2_X1 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.38 0.7 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.82 0.525 0.95 0.7 ;
    END
  END B
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.765 0.595 0.835 ;
        RECT 0.525 0.535 0.595 0.835 ;
        RECT 0.06 0.525 0.185 0.835 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.18 0.19 1.27 1.23 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.33 1.485 ;
        RECT 0.985 0.975 1.055 1.485 ;
        RECT 0.225 1.035 0.295 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.33 0.085 ;
        RECT 0.985 -0.085 1.055 0.24 ;
        RECT 0.225 -0.085 0.295 0.24 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.58 1.07 0.92 1.14 ;
      RECT 0.85 0.84 0.92 1.14 ;
      RECT 0.85 0.84 1.115 0.91 ;
      RECT 1.045 0.39 1.115 0.91 ;
      RECT 0.83 0.39 1.115 0.46 ;
      RECT 0.83 0.22 0.9 0.46 ;
      RECT 0.58 0.22 0.9 0.29 ;
      RECT 0.045 0.9 0.115 1.25 ;
      RECT 0.045 0.9 0.755 0.97 ;
      RECT 0.685 0.39 0.755 0.97 ;
      RECT 0.045 0.39 0.755 0.46 ;
      RECT 0.045 0.19 0.115 0.46 ;
  END
END MUX2_X1

MACRO MUX2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2_X2 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.225 0.7 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.575 0.525 0.7 0.7 ;
    END
  END B
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.925 0.85 1.535 0.92 ;
        RECT 1.465 0.525 1.535 0.92 ;
        RECT 0.925 0.525 0.995 0.92 ;
        RECT 0.77 0.525 0.995 0.7 ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.2 0.15 1.29 0.785 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.71 1.485 ;
        RECT 1.405 1.205 1.475 1.485 ;
        RECT 1.035 1.205 1.105 1.485 ;
        RECT 0.24 1.24 0.375 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.71 0.085 ;
        RECT 1.405 -0.085 1.475 0.285 ;
        RECT 1.03 -0.085 1.1 0.285 ;
        RECT 0.46 -0.085 0.53 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.6 0.15 1.67 1.25 ;
      RECT 0.79 0.985 1.67 1.055 ;
      RECT 0.79 0.765 0.86 1.055 ;
      RECT 0.425 0.765 0.86 0.835 ;
      RECT 0.425 0.525 0.495 0.835 ;
      RECT 0.655 0.9 0.725 1.075 ;
      RECT 0.29 0.9 0.725 0.97 ;
      RECT 0.29 0.385 0.36 0.97 ;
      RECT 1.065 0.385 1.135 0.66 ;
      RECT 0.09 0.385 1.135 0.455 ;
      RECT 0.845 0.15 0.915 0.455 ;
      RECT 0.09 0.15 0.16 0.455 ;
      RECT 0.46 1.175 0.955 1.245 ;
      RECT 0.46 1.065 0.53 1.245 ;
      RECT 0.09 1.065 0.53 1.135 ;
      RECT 0.09 0.86 0.16 1.135 ;
  END
END MUX2_X2

MACRO NAND2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_X1 0 0 ;
  SIZE 0.57 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.385 0.525 0.51 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.355 0.5 0.425 ;
        RECT 0.43 0.15 0.5 0.425 ;
        RECT 0.25 0.355 0.32 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.57 1.485 ;
        RECT 0.43 0.975 0.5 1.485 ;
        RECT 0.055 0.975 0.125 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.57 0.085 ;
        RECT 0.055 -0.085 0.125 0.425 ;
    END
  END VSS
END NAND2_X1

MACRO NAND2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_X2 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.51 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.77 0.81 0.84 ;
        RECT 0.74 0.525 0.81 0.84 ;
        RECT 0.25 0.525 0.32 0.84 ;
        RECT 0.175 0.525 0.32 0.66 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.905 0.7 1.25 ;
        RECT 0.04 0.905 0.7 0.975 ;
        RECT 0.04 0.39 0.51 0.46 ;
        RECT 0.44 0.15 0.51 0.46 ;
        RECT 0.25 0.905 0.32 1.25 ;
        RECT 0.04 0.39 0.11 0.975 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.95 1.485 ;
        RECT 0.82 1.04 0.89 1.485 ;
        RECT 0.44 1.04 0.51 1.485 ;
        RECT 0.065 1.04 0.135 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.95 0.085 ;
        RECT 0.82 -0.085 0.89 0.425 ;
        RECT 0.065 -0.085 0.135 0.285 ;
    END
  END VSS
END NAND2_X2

MACRO NAND2_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_X4 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.01 0.525 1.14 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.38 0.525 0.51 0.7 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.405 0.35 1.475 1.07 ;
        RECT 0.275 0.785 1.475 0.855 ;
        RECT 1.39 0.35 1.475 0.855 ;
        RECT 1 0.35 1.475 0.42 ;
        RECT 1.025 0.785 1.095 1.07 ;
        RECT 0.645 0.785 0.715 1.07 ;
        RECT 0.275 0.785 0.345 1.07 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.71 1.485 ;
        RECT 1.595 1.04 1.665 1.485 ;
        RECT 1.215 1.04 1.285 1.485 ;
        RECT 0.835 1.04 0.905 1.485 ;
        RECT 0.455 1.04 0.525 1.485 ;
        RECT 0.08 1.04 0.15 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.71 0.085 ;
        RECT 0.645 -0.085 0.715 0.285 ;
        RECT 0.265 -0.085 0.335 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.595 0.15 1.665 0.425 ;
      RECT 0.085 0.355 0.905 0.425 ;
      RECT 0.835 0.15 0.905 0.425 ;
      RECT 0.455 0.15 0.525 0.425 ;
      RECT 0.085 0.15 0.155 0.425 ;
      RECT 0.835 0.15 1.665 0.22 ;
  END
END NAND2_X4

MACRO NAND3_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3_X1 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.54 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.375 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.605 0.15 0.675 1.25 ;
        RECT 0.235 0.8 0.675 0.87 ;
        RECT 0.235 0.8 0.32 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
        RECT 0.415 0.975 0.485 1.485 ;
        RECT 0.04 0.975 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
        RECT 0.04 -0.085 0.11 0.425 ;
    END
  END VSS
END NAND3_X1

MACRO NAND3_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3_X2 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.595 0.56 0.73 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.95 0.42 1.08 0.7 ;
        RECT 0.38 0.42 1.08 0.49 ;
        RECT 0.38 0.42 0.45 0.66 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.195 0.77 1.215 0.84 ;
        RECT 1.145 0.525 1.215 0.84 ;
        RECT 0.195 0.7 0.32 0.84 ;
        RECT 0.195 0.525 0.265 0.84 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.025 0.905 1.095 1.25 ;
        RECT 0.06 0.905 1.095 0.975 ;
        RECT 0.06 0.265 0.75 0.335 ;
        RECT 0.645 0.905 0.715 1.25 ;
        RECT 0.265 0.905 0.335 1.25 ;
        RECT 0.06 0.265 0.13 0.975 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.33 1.485 ;
        RECT 1.215 1.04 1.285 1.485 ;
        RECT 0.835 1.04 0.905 1.485 ;
        RECT 0.455 1.04 0.525 1.485 ;
        RECT 0.08 1.04 0.15 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.33 0.085 ;
        RECT 1.215 -0.085 1.285 0.335 ;
        RECT 0.08 -0.085 0.15 0.195 ;
    END
  END VSS
END NAND3_X2

MACRO NAND3_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3_X4 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.66 0.555 1.89 0.625 ;
        RECT 1.66 0.29 1.73 0.625 ;
        RECT 0.82 0.29 1.73 0.36 ;
        RECT 0.625 0.555 0.89 0.625 ;
        RECT 0.82 0.29 0.89 0.625 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.525 0.69 2.13 0.76 ;
        RECT 2.06 0.525 2.13 0.76 ;
        RECT 1.525 0.425 1.595 0.76 ;
        RECT 0.955 0.425 1.595 0.495 ;
        RECT 0.38 0.69 1.08 0.76 ;
        RECT 0.955 0.425 1.08 0.76 ;
        RECT 0.38 0.525 0.45 0.76 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.19 0.825 2.3 0.895 ;
        RECT 2.23 0.525 2.3 0.895 ;
        RECT 1.19 0.56 1.325 0.895 ;
        RECT 0.19 0.525 0.26 0.895 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.055 0.98 2.435 1.05 ;
        RECT 2.365 0.355 2.435 1.05 ;
        RECT 1.795 0.355 2.435 0.425 ;
        RECT 2.165 0.98 2.235 1.22 ;
        RECT 0.265 0.98 2.235 1.12 ;
        RECT 1.795 0.15 1.865 0.425 ;
        RECT 1.785 0.98 1.855 1.22 ;
        RECT 1.405 0.98 1.475 1.22 ;
        RECT 1.025 0.98 1.095 1.22 ;
        RECT 0.645 0.98 0.715 1.22 ;
        RECT 0.055 0.355 0.715 0.425 ;
        RECT 0.645 0.15 0.715 0.425 ;
        RECT 0.265 0.98 0.335 1.22 ;
        RECT 0.055 0.355 0.125 1.05 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.47 1.485 ;
        RECT 2.355 1.17 2.425 1.485 ;
        RECT 1.945 1.205 2.08 1.485 ;
        RECT 1.565 1.205 1.7 1.485 ;
        RECT 1.185 1.205 1.32 1.485 ;
        RECT 0.805 1.195 0.94 1.485 ;
        RECT 0.425 1.195 0.56 1.485 ;
        RECT 0.08 1.16 0.15 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.47 0.085 ;
        RECT 2.355 -0.085 2.425 0.195 ;
        RECT 1.215 -0.085 1.285 0.195 ;
        RECT 0.08 -0.085 0.15 0.195 ;
    END
  END VSS
END NAND3_X4

MACRO NAND4_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4_X1 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765 0.525 0.89 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.42 0.555 0.66 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.42 0.375 0.66 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.42 0.185 0.66 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.355 0.865 0.425 ;
        RECT 0.795 0.15 0.865 0.425 ;
        RECT 0.615 0.84 0.7 1.25 ;
        RECT 0.63 0.355 0.7 1.25 ;
        RECT 0.235 0.84 0.7 0.91 ;
        RECT 0.235 0.84 0.305 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.95 1.485 ;
        RECT 0.795 0.975 0.865 1.485 ;
        RECT 0.415 0.975 0.485 1.485 ;
        RECT 0.04 0.975 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.95 0.085 ;
        RECT 0.04 -0.085 0.11 0.355 ;
    END
  END VSS
END NAND4_X1

MACRO NAND4_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4_X2 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.81 0.42 0.945 0.625 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.145 0.285 1.27 0.66 ;
        RECT 0.575 0.285 1.27 0.355 ;
        RECT 0.575 0.285 0.645 0.66 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.39 0.725 1.405 0.795 ;
        RECT 1.335 0.525 1.405 0.795 ;
        RECT 0.39 0.525 0.51 0.795 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.195 0.86 1.59 0.93 ;
        RECT 1.52 0.525 1.59 0.93 ;
        RECT 0.195 0.525 0.32 0.93 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.375 0.995 1.51 1.25 ;
        RECT 0.06 0.995 1.51 1.065 ;
        RECT 0.995 0.995 1.13 1.25 ;
        RECT 0.285 0.15 0.94 0.22 ;
        RECT 0.615 0.995 0.75 1.25 ;
        RECT 0.235 0.995 0.37 1.25 ;
        RECT 0.06 0.39 0.355 0.46 ;
        RECT 0.285 0.15 0.355 0.46 ;
        RECT 0.06 0.39 0.13 1.065 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.71 1.485 ;
        RECT 1.595 1.065 1.665 1.485 ;
        RECT 1.215 1.13 1.285 1.485 ;
        RECT 0.835 1.13 0.905 1.485 ;
        RECT 0.455 1.13 0.525 1.485 ;
        RECT 0.08 1.13 0.15 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.71 0.085 ;
        RECT 1.595 -0.085 1.665 0.39 ;
        RECT 0.08 -0.085 0.15 0.25 ;
    END
  END VSS
END NAND4_X2

MACRO NAND4_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4_X4 0 0 ;
  SIZE 3.42 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.405 0.525 0.51 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.17 0.525 1.27 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.15 0.525 2.22 0.7 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.91 0.525 2.98 0.7 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.27 0.84 3.34 1.155 ;
        RECT 0.09 0.84 3.34 0.98 ;
        RECT 2.89 0.84 2.96 1.155 ;
        RECT 2.51 0.84 2.58 1.155 ;
        RECT 2.13 0.84 2.2 1.155 ;
        RECT 1.68 0.84 1.75 1.155 ;
        RECT 1.22 0.84 1.29 1.155 ;
        RECT 0.84 0.84 0.91 1.155 ;
        RECT 0.685 0.285 0.755 0.98 ;
        RECT 0.225 0.285 0.755 0.355 ;
        RECT 0.46 0.84 0.53 1.155 ;
        RECT 0.09 0.84 0.16 1.155 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 3.42 1.485 ;
        RECT 3.05 1.095 3.185 1.485 ;
        RECT 2.67 1.095 2.805 1.485 ;
        RECT 2.29 1.095 2.425 1.485 ;
        RECT 1.91 1.095 2.045 1.485 ;
        RECT 1.38 1.095 1.515 1.485 ;
        RECT 1 1.095 1.135 1.485 ;
        RECT 0.62 1.095 0.755 1.485 ;
        RECT 0.24 1.095 0.375 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 3.42 0.085 ;
        RECT 3.05 -0.085 3.185 0.3 ;
        RECT 2.67 -0.085 2.805 0.3 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 2.51 0.39 3.34 0.46 ;
      RECT 3.27 0.185 3.34 0.46 ;
      RECT 1.76 0.15 1.83 0.46 ;
      RECT 2.89 0.185 2.96 0.46 ;
      RECT 2.51 0.15 2.58 0.46 ;
      RECT 1.76 0.15 2.58 0.22 ;
      RECT 1.38 0.525 2.045 0.595 ;
      RECT 1.91 0.285 2.045 0.595 ;
      RECT 1.38 0.285 1.515 0.595 ;
      RECT 1.91 0.285 2.425 0.355 ;
      RECT 1.005 0.285 1.515 0.355 ;
      RECT 1.6 0.15 1.67 0.46 ;
      RECT 0.84 0.15 0.91 0.46 ;
      RECT 0.09 0.15 0.16 0.46 ;
      RECT 0.09 0.15 1.67 0.22 ;
  END
END NAND4_X4

MACRO NOR2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_X1 0 0 ;
  SIZE 0.57 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.385 0.525 0.51 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.43 0.975 0.5 1.25 ;
        RECT 0.25 0.975 0.5 1.045 ;
        RECT 0.25 0.15 0.32 1.045 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.57 1.485 ;
        RECT 0.055 0.975 0.125 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.57 0.085 ;
        RECT 0.43 -0.085 0.5 0.425 ;
        RECT 0.055 -0.085 0.125 0.425 ;
    END
  END VSS
END NOR2_X1

MACRO NOR2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_X2 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.42 0.51 0.66 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.195 0.725 0.89 0.795 ;
        RECT 0.76 0.525 0.89 0.795 ;
        RECT 0.195 0.525 0.265 0.795 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.26 0.75 0.33 ;
        RECT 0.455 0.91 0.525 1.25 ;
        RECT 0.06 0.91 0.525 0.98 ;
        RECT 0.06 0.26 0.13 0.98 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.95 1.485 ;
        RECT 0.835 1.045 0.905 1.485 ;
        RECT 0.08 1.045 0.15 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.95 0.085 ;
        RECT 0.835 -0.085 0.905 0.335 ;
        RECT 0.455 -0.085 0.525 0.195 ;
        RECT 0.08 -0.085 0.15 0.195 ;
    END
  END VSS
END NOR2_X2

MACRO NOR2_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_X4 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.09 0.42 1.16 0.66 ;
        RECT 0.59 0.42 1.16 0.49 ;
        RECT 0.59 0.42 0.7 0.66 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.215 0.91 1.535 0.98 ;
        RECT 1.465 0.525 1.535 0.98 ;
        RECT 0.805 0.56 0.94 0.98 ;
        RECT 0.215 0.525 0.285 0.98 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.24 0.28 1.51 0.35 ;
        RECT 1.225 0.28 1.295 0.845 ;
        RECT 0.44 0.28 0.525 0.845 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.71 1.485 ;
        RECT 1.6 0.71 1.67 1.485 ;
        RECT 0.835 1.045 0.905 1.485 ;
        RECT 0.08 0.71 0.15 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.71 0.085 ;
        RECT 1.595 -0.085 1.665 0.39 ;
        RECT 1.215 -0.085 1.285 0.195 ;
        RECT 0.835 -0.085 0.905 0.195 ;
        RECT 0.455 -0.085 0.525 0.195 ;
        RECT 0.08 -0.085 0.15 0.39 ;
    END
  END VSS
END NOR2_X4

MACRO NOR3_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3_X1 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.545 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.375 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.175 0.7 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.61 0.15 0.7 1 ;
        RECT 0.235 0.355 0.7 0.425 ;
        RECT 0.235 0.15 0.305 0.425 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
        RECT 0.04 0.975 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
        RECT 0.415 -0.085 0.485 0.22 ;
        RECT 0.04 -0.085 0.11 0.425 ;
    END
  END VSS
END NOR3_X1

MACRO NOR3_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3_X2 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.62 0.56 0.755 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.92 0.425 0.99 0.66 ;
        RECT 0.39 0.425 0.99 0.495 ;
        RECT 0.39 0.425 0.51 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.195 0.77 1.27 0.84 ;
        RECT 1.145 0.525 1.27 0.84 ;
        RECT 0.195 0.525 0.265 0.84 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.285 1.13 0.355 ;
        RECT 0.645 0.905 0.715 1.18 ;
        RECT 0.06 0.905 0.715 0.975 ;
        RECT 0.06 0.285 0.13 0.975 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.33 1.485 ;
        RECT 1.215 1.065 1.285 1.485 ;
        RECT 0.08 1.065 0.15 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.33 0.085 ;
        RECT 1.215 -0.085 1.285 0.335 ;
        RECT 0.835 -0.085 0.905 0.195 ;
        RECT 0.455 -0.085 0.525 0.195 ;
        RECT 0.08 -0.085 0.15 0.195 ;
    END
  END VSS
END NOR3_X2

MACRO NOR3_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3_X4 0 0 ;
  SIZE 2.66 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425 0.525 0.51 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.185 0.525 1.27 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.13 0.525 2.23 0.7 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235 0.39 2.38 0.46 ;
        RECT 2.31 0.15 2.38 0.46 ;
        RECT 1.93 0.15 2 0.46 ;
        RECT 1.365 0.15 1.435 0.46 ;
        RECT 0.985 0.15 1.055 0.46 ;
        RECT 0.605 0.765 0.675 1.115 ;
        RECT 0.605 0.15 0.675 0.46 ;
        RECT 0.235 0.765 0.675 0.835 ;
        RECT 0.235 0.39 0.32 0.835 ;
        RECT 0.235 0.15 0.305 1.115 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.66 1.485 ;
        RECT 2.5 0.9 2.57 1.485 ;
        RECT 2.09 0.935 2.225 1.485 ;
        RECT 1.745 0.9 1.815 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.66 0.085 ;
        RECT 2.505 -0.085 2.575 0.425 ;
        RECT 2.09 -0.085 2.225 0.325 ;
        RECT 1.525 -0.085 1.85 0.325 ;
        RECT 1.145 -0.085 1.28 0.325 ;
        RECT 0.765 -0.085 0.9 0.325 ;
        RECT 0.385 -0.085 0.52 0.325 ;
        RECT 0.04 -0.085 0.11 0.425 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 2.31 0.765 2.38 1.175 ;
      RECT 1.93 0.765 2 1.175 ;
      RECT 1.365 0.765 1.435 1.115 ;
      RECT 0.995 0.765 1.065 1.115 ;
      RECT 0.995 0.765 2.38 0.835 ;
      RECT 0.045 1.18 1.625 1.25 ;
      RECT 1.555 0.9 1.625 1.25 ;
      RECT 1.175 0.9 1.245 1.25 ;
      RECT 0.795 0.9 0.865 1.25 ;
      RECT 0.415 0.9 0.485 1.25 ;
      RECT 0.045 0.9 0.115 1.25 ;
  END
END NOR3_X4

MACRO NOR4_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4_X1 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765 0.525 0.89 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.565 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.375 0.7 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.795 0.975 0.865 1.25 ;
        RECT 0.63 0.975 0.865 1.045 ;
        RECT 0.63 0.15 0.7 1.045 ;
        RECT 0.235 0.355 0.7 0.425 ;
        RECT 0.61 0.15 0.7 0.425 ;
        RECT 0.235 0.15 0.305 0.425 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.95 1.485 ;
        RECT 0.04 0.975 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.95 0.085 ;
        RECT 0.795 -0.085 0.865 0.425 ;
        RECT 0.415 -0.085 0.485 0.285 ;
        RECT 0.04 -0.085 0.11 0.425 ;
    END
  END VSS
END NOR4_X1

MACRO NOR4_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4_X2 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.81 0.56 0.945 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.11 0.42 1.18 0.66 ;
        RECT 0.57 0.42 1.18 0.49 ;
        RECT 0.57 0.42 0.7 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.38 0.765 1.46 0.835 ;
        RECT 1.33 0.525 1.46 0.835 ;
        RECT 0.38 0.525 0.45 0.835 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.2 0.91 1.65 0.98 ;
        RECT 1.525 0.84 1.65 0.98 ;
        RECT 1.525 0.525 1.595 0.98 ;
        RECT 0.2 0.525 0.27 0.98 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.405 0.15 1.475 0.425 ;
        RECT 0.055 0.26 1.475 0.33 ;
        RECT 0.055 1.055 0.94 1.125 ;
        RECT 0.055 0.26 0.13 1.125 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.71 1.485 ;
        RECT 1.595 1.065 1.665 1.485 ;
        RECT 0.08 1.205 0.15 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.71 0.085 ;
        RECT 1.595 -0.085 1.665 0.335 ;
        RECT 1.185 -0.085 1.32 0.16 ;
        RECT 0.805 -0.085 0.94 0.16 ;
        RECT 0.425 -0.085 0.56 0.16 ;
        RECT 0.08 -0.085 0.15 0.195 ;
    END
  END VSS
END NOR4_X2

MACRO NOR4_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4_X4 0 0 ;
  SIZE 3.42 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425 0.525 0.51 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.18 0.525 1.27 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.15 0.525 2.245 0.7 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.91 0.525 3 0.7 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235 0.39 3.375 0.46 ;
        RECT 3.305 0.15 3.375 0.46 ;
        RECT 2.925 0.15 2.995 0.46 ;
        RECT 2.545 0.15 2.615 0.46 ;
        RECT 2.165 0.15 2.235 0.46 ;
        RECT 1.79 0.15 1.86 0.46 ;
        RECT 1.37 0.15 1.44 0.46 ;
        RECT 0.985 0.15 1.055 0.46 ;
        RECT 0.605 0.765 0.675 1.115 ;
        RECT 0.605 0.15 0.675 0.46 ;
        RECT 0.235 0.765 0.675 0.835 ;
        RECT 0.235 0.39 0.32 0.835 ;
        RECT 0.235 0.15 0.305 1.115 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 3.42 1.485 ;
        RECT 3.085 0.935 3.22 1.485 ;
        RECT 2.705 0.935 2.84 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 3.42 0.085 ;
        RECT 3.085 -0.085 3.22 0.325 ;
        RECT 2.705 -0.085 2.84 0.325 ;
        RECT 2.325 -0.085 2.46 0.325 ;
        RECT 1.945 -0.085 2.08 0.325 ;
        RECT 1.525 -0.085 1.66 0.325 ;
        RECT 1.145 -0.085 1.28 0.325 ;
        RECT 0.765 -0.085 0.9 0.325 ;
        RECT 0.385 -0.085 0.52 0.325 ;
        RECT 0.04 -0.085 0.11 0.36 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 3.305 0.765 3.375 1.175 ;
      RECT 2.925 0.765 2.995 1.175 ;
      RECT 2.545 0.765 2.615 1.175 ;
      RECT 2.165 0.765 2.235 1.115 ;
      RECT 1.795 0.765 1.865 1.115 ;
      RECT 1.795 0.765 3.375 0.835 ;
      RECT 0.995 1.18 2.425 1.25 ;
      RECT 2.355 0.9 2.425 1.25 ;
      RECT 1.975 0.9 2.045 1.25 ;
      RECT 1.365 0.9 1.435 1.25 ;
      RECT 0.995 0.9 1.065 1.25 ;
      RECT 0.045 1.18 0.865 1.25 ;
      RECT 0.795 0.765 0.865 1.25 ;
      RECT 0.415 0.9 0.485 1.25 ;
      RECT 0.045 0.9 0.115 1.25 ;
      RECT 1.555 0.765 1.625 1.115 ;
      RECT 1.175 0.765 1.245 1.115 ;
      RECT 0.795 0.765 1.625 0.835 ;
  END
END NOR4_X4

MACRO OAI211_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211_X1 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.575 0.525 0.7 0.7 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.79 0.525 0.89 0.7 ;
    END
  END B
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.4 0.525 0.51 0.7 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.835 0.78 0.905 1.055 ;
        RECT 0.25 0.78 0.905 0.85 ;
        RECT 0.455 0.78 0.525 1.055 ;
        RECT 0.25 0.78 0.525 0.855 ;
        RECT 0.25 0.285 0.335 0.855 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.95 1.485 ;
        RECT 0.645 1.04 0.715 1.485 ;
        RECT 0.08 1.04 0.15 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.95 0.085 ;
        RECT 0.835 -0.085 0.905 0.46 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.455 0.15 0.525 0.425 ;
      RECT 0.085 0.15 0.155 0.425 ;
      RECT 0.085 0.15 0.525 0.22 ;
  END
END OAI211_X1

MACRO OAI211_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211_X2 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.185 0.765 0.755 0.835 ;
        RECT 0.685 0.525 0.755 0.835 ;
        RECT 0.185 0.525 0.32 0.835 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.53 0.7 ;
    END
  END B
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.19 0.525 1.29 0.7 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.96 0.77 1.65 0.84 ;
        RECT 1.525 0.525 1.65 0.84 ;
        RECT 0.96 0.525 1.03 0.84 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.82 0.39 1.51 0.46 ;
        RECT 1.215 0.905 1.285 1.25 ;
        RECT 0.27 0.905 1.285 0.975 ;
        RECT 0.82 0.39 0.89 0.975 ;
        RECT 0.645 0.905 0.715 1.25 ;
        RECT 0.27 0.905 0.34 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.71 1.485 ;
        RECT 1.595 1.04 1.665 1.485 ;
        RECT 0.835 1.04 0.905 1.485 ;
        RECT 0.455 1.04 0.525 1.485 ;
        RECT 0.08 1.04 0.15 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.71 0.085 ;
        RECT 0.45 -0.085 0.52 0.32 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.595 0.185 1.665 0.46 ;
      RECT 0.08 0.39 0.66 0.46 ;
      RECT 0.59 0.185 0.66 0.46 ;
      RECT 0.08 0.185 0.15 0.46 ;
      RECT 0.59 0.185 1.665 0.255 ;
  END
END OAI211_X2

MACRO OAI211_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211_X4 0 0 ;
  SIZE 3.23 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.39 0.39 1.52 0.66 ;
        RECT 0.125 0.39 1.52 0.46 ;
        RECT 0.805 0.39 0.875 0.66 ;
        RECT 0.125 0.39 0.195 0.66 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.42 0.77 1.245 0.84 ;
        RECT 1.175 0.525 1.245 0.84 ;
        RECT 0.42 0.525 0.51 0.84 ;
    END
  END B
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.91 0.77 2.8 0.84 ;
        RECT 2.665 0.56 2.8 0.84 ;
        RECT 1.91 0.56 2.045 0.84 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.965 0.425 3.035 0.66 ;
        RECT 1.67 0.425 3.035 0.495 ;
        RECT 2.31 0.425 2.41 0.7 ;
        RECT 1.67 0.425 1.74 0.66 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235 0.905 3.17 0.975 ;
        RECT 3.1 0.29 3.17 0.975 ;
        RECT 1.72 0.29 3.17 0.36 ;
        RECT 2.695 0.905 2.765 1.25 ;
        RECT 1.935 0.905 2.005 1.25 ;
        RECT 1.365 0.905 1.435 1.25 ;
        RECT 0.985 0.905 1.055 1.25 ;
        RECT 0.605 0.905 0.675 1.25 ;
        RECT 0.235 0.905 0.305 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 3.23 1.485 ;
        RECT 3.075 1.04 3.145 1.485 ;
        RECT 2.315 1.04 2.385 1.485 ;
        RECT 1.555 1.04 1.625 1.485 ;
        RECT 1.175 1.04 1.245 1.485 ;
        RECT 0.795 1.04 0.865 1.485 ;
        RECT 0.415 1.04 0.485 1.485 ;
        RECT 0.04 1.04 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 3.23 0.085 ;
        RECT 1.145 -0.085 1.28 0.16 ;
        RECT 0.385 -0.085 0.52 0.16 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.225 1.625 0.295 ;
      RECT 1.555 0.15 1.625 0.295 ;
      RECT 0.045 0.15 0.115 0.295 ;
      RECT 1.555 0.15 3.18 0.22 ;
  END
END OAI211_X4

MACRO OAI21_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21_X1 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.575 0.525 0.7 0.7 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.385 0.525 0.51 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.765 0.51 1.25 ;
        RECT 0.25 0.765 0.51 0.835 ;
        RECT 0.25 0.285 0.32 0.835 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
        RECT 0.63 0.975 0.7 1.485 ;
        RECT 0.065 0.975 0.135 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
        RECT 0.63 -0.085 0.7 0.46 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.44 0.15 0.51 0.425 ;
      RECT 0.07 0.15 0.14 0.425 ;
      RECT 0.07 0.15 0.51 0.22 ;
  END
END OAI21_X1

MACRO OAI21_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21_X2 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.19 0.7 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.805 0.525 0.89 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.77 1.135 0.84 ;
        RECT 1.065 0.525 1.135 0.84 ;
        RECT 0.44 0.525 0.57 0.84 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235 0.905 1.27 0.975 ;
        RECT 1.2 0.355 1.27 0.975 ;
        RECT 0.58 0.355 1.27 0.425 ;
        RECT 0.795 0.905 0.865 1.25 ;
        RECT 0.235 0.905 0.305 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.33 1.485 ;
        RECT 1.175 1.04 1.245 1.485 ;
        RECT 0.415 1.04 0.485 1.485 ;
        RECT 0.04 1.04 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.33 0.085 ;
        RECT 0.225 -0.085 0.295 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.355 0.485 0.425 ;
      RECT 0.415 0.15 0.485 0.425 ;
      RECT 0.045 0.15 0.115 0.425 ;
      RECT 0.415 0.15 1.28 0.22 ;
  END
END OAI21_X2

MACRO OAI21_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21_X4 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.43 0.525 0.515 0.7 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.15 0.69 2.04 0.76 ;
        RECT 1.905 0.56 2.04 0.76 ;
        RECT 1.15 0.56 1.285 0.76 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.15 0.42 2.275 0.66 ;
        RECT 0.91 0.42 2.275 0.49 ;
        RECT 1.525 0.42 1.66 0.625 ;
        RECT 0.91 0.42 0.98 0.66 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235 0.845 2.41 0.915 ;
        RECT 2.34 0.285 2.41 0.915 ;
        RECT 0.96 0.285 2.41 0.355 ;
        RECT 1.935 0.845 2.005 1.19 ;
        RECT 1.175 0.845 1.245 1.19 ;
        RECT 0.605 0.845 0.675 1.19 ;
        RECT 0.235 0.845 0.305 1.19 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.47 1.485 ;
        RECT 2.315 1.04 2.385 1.485 ;
        RECT 1.555 1.04 1.625 1.485 ;
        RECT 0.795 1.04 0.865 1.485 ;
        RECT 0.415 1.04 0.485 1.485 ;
        RECT 0.04 1.04 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.47 0.085 ;
        RECT 0.605 -0.085 0.675 0.285 ;
        RECT 0.225 -0.085 0.295 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.355 0.83 0.425 ;
      RECT 0.76 0.15 0.83 0.425 ;
      RECT 0.42 0.15 0.49 0.425 ;
      RECT 0.045 0.15 0.115 0.425 ;
      RECT 0.76 0.15 2.42 0.22 ;
  END
END OAI21_X4

MACRO OAI221_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221_X1 0 0 ;
  SIZE 1.14 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.565 0.7 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.375 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.955 0.525 1.08 0.7 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.525 0.74 0.7 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.985 0.85 1.055 1.25 ;
        RECT 0.425 0.85 1.055 0.92 ;
        RECT 0.805 0.4 0.89 0.92 ;
        RECT 0.425 0.85 0.495 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.14 1.485 ;
        RECT 0.605 1.04 0.675 1.485 ;
        RECT 0.04 1.04 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.14 0.085 ;
        RECT 0.225 -0.085 0.295 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.985 0.15 1.055 0.425 ;
      RECT 0.615 0.15 0.685 0.425 ;
      RECT 0.615 0.15 1.055 0.22 ;
      RECT 0.045 0.355 0.485 0.425 ;
      RECT 0.415 0.15 0.485 0.425 ;
      RECT 0.045 0.15 0.115 0.425 ;
  END
END OAI221_X1

MACRO OAI221_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221_X2 0 0 ;
  SIZE 2.09 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.955 0.9 2.03 0.97 ;
        RECT 1.93 0.525 2.03 0.97 ;
        RECT 0.955 0.525 1.025 0.97 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.155 0.765 1.84 0.835 ;
        RECT 1.715 0.525 1.84 0.835 ;
        RECT 1.155 0.525 1.225 0.835 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.38 0.525 1.48 0.7 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.525 0.7 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.195 0.77 0.89 0.84 ;
        RECT 0.76 0.525 0.89 0.84 ;
        RECT 0.195 0.525 0.265 0.84 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.755 1.035 1.89 1.245 ;
        RECT 0.06 1.035 1.89 1.105 ;
        RECT 0.995 1.035 1.13 1.245 ;
        RECT 0.06 0.39 0.75 0.46 ;
        RECT 0.425 1.035 0.56 1.245 ;
        RECT 0.06 0.39 0.13 1.105 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.09 1.485 ;
        RECT 1.975 1.065 2.045 1.485 ;
        RECT 1.405 1.17 1.475 1.485 ;
        RECT 0.835 1.17 0.905 1.485 ;
        RECT 0.085 1.17 0.155 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.09 0.085 ;
        RECT 1.565 -0.085 1.7 0.19 ;
        RECT 1.185 -0.085 1.32 0.19 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.975 0.15 2.045 0.425 ;
      RECT 0.05 0.255 2.045 0.325 ;
      RECT 1 0.39 1.89 0.46 ;
  END
END OAI221_X2

MACRO OAI221_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221_X4 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.585 0.525 0.7 0.7 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.775 0.525 0.9 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.01 0.525 1.155 0.7 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.245 0.7 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.395 0.525 0.51 0.7 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.165 0.185 2.235 1.25 ;
        RECT 1.795 0.7 2.235 0.84 ;
        RECT 1.795 0.185 1.865 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.47 1.485 ;
        RECT 2.355 0.975 2.425 1.485 ;
        RECT 1.975 0.975 2.045 1.485 ;
        RECT 1.595 0.975 1.665 1.485 ;
        RECT 1.19 1.04 1.26 1.485 ;
        RECT 0.47 1.04 0.54 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.47 0.085 ;
        RECT 2.355 -0.085 2.425 0.46 ;
        RECT 1.975 -0.085 2.045 0.46 ;
        RECT 1.595 -0.085 1.665 0.335 ;
        RECT 1.19 -0.085 1.26 0.2 ;
        RECT 0.82 -0.085 0.955 0.16 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.415 0.185 1.485 1.25 ;
      RECT 1.415 0.525 1.73 0.66 ;
      RECT 0.66 0.775 0.73 1.12 ;
      RECT 0.1 0.775 0.17 1.12 ;
      RECT 0.1 0.775 1.35 0.845 ;
      RECT 1.28 0.39 1.35 0.845 ;
      RECT 0.29 0.39 1.35 0.46 ;
      RECT 0.29 0.285 0.36 0.46 ;
      RECT 0.67 0.255 1.11 0.325 ;
      RECT 0.67 0.15 0.74 0.325 ;
      RECT 0.47 0.15 0.54 0.285 ;
      RECT 0.1 0.15 0.17 0.285 ;
      RECT 0.1 0.15 0.54 0.22 ;
  END
END OAI221_X4

MACRO OAI222_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222_X1 0 0 ;
  SIZE 1.52 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.34 0.525 1.46 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.01 0.525 1.115 0.7 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.525 0.755 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.82 0.525 0.945 0.7 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.35 0.525 0.51 0.7 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.2 0.7 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.36 0.795 1.43 1.14 ;
        RECT 0.52 0.795 1.43 0.865 ;
        RECT 1.18 0.4 1.27 0.865 ;
        RECT 0.52 0.795 0.59 1.14 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.52 1.485 ;
        RECT 0.98 1.04 1.05 1.485 ;
        RECT 0.05 1.04 0.12 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.52 0.085 ;
        RECT 0.395 -0.085 0.53 0.19 ;
        RECT 0.05 -0.085 0.12 0.425 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.575 0.39 1.05 0.46 ;
      RECT 0.98 0.15 1.05 0.46 ;
      RECT 1.36 0.15 1.43 0.425 ;
      RECT 0.98 0.265 1.43 0.335 ;
      RECT 0.245 0.15 0.315 0.425 ;
      RECT 0.245 0.255 0.86 0.325 ;
      RECT 0.79 0.15 0.86 0.325 ;
  END
END OAI222_X1

MACRO OAI222_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222_X2 0 0 ;
  SIZE 2.66 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.85 0.725 2.465 0.795 ;
        RECT 2.34 0.525 2.465 0.795 ;
        RECT 1.85 0.525 1.92 0.795 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.15 0.42 2.22 0.66 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.955 0.77 1.65 0.84 ;
        RECT 1.525 0.525 1.65 0.84 ;
        RECT 0.955 0.525 1.025 0.84 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.2 0.525 1.29 0.7 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.195 0.77 0.83 0.84 ;
        RECT 0.76 0.525 0.83 0.84 ;
        RECT 0.195 0.525 0.32 0.84 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.53 0.7 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.53 0.285 2.6 1.25 ;
        RECT 0.09 0.905 2.6 0.975 ;
        RECT 1.925 0.285 2.6 0.355 ;
        RECT 1.605 0.905 1.675 1.25 ;
        RECT 0.84 0.905 0.91 1.25 ;
        RECT 0.09 0.905 0.16 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.66 1.485 ;
        RECT 2.14 1.04 2.21 1.485 ;
        RECT 1.22 1.04 1.29 1.485 ;
        RECT 0.46 1.04 0.53 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.66 0.085 ;
        RECT 0.65 -0.085 0.72 0.285 ;
        RECT 0.27 -0.085 0.34 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.005 0.355 1.84 0.425 ;
      RECT 1.77 0.15 1.84 0.425 ;
      RECT 1.77 0.15 2.625 0.22 ;
      RECT 0.09 0.355 0.91 0.425 ;
      RECT 0.84 0.15 0.91 0.425 ;
      RECT 0.465 0.15 0.535 0.425 ;
      RECT 0.09 0.15 0.16 0.425 ;
      RECT 0.84 0.15 1.705 0.22 ;
  END
END OAI222_X2

MACRO OAI222_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222_X4 0 0 ;
  SIZE 2.66 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.38 0.7 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765 0.56 0.9 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.495 0.56 0.7 0.7 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.995 0.56 1.13 0.7 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.195 0.56 1.33 0.7 ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.29 0.15 2.36 1.25 ;
        RECT 1.915 0.56 2.36 0.7 ;
        RECT 1.915 0.15 1.985 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.66 1.485 ;
        RECT 2.475 0.975 2.545 1.485 ;
        RECT 2.095 0.975 2.165 1.485 ;
        RECT 1.715 0.975 1.785 1.485 ;
        RECT 1.335 1.04 1.405 1.485 ;
        RECT 0.415 1.03 0.485 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.66 0.085 ;
        RECT 2.475 -0.085 2.545 0.425 ;
        RECT 2.095 -0.085 2.165 0.425 ;
        RECT 1.715 -0.085 1.785 0.335 ;
        RECT 1.335 -0.085 1.405 0.22 ;
        RECT 0.965 -0.085 1.035 0.22 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.535 0.15 1.605 1.16 ;
      RECT 1.535 0.525 1.85 0.66 ;
      RECT 0.88 0.785 0.95 1.075 ;
      RECT 0.045 0.785 0.115 1.075 ;
      RECT 0.045 0.785 1.465 0.855 ;
      RECT 1.395 0.285 1.465 0.855 ;
      RECT 0.2 0.285 1.465 0.355 ;
      RECT 0.045 0.15 0.115 0.425 ;
      RECT 0.045 0.15 0.9 0.22 ;
      RECT 0.58 0.42 1.25 0.49 ;
  END
END OAI222_X4

MACRO OAI22_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22_X1 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.575 0.525 0.7 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765 0.525 0.89 0.7 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.375 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.39 0.725 0.46 ;
        RECT 0.44 0.39 0.51 1.05 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.95 1.485 ;
        RECT 0.81 0.975 0.88 1.485 ;
        RECT 0.055 0.975 0.125 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.95 0.085 ;
        RECT 0.21 -0.085 0.345 0.16 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.81 0.185 0.88 0.46 ;
      RECT 0.06 0.185 0.13 0.46 ;
      RECT 0.06 0.245 0.88 0.315 ;
  END
END OAI22_X1

MACRO OAI22_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22_X2 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.185 0.525 1.27 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.82 0.765 1.515 0.835 ;
        RECT 1.445 0.525 1.515 0.835 ;
        RECT 0.82 0.525 0.95 0.835 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425 0.525 0.525 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.765 0.75 0.835 ;
        RECT 0.68 0.525 0.75 0.835 ;
        RECT 0.06 0.525 0.185 0.835 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425 0.9 1.65 0.97 ;
        RECT 1.58 0.39 1.65 0.97 ;
        RECT 0.96 0.39 1.65 0.46 ;
        RECT 1.185 0.9 1.255 1.25 ;
        RECT 0.425 0.9 0.495 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.71 1.485 ;
        RECT 1.555 1.035 1.625 1.485 ;
        RECT 0.795 1.035 0.865 1.485 ;
        RECT 0.04 1.035 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.71 0.085 ;
        RECT 0.605 -0.085 0.675 0.285 ;
        RECT 0.225 -0.085 0.295 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.355 0.865 0.425 ;
      RECT 0.795 0.15 0.865 0.425 ;
      RECT 0.415 0.15 0.485 0.425 ;
      RECT 0.045 0.15 0.115 0.425 ;
      RECT 0.795 0.15 1.66 0.22 ;
  END
END OAI22_X2

MACRO OAI22_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22_X4 0 0 ;
  SIZE 3.23 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.91 0.725 2.805 0.795 ;
        RECT 2.67 0.56 2.805 0.795 ;
        RECT 1.91 0.56 2.045 0.795 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.91 0.425 3.035 0.7 ;
        RECT 1.645 0.425 3.035 0.495 ;
        RECT 2.32 0.425 2.39 0.66 ;
        RECT 1.645 0.425 1.715 0.66 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.385 0.725 1.28 0.795 ;
        RECT 1.145 0.56 1.28 0.795 ;
        RECT 0.385 0.56 0.52 0.795 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.39 0.425 1.52 0.7 ;
        RECT 0.15 0.425 1.52 0.495 ;
        RECT 0.795 0.425 0.865 0.66 ;
        RECT 0.15 0.425 0.22 0.66 ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425 0.865 3.17 0.935 ;
        RECT 3.1 0.29 3.17 0.935 ;
        RECT 1.72 0.29 3.17 0.36 ;
        RECT 2.695 0.865 2.765 1.21 ;
        RECT 1.935 0.865 2.005 1.21 ;
        RECT 1.175 0.865 1.245 1.21 ;
        RECT 0.425 0.865 0.495 1.21 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 3.23 1.485 ;
        RECT 3.075 1.04 3.145 1.485 ;
        RECT 2.315 1.04 2.385 1.485 ;
        RECT 1.555 1.04 1.625 1.485 ;
        RECT 0.795 1.04 0.865 1.485 ;
        RECT 0.04 1.04 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 3.23 0.085 ;
        RECT 1.365 -0.085 1.435 0.195 ;
        RECT 0.985 -0.085 1.055 0.195 ;
        RECT 0.605 -0.085 0.675 0.195 ;
        RECT 0.225 -0.085 0.295 0.195 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.26 1.595 0.33 ;
      RECT 1.525 0.15 1.595 0.33 ;
      RECT 0.045 0.185 0.115 0.33 ;
      RECT 1.525 0.15 3.18 0.22 ;
  END
END OAI22_X4

MACRO OAI33_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33_X1 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765 0.525 0.89 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.955 0.525 1.08 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.145 0.525 1.27 0.7 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.565 0.7 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.375 0.7 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.365 1.26 0.435 ;
        RECT 1.19 0.15 1.26 0.435 ;
        RECT 0.63 0.365 0.7 1 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.33 1.485 ;
        RECT 1.19 0.975 1.26 1.485 ;
        RECT 0.055 0.975 0.125 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.33 0.085 ;
        RECT 0.4 -0.085 0.535 0.16 ;
        RECT 0.055 -0.085 0.125 0.335 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.215 0.225 1.105 0.295 ;
  END
END OAI33_X1

MACRO OR2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2_X1 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.38 0.7 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.61 0.15 0.7 1.24 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
        RECT 0.415 0.965 0.485 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
        RECT 0.415 -0.085 0.485 0.285 ;
        RECT 0.04 -0.085 0.11 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.83 0.115 1.24 ;
      RECT 0.045 0.83 0.54 0.9 ;
      RECT 0.47 0.35 0.54 0.9 ;
      RECT 0.235 0.35 0.54 0.42 ;
      RECT 0.235 0.15 0.305 0.42 ;
  END
END OR2_X1

MACRO OR2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2_X2 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.38 0.7 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.615 0.15 0.7 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.95 1.485 ;
        RECT 0.795 0.975 0.865 1.485 ;
        RECT 0.415 1.04 0.485 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.95 0.085 ;
        RECT 0.795 -0.085 0.865 0.425 ;
        RECT 0.415 -0.085 0.485 0.285 ;
        RECT 0.04 -0.085 0.11 0.425 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.905 0.115 1.25 ;
      RECT 0.045 0.905 0.545 0.975 ;
      RECT 0.475 0.355 0.545 0.975 ;
      RECT 0.235 0.355 0.545 0.425 ;
      RECT 0.235 0.15 0.305 0.425 ;
  END
END OR2_X2

MACRO OR2_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2_X4 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.38 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.765 0.76 0.835 ;
        RECT 0.69 0.525 0.76 0.835 ;
        RECT 0.06 0.525 0.15 0.835 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.365 0.15 1.435 1.095 ;
        RECT 0.995 0.56 1.435 0.7 ;
        RECT 0.995 0.15 1.075 0.7 ;
        RECT 0.995 0.15 1.065 1.095 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.71 1.485 ;
        RECT 1.555 1.035 1.625 1.485 ;
        RECT 1.175 1.035 1.245 1.485 ;
        RECT 0.795 1.035 0.865 1.485 ;
        RECT 0.04 1.035 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.71 0.085 ;
        RECT 1.555 -0.085 1.625 0.425 ;
        RECT 1.175 -0.085 1.245 0.425 ;
        RECT 0.795 -0.085 0.865 0.285 ;
        RECT 0.415 -0.085 0.485 0.285 ;
        RECT 0.04 -0.085 0.11 0.425 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.425 0.9 0.495 1.25 ;
      RECT 0.425 0.9 0.925 0.97 ;
      RECT 0.855 0.355 0.925 0.97 ;
      RECT 0.235 0.355 0.925 0.425 ;
      RECT 0.605 0.15 0.675 0.425 ;
      RECT 0.235 0.15 0.305 0.425 ;
  END
END OR2_X4

MACRO OR3_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3_X1 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.375 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.57 0.7 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.8 0.15 0.89 1.24 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.95 1.485 ;
        RECT 0.605 0.965 0.675 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.95 0.085 ;
        RECT 0.605 -0.085 0.675 0.285 ;
        RECT 0.225 -0.085 0.295 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.83 0.115 1.24 ;
      RECT 0.045 0.83 0.73 0.9 ;
      RECT 0.66 0.35 0.73 0.9 ;
      RECT 0.045 0.35 0.73 0.42 ;
      RECT 0.415 0.15 0.485 0.42 ;
      RECT 0.045 0.15 0.115 0.42 ;
  END
END OR3_X1

MACRO OR3_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3_X2 0 0 ;
  SIZE 1.14 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.375 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.57 0.7 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.805 0.15 0.89 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.14 1.485 ;
        RECT 0.985 0.975 1.055 1.485 ;
        RECT 0.605 0.975 0.675 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.14 0.085 ;
        RECT 0.985 -0.085 1.055 0.425 ;
        RECT 0.605 -0.085 0.675 0.285 ;
        RECT 0.225 -0.085 0.295 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.84 0.115 1.25 ;
      RECT 0.045 0.84 0.73 0.91 ;
      RECT 0.66 0.39 0.73 0.91 ;
      RECT 0.045 0.39 0.73 0.46 ;
      RECT 0.415 0.15 0.485 0.46 ;
      RECT 0.045 0.15 0.115 0.46 ;
  END
END OR3_X2

MACRO OR3_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3_X4 0 0 ;
  SIZE 2.09 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.61 0.56 0.745 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.915 0.42 0.985 0.66 ;
        RECT 0.375 0.42 0.985 0.49 ;
        RECT 0.375 0.42 0.51 0.66 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.185 0.77 1.2 0.84 ;
        RECT 1.13 0.525 1.2 0.84 ;
        RECT 0.185 0.7 0.32 0.84 ;
        RECT 0.185 0.525 0.255 0.84 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.79 0.26 1.86 1.25 ;
        RECT 1.415 0.56 1.86 0.7 ;
        RECT 1.415 0.26 1.485 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.09 1.485 ;
        RECT 1.975 1.035 2.045 1.485 ;
        RECT 1.595 1.035 1.665 1.485 ;
        RECT 1.21 1.045 1.28 1.485 ;
        RECT 0.075 1.035 0.145 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.09 0.085 ;
        RECT 1.975 -0.085 2.045 0.335 ;
        RECT 1.595 -0.085 1.665 0.335 ;
        RECT 1.21 -0.085 1.28 0.195 ;
        RECT 0.83 -0.085 0.9 0.195 ;
        RECT 0.45 -0.085 0.52 0.195 ;
        RECT 0.075 -0.085 0.145 0.335 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.65 0.91 0.72 1.25 ;
      RECT 0.65 0.91 1.35 0.98 ;
      RECT 1.28 0.26 1.35 0.98 ;
      RECT 0.235 0.26 1.35 0.33 ;
  END
END OR3_X4

MACRO OR4_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4_X1 0 0 ;
  SIZE 1.14 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.375 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.565 0.7 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.525 0.76 0.7 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.99 0.15 1.08 1.24 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.14 1.485 ;
        RECT 0.795 0.965 0.865 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.14 0.085 ;
        RECT 0.795 -0.085 0.865 0.285 ;
        RECT 0.415 -0.085 0.485 0.285 ;
        RECT 0.04 -0.085 0.11 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.83 0.115 1.24 ;
      RECT 0.045 0.83 0.92 0.9 ;
      RECT 0.85 0.35 0.92 0.9 ;
      RECT 0.235 0.35 0.92 0.42 ;
      RECT 0.605 0.15 0.675 0.42 ;
      RECT 0.235 0.15 0.305 0.42 ;
  END
END OR4_X1

MACRO OR4_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4_X2 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.525 0.375 0.7 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.525 0.565 0.7 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.525 0.76 0.7 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.995 0.15 1.08 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.33 1.485 ;
        RECT 1.175 0.975 1.245 1.485 ;
        RECT 0.795 0.975 0.865 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.33 0.085 ;
        RECT 1.175 -0.085 1.245 0.425 ;
        RECT 0.795 -0.085 0.865 0.285 ;
        RECT 0.415 -0.085 0.485 0.285 ;
        RECT 0.04 -0.085 0.11 0.425 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.84 0.115 1.25 ;
      RECT 0.045 0.84 0.925 0.91 ;
      RECT 0.855 0.355 0.925 0.91 ;
      RECT 0.235 0.355 0.925 0.425 ;
      RECT 0.605 0.15 0.675 0.425 ;
      RECT 0.235 0.15 0.305 0.425 ;
  END
END OR4_X2

MACRO OR4_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4_X4 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.805 0.525 0.89 0.7 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.01 0.39 1.14 0.66 ;
        RECT 0.505 0.39 1.14 0.46 ;
        RECT 0.505 0.39 0.575 0.66 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.31 0.77 1.33 0.84 ;
        RECT 1.26 0.525 1.33 0.84 ;
        RECT 0.31 0.525 0.38 0.84 ;
        RECT 0.25 0.525 0.38 0.7 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.115 0.905 1.52 0.975 ;
        RECT 1.45 0.525 1.52 0.975 ;
        RECT 0.115 0.525 0.185 0.975 ;
        RECT 0.06 0.525 0.185 0.7 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.13 0.15 2.2 1.25 ;
        RECT 1.755 0.56 2.2 0.7 ;
        RECT 1.755 0.15 1.825 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.47 1.485 ;
        RECT 2.315 1.045 2.385 1.485 ;
        RECT 1.935 1.045 2.005 1.485 ;
        RECT 1.555 1.205 1.625 1.485 ;
        RECT 0.04 1.045 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.47 0.085 ;
        RECT 2.315 -0.085 2.385 0.4 ;
        RECT 1.905 -0.085 2.04 0.365 ;
        RECT 1.525 -0.085 1.66 0.325 ;
        RECT 1.145 -0.085 1.28 0.16 ;
        RECT 0.765 -0.085 0.9 0.16 ;
        RECT 0.385 -0.085 0.52 0.16 ;
        RECT 0.04 -0.085 0.11 0.4 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.77 1.04 1.685 1.11 ;
      RECT 1.615 0.39 1.685 1.11 ;
      RECT 1.37 0.39 1.685 0.46 ;
      RECT 0.235 0.15 0.305 0.425 ;
      RECT 1.37 0.15 1.44 0.46 ;
      RECT 0.235 0.225 1.44 0.295 ;
  END
END OR4_X4

MACRO SDFFRS_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRS_X1 0 0 ;
  SIZE 5.51 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 5.07 0.765 5.26 0.98 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.82 0.525 0.92 0.7 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 5.19 0.39 5.335 0.56 ;
        RECT 4.76 0.39 5.335 0.46 ;
        RECT 4.76 0.765 5.005 0.835 ;
        RECT 4.76 0.39 4.83 0.835 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.56 0.695 4.69 0.84 ;
    END
  END SI
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.01 0.525 1.11 0.7 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.575 0.7 1.67 0.84 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.26 0.13 1.105 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425 0.36 0.51 0.8 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 5.51 1.485 ;
        RECT 5.175 1.095 5.31 1.485 ;
        RECT 4.415 1.13 4.55 1.485 ;
        RECT 3.585 1.03 3.72 1.485 ;
        RECT 3.045 0.865 3.18 1.485 ;
        RECT 2.665 0.99 2.8 1.485 ;
        RECT 1.945 0.83 2.015 1.485 ;
        RECT 1.305 1.105 1.44 1.485 ;
        RECT 0.925 1.105 1.06 1.485 ;
        RECT 0.545 1.035 0.68 1.485 ;
        RECT 0.195 1.18 0.33 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 5.51 0.085 ;
        RECT 5.175 -0.085 5.31 0.225 ;
        RECT 4.415 -0.085 4.55 0.225 ;
        RECT 3.4 -0.085 3.535 0.285 ;
        RECT 2.665 -0.085 2.8 0.285 ;
        RECT 1.755 -0.085 1.825 0.32 ;
        RECT 0.92 -0.085 1.055 0.285 ;
        RECT 0.195 -0.085 0.33 0.16 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 5.4 0.215 5.47 1.235 ;
      RECT 4.9 0.625 5.47 0.695 ;
      RECT 4.9 0.56 4.975 0.695 ;
      RECT 4.37 0.945 4.93 1.015 ;
      RECT 4.37 0.41 4.44 1.015 ;
      RECT 4.37 0.41 4.685 0.48 ;
      RECT 4.615 0.22 4.685 0.48 ;
      RECT 4.615 0.22 4.93 0.29 ;
      RECT 3.94 1.18 4.28 1.25 ;
      RECT 4.21 0.16 4.28 1.25 ;
      RECT 3.94 0.76 4.01 1.25 ;
      RECT 2.18 1.035 2.525 1.105 ;
      RECT 2.455 0.35 2.525 1.105 ;
      RECT 3.27 0.76 3.34 1.09 ;
      RECT 3.27 0.76 4.01 0.83 ;
      RECT 3.865 0.16 3.935 0.51 ;
      RECT 3.265 0.35 3.935 0.42 ;
      RECT 2.455 0.35 2.98 0.42 ;
      RECT 2.91 0.16 2.98 0.42 ;
      RECT 3.265 0.16 3.335 0.42 ;
      RECT 3.865 0.16 4.28 0.23 ;
      RECT 2.91 0.16 3.335 0.23 ;
      RECT 4.075 0.295 4.145 1.115 ;
      RECT 2.75 0.62 4.145 0.69 ;
      RECT 4 0.295 4.145 0.69 ;
      RECT 3.805 0.895 3.875 1.115 ;
      RECT 3.435 0.895 3.505 1.115 ;
      RECT 3.435 0.895 3.875 0.965 ;
      RECT 2.615 0.755 2.99 0.825 ;
      RECT 2.615 0.485 2.685 0.825 ;
      RECT 2.615 0.485 3.8 0.555 ;
      RECT 3.045 0.295 3.18 0.555 ;
      RECT 2.315 0.2 2.385 0.965 ;
      RECT 1.415 0.555 2.385 0.625 ;
      RECT 2.125 0.695 2.195 0.965 ;
      RECT 1.755 0.695 1.825 0.965 ;
      RECT 1.755 0.695 2.195 0.765 ;
      RECT 1.145 0.765 1.215 1.105 ;
      RECT 0.61 0.765 1.215 0.835 ;
      RECT 0.61 0.39 0.68 0.835 ;
      RECT 0.61 0.39 1.19 0.46 ;
      RECT 1.12 0.25 1.19 0.46 ;
      RECT 1.62 0.385 2.15 0.455 ;
      RECT 1.62 0.15 1.69 0.455 ;
      RECT 1.12 0.25 1.4 0.32 ;
      RECT 1.33 0.15 1.4 0.32 ;
      RECT 1.33 0.15 1.69 0.22 ;
      RECT 1.585 1.165 1.815 1.235 ;
      RECT 1.585 0.905 1.655 1.235 ;
      RECT 1.28 0.905 1.655 0.975 ;
      RECT 1.28 0.41 1.35 0.975 ;
      RECT 1.28 0.41 1.555 0.48 ;
      RECT 1.485 0.285 1.555 0.48 ;
      RECT 0.195 0.9 0.865 0.97 ;
      RECT 0.195 0.225 0.265 0.97 ;
      RECT 0.195 0.225 0.68 0.295 ;
  END
END SDFFRS_X1

MACRO SDFFRS_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRS_X2 0 0 ;
  SIZE 5.89 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 5.495 0.42 5.64 0.56 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.01 0.545 1.165 0.7 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 5.57 0.675 5.7 0.84 ;
        RECT 5.135 0.72 5.7 0.79 ;
        RECT 5.135 0.385 5.205 0.79 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.925 0.56 5.07 0.7 ;
    END
  END SI
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.365 0.545 1.46 0.7 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.9 0.175 2.065 0.245 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.24 0.15 0.32 1.125 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6 0.435 0.735 0.9 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 5.89 1.485 ;
        RECT 5.54 1.195 5.675 1.485 ;
        RECT 4.78 1.09 4.915 1.485 ;
        RECT 3.95 1.09 4.085 1.485 ;
        RECT 3.42 0.985 3.555 1.485 ;
        RECT 3.04 0.985 3.175 1.485 ;
        RECT 2.285 0.965 2.42 1.485 ;
        RECT 1.64 1.115 1.775 1.485 ;
        RECT 1.18 1.12 1.315 1.485 ;
        RECT 0.79 1.1 0.925 1.485 ;
        RECT 0.41 1.1 0.545 1.485 ;
        RECT 0.065 0.85 0.135 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 5.89 0.085 ;
        RECT 5.54 -0.085 5.675 0.18 ;
        RECT 4.81 -0.085 4.88 0.27 ;
        RECT 3.76 -0.085 3.895 0.285 ;
        RECT 3.04 -0.085 3.175 0.285 ;
        RECT 2.13 -0.085 2.2 0.32 ;
        RECT 1.7 -0.085 1.835 0.285 ;
        RECT 0.79 -0.085 0.925 0.16 ;
        RECT 0.41 -0.085 0.545 0.16 ;
        RECT 0.065 -0.085 0.135 0.41 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 5.765 0.15 5.835 1.09 ;
      RECT 5.27 0.565 5.41 0.635 ;
      RECT 5.34 0.285 5.41 0.635 ;
      RECT 5.34 0.285 5.835 0.355 ;
      RECT 4.74 0.95 5.295 1.02 ;
      RECT 4.74 0.375 4.81 1.02 ;
      RECT 4.74 0.375 5.045 0.445 ;
      RECT 4.975 0.165 5.045 0.445 ;
      RECT 4.975 0.165 5.295 0.235 ;
      RECT 4.305 1.155 4.675 1.225 ;
      RECT 4.605 0.15 4.675 1.225 ;
      RECT 2.555 1.115 2.915 1.185 ;
      RECT 2.845 0.35 2.915 1.185 ;
      RECT 4.305 0.765 4.375 1.225 ;
      RECT 3.615 0.765 4.375 0.835 ;
      RECT 4.575 0.69 4.675 0.825 ;
      RECT 3.61 0.355 4.34 0.425 ;
      RECT 4.27 0.15 4.34 0.425 ;
      RECT 2.845 0.35 3.39 0.42 ;
      RECT 3.32 0.15 3.39 0.42 ;
      RECT 3.61 0.15 3.68 0.425 ;
      RECT 4.27 0.15 4.675 0.22 ;
      RECT 3.32 0.15 3.68 0.22 ;
      RECT 4.44 0.625 4.51 1.09 ;
      RECT 3.125 0.625 4.51 0.695 ;
      RECT 4.405 0.285 4.475 0.695 ;
      RECT 4.405 0.285 4.54 0.355 ;
      RECT 4.17 0.955 4.24 1.175 ;
      RECT 3.8 0.955 3.87 1.175 ;
      RECT 3.8 0.955 4.24 1.025 ;
      RECT 2.99 0.765 3.37 0.835 ;
      RECT 2.99 0.485 3.06 0.835 ;
      RECT 2.99 0.49 4.17 0.56 ;
      RECT 2.99 0.485 3.525 0.56 ;
      RECT 3.455 0.32 3.525 0.56 ;
      RECT 2.7 0.2 2.77 1.05 ;
      RECT 1.665 0.485 1.735 0.68 ;
      RECT 1.665 0.485 2.77 0.555 ;
      RECT 1.53 0.84 2.04 0.91 ;
      RECT 1.97 0.685 2.04 0.91 ;
      RECT 1.53 0.35 1.6 0.91 ;
      RECT 1.97 0.685 2.635 0.755 ;
      RECT 2.565 0.62 2.635 0.755 ;
      RECT 1.53 0.35 2.04 0.42 ;
      RECT 2.5 0.83 2.57 1.05 ;
      RECT 2.13 0.83 2.2 1.05 ;
      RECT 2.13 0.83 2.57 0.9 ;
      RECT 1.84 1.16 2.22 1.23 ;
      RECT 1.84 0.975 1.91 1.23 ;
      RECT 1.395 0.975 1.91 1.045 ;
      RECT 1.395 0.765 1.465 1.045 ;
      RECT 0.87 0.765 1.465 0.835 ;
      RECT 0.87 0.41 0.94 0.835 ;
      RECT 0.87 0.41 1.46 0.48 ;
      RECT 0.39 0.965 1.12 1.035 ;
      RECT 0.39 0.23 0.46 1.035 ;
      RECT 0.39 0.23 1.305 0.3 ;
  END
END SDFFRS_X2

MACRO SDFFR_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFR_X1 0 0 ;
  SIZE 4.75 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.24 0.56 4.365 0.7 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.82 0.84 0.925 0.98 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.105 0.77 4.53 0.84 ;
        RECT 4.43 0.56 4.53 0.84 ;
        RECT 4.105 0.565 4.175 0.84 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.67 0.655 3.765 0.84 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.77 0.66 1.995 0.84 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.435 0.185 0.51 1.015 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.185 0.13 1.065 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 4.75 1.485 ;
        RECT 4.4 1.045 4.47 1.485 ;
        RECT 3.64 1.08 3.71 1.485 ;
        RECT 3.27 1.08 3.34 1.485 ;
        RECT 2.4 0.995 2.47 1.485 ;
        RECT 1.84 1.06 1.975 1.485 ;
        RECT 1.15 1.205 1.22 1.485 ;
        RECT 0.74 1.24 0.875 1.485 ;
        RECT 0.21 1.24 0.345 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 4.75 0.085 ;
        RECT 4.4 -0.085 4.47 0.32 ;
        RECT 3.64 -0.085 3.71 0.32 ;
        RECT 3.11 -0.085 3.18 0.32 ;
        RECT 2.27 -0.085 2.34 0.425 ;
        RECT 1.71 -0.085 1.845 0.285 ;
        RECT 0.77 -0.085 0.84 0.32 ;
        RECT 0.24 -0.085 0.31 0.46 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 4.595 0.185 4.665 1.22 ;
      RECT 3.965 0.905 4.665 0.975 ;
      RECT 3.965 0.715 4.035 0.975 ;
      RECT 4.1 0.415 4.665 0.485 ;
      RECT 3.83 1.04 4.125 1.11 ;
      RECT 3.83 0.22 3.9 1.11 ;
      RECT 3.12 0.52 3.9 0.59 ;
      RECT 3.83 0.22 4.125 0.29 ;
      RECT 2.54 1.18 3.205 1.25 ;
      RECT 3.135 0.945 3.205 1.25 ;
      RECT 3.45 0.945 3.52 1.2 ;
      RECT 2.54 0.505 2.61 1.25 ;
      RECT 3.135 0.945 3.585 1.015 ;
      RECT 3.515 0.655 3.585 1.015 ;
      RECT 2.985 0.655 3.585 0.725 ;
      RECT 2.985 0.385 3.055 0.725 ;
      RECT 2.985 0.385 3.335 0.455 ;
      RECT 3.265 0.185 3.335 0.455 ;
      RECT 2.69 1.015 3.065 1.085 ;
      RECT 2.995 0.81 3.065 1.085 ;
      RECT 2.69 0.305 2.76 1.085 ;
      RECT 2.995 0.81 3.45 0.88 ;
      RECT 2.22 0.855 2.29 1.13 ;
      RECT 2.22 0.855 2.405 0.925 ;
      RECT 2.335 0.49 2.405 0.925 ;
      RECT 2.85 0.17 2.92 0.835 ;
      RECT 1.43 0.49 1.5 0.7 ;
      RECT 1.43 0.49 2.475 0.56 ;
      RECT 2.405 0.17 2.475 0.56 ;
      RECT 2.09 0.185 2.16 0.56 ;
      RECT 2.405 0.17 2.92 0.24 ;
      RECT 1.545 1.18 1.695 1.25 ;
      RECT 1.625 0.765 1.695 1.25 ;
      RECT 2.065 0.655 2.135 1.065 ;
      RECT 1.625 0.905 2.135 0.975 ;
      RECT 1.28 0.765 1.695 0.835 ;
      RECT 2.065 0.655 2.26 0.79 ;
      RECT 1.28 0.35 1.35 0.835 ;
      RECT 1.28 0.35 2 0.42 ;
      RECT 1.93 0.185 2 0.42 ;
      RECT 1.49 0.905 1.56 1.04 ;
      RECT 1.14 0.905 1.56 0.975 ;
      RECT 1.14 0.215 1.21 0.975 ;
      RECT 0.72 0.705 1.21 0.775 ;
      RECT 0.72 0.525 0.79 0.775 ;
      RECT 1.14 0.215 1.46 0.285 ;
      RECT 0.585 0.185 0.655 1.24 ;
      RECT 0.195 1.08 0.655 1.15 ;
      RECT 0.195 0.525 0.265 1.15 ;
      RECT 1.005 0.39 1.075 0.635 ;
      RECT 0.585 0.39 1.075 0.46 ;
      RECT 0.935 1.045 1.41 1.115 ;
  END
END SDFFR_X1

MACRO SDFFR_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFR_X2 0 0 ;
  SIZE 4.94 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.565 0.42 4.69 0.625 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.145 0.84 1.27 0.98 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.345 0.7 4.765 0.845 ;
        RECT 4.345 0.565 4.415 0.845 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.86 0.67 4.005 0.84 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.145 0.695 2.28 0.84 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425 0.395 0.51 1.005 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.795 0.56 0.89 1.005 ;
        RECT 0.795 0.395 0.865 1.005 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 4.94 1.485 ;
        RECT 4.635 1.045 4.705 1.485 ;
        RECT 3.875 1.08 3.945 1.485 ;
        RECT 3.46 1.115 3.595 1.485 ;
        RECT 2.66 0.995 2.73 1.485 ;
        RECT 2.06 1.06 2.195 1.485 ;
        RECT 1.37 1.205 1.44 1.485 ;
        RECT 0.985 1.205 1.055 1.485 ;
        RECT 0.575 1.24 0.71 1.485 ;
        RECT 0.225 1.205 0.295 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 4.94 0.085 ;
        RECT 4.635 -0.085 4.705 0.195 ;
        RECT 3.875 -0.085 3.945 0.32 ;
        RECT 3.295 -0.085 3.365 0.32 ;
        RECT 2.535 -0.085 2.605 0.42 ;
        RECT 2.005 -0.085 2.075 0.32 ;
        RECT 1.065 -0.085 1.135 0.32 ;
        RECT 0.575 -0.085 0.71 0.16 ;
        RECT 0.195 -0.085 0.33 0.16 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 4.83 0.195 4.9 1.22 ;
      RECT 4.205 0.91 4.9 0.98 ;
      RECT 4.205 0.715 4.275 0.98 ;
      RECT 4.36 0.415 4.495 0.485 ;
      RECT 4.425 0.285 4.495 0.485 ;
      RECT 4.425 0.285 4.9 0.355 ;
      RECT 4.07 1.045 4.36 1.115 ;
      RECT 4.07 0.23 4.14 1.115 ;
      RECT 3.42 0.52 4.14 0.59 ;
      RECT 4.07 0.23 4.36 0.3 ;
      RECT 2.805 1.18 3.255 1.25 ;
      RECT 3.185 0.975 3.255 1.25 ;
      RECT 3.69 0.655 3.76 1.2 ;
      RECT 2.805 0.5 2.875 1.25 ;
      RECT 3.185 0.975 3.76 1.045 ;
      RECT 3.285 0.655 3.76 0.725 ;
      RECT 3.285 0.385 3.355 0.725 ;
      RECT 3.285 0.385 3.57 0.455 ;
      RECT 3.5 0.2 3.57 0.455 ;
      RECT 3.04 0.84 3.11 1.115 ;
      RECT 2.955 0.84 3.11 0.915 ;
      RECT 2.955 0.84 3.625 0.91 ;
      RECT 2.955 0.33 3.025 0.915 ;
      RECT 2.89 0.33 3.025 0.4 ;
      RECT 2.48 0.815 2.55 1.09 ;
      RECT 2.48 0.815 2.74 0.885 ;
      RECT 2.67 0.165 2.74 0.885 ;
      RECT 3.15 0.165 3.22 0.775 ;
      RECT 1.715 0.545 1.785 0.685 ;
      RECT 1.715 0.545 2.74 0.615 ;
      RECT 2.35 0.285 2.42 0.615 ;
      RECT 2.67 0.165 3.22 0.235 ;
      RECT 1.79 1.18 1.95 1.25 ;
      RECT 1.88 0.75 1.95 1.25 ;
      RECT 1.88 0.915 2.415 0.985 ;
      RECT 2.345 0.68 2.415 0.985 ;
      RECT 1.56 0.75 1.95 0.82 ;
      RECT 2.345 0.68 2.56 0.75 ;
      RECT 1.56 0.41 1.63 0.82 ;
      RECT 1.56 0.41 2.265 0.48 ;
      RECT 2.195 0.26 2.265 0.48 ;
      RECT 1.425 0.885 1.815 0.955 ;
      RECT 1.425 0.265 1.495 0.955 ;
      RECT 0.29 0.26 0.36 0.66 ;
      RECT 0.93 0.385 1.495 0.455 ;
      RECT 0.93 0.26 1 0.455 ;
      RECT 1.425 0.265 1.73 0.335 ;
      RECT 0.29 0.26 1 0.33 ;
      RECT 1.155 1.045 1.29 1.25 ;
      RECT 1.155 1.045 1.63 1.115 ;
      RECT 0.045 1.07 1.08 1.14 ;
      RECT 1.01 0.64 1.08 1.14 ;
      RECT 0.66 0.525 0.73 1.14 ;
      RECT 0.045 0.26 0.115 1.14 ;
      RECT 1.01 0.64 1.36 0.775 ;
  END
END SDFFR_X2

MACRO SDFFS_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFS_X1 0 0 ;
  SIZE 4.75 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.55 0.38 0.7 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.765 0.57 0.835 ;
        RECT 0.5 0.55 0.57 0.835 ;
        RECT 0.06 0.55 0.185 0.835 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.91 0.42 1.08 0.56 ;
    END
  END SI
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.84 0.42 3.93 0.575 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.01 0.785 1.115 0.98 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.24 0.98 4.335 1.25 ;
        RECT 4.265 0.4 4.335 1.25 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.62 0.98 4.705 1.25 ;
        RECT 4.635 0.15 4.705 1.25 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 4.75 1.485 ;
        RECT 4.445 0.975 4.515 1.485 ;
        RECT 4.105 0.975 4.175 1.485 ;
        RECT 3.735 1.07 3.805 1.485 ;
        RECT 2.83 1.07 2.9 1.485 ;
        RECT 2.3 1.155 2.37 1.485 ;
        RECT 1.52 1.04 1.59 1.485 ;
        RECT 0.985 1.045 1.055 1.485 ;
        RECT 0.225 1.035 0.295 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 4.75 0.085 ;
        RECT 4.445 -0.085 4.515 0.195 ;
        RECT 3.735 -0.085 3.805 0.32 ;
        RECT 2.805 -0.085 2.94 0.285 ;
        RECT 2.485 -0.085 2.555 0.37 ;
        RECT 1.49 -0.085 1.625 0.215 ;
        RECT 0.985 -0.085 1.055 0.285 ;
        RECT 0.225 -0.085 0.295 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 3.915 0.775 3.985 1.25 ;
      RECT 3.69 0.775 3.985 0.915 ;
      RECT 3.69 0.775 4.2 0.845 ;
      RECT 4.13 0.265 4.2 0.845 ;
      RECT 4.495 0.265 4.565 0.66 ;
      RECT 4.075 0.265 4.565 0.335 ;
      RECT 3.255 1.1 3.625 1.17 ;
      RECT 3.555 0.215 3.625 1.17 ;
      RECT 3.555 0.64 4.065 0.71 ;
      RECT 3.995 0.525 4.065 0.71 ;
      RECT 3.25 0.215 3.625 0.285 ;
      RECT 2.615 0.93 3.49 1 ;
      RECT 3.42 0.35 3.49 1 ;
      RECT 2.615 0.805 2.685 1 ;
      RECT 2.225 0.805 2.685 0.875 ;
      RECT 2.65 0.35 3.49 0.42 ;
      RECT 2.65 0.2 2.72 0.42 ;
      RECT 1.34 0.905 1.41 1.25 ;
      RECT 1.34 0.905 1.865 0.975 ;
      RECT 1.795 0.74 1.865 0.975 ;
      RECT 3.285 0.485 3.355 0.86 ;
      RECT 1.795 0.74 2.025 0.81 ;
      RECT 1.955 0.42 2.025 0.81 ;
      RECT 2.225 0.485 3.355 0.555 ;
      RECT 1.74 0.42 2.025 0.49 ;
      RECT 2.225 0.15 2.295 0.555 ;
      RECT 1.74 0.15 1.81 0.49 ;
      RECT 1.34 0.28 1.81 0.35 ;
      RECT 1.34 0.15 1.41 0.35 ;
      RECT 1.74 0.15 2.295 0.22 ;
      RECT 1.87 1.17 2.005 1.24 ;
      RECT 1.935 0.88 2.005 1.24 ;
      RECT 1.935 0.88 2.16 0.95 ;
      RECT 2.09 0.285 2.16 0.95 ;
      RECT 2.09 0.665 2.945 0.735 ;
      RECT 1.875 0.285 2.16 0.355 ;
      RECT 2.455 1.17 2.59 1.24 ;
      RECT 2.07 1.17 2.205 1.24 ;
      RECT 2.135 1.02 2.205 1.24 ;
      RECT 2.455 1.02 2.525 1.24 ;
      RECT 2.135 1.02 2.525 1.09 ;
      RECT 1.18 0.77 1.25 1.25 ;
      RECT 1.18 0.77 1.675 0.84 ;
      RECT 1.605 0.415 1.675 0.84 ;
      RECT 1.605 0.6 1.89 0.67 ;
      RECT 1.18 0.415 1.675 0.485 ;
      RECT 1.18 0.15 1.25 0.485 ;
      RECT 0.58 1.035 0.715 1.24 ;
      RECT 0.58 1.035 0.9 1.105 ;
      RECT 0.83 0.625 0.9 1.105 ;
      RECT 0.775 0.625 1.54 0.695 ;
      RECT 0.775 0.15 0.845 0.695 ;
      RECT 0.615 0.15 0.845 0.285 ;
      RECT 0.045 0.9 0.115 1.25 ;
      RECT 0.045 0.9 0.765 0.97 ;
      RECT 0.635 0.835 0.765 0.97 ;
      RECT 0.635 0.415 0.705 0.97 ;
      RECT 0.045 0.415 0.705 0.485 ;
      RECT 0.045 0.15 0.115 0.485 ;
  END
END SDFFS_X1

MACRO SDFFS_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFS_X2 0 0 ;
  SIZE 5.13 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.25 0.67 0.375 0.84 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.91 0.595 0.98 ;
        RECT 0.525 0.67 0.595 0.98 ;
        RECT 0.06 0.795 0.185 0.98 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.965 0.42 1.08 0.64 ;
    END
  END SI
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.34 0.56 4.03 0.63 ;
        RECT 3.34 0.28 3.41 0.63 ;
        RECT 2.91 0.28 3.41 0.35 ;
        RECT 2.42 0.425 2.98 0.495 ;
        RECT 2.91 0.28 2.98 0.495 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.01 0.84 1.13 0.98 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.43 0.395 4.5 0.785 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.81 0.395 4.88 0.785 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 5.13 1.485 ;
        RECT 4.99 1.125 5.06 1.485 ;
        RECT 4.58 1.15 4.715 1.485 ;
        RECT 4.2 1.15 4.335 1.485 ;
        RECT 3.825 1.15 3.96 1.485 ;
        RECT 3.51 1.12 3.58 1.485 ;
        RECT 2.64 1.03 2.71 1.485 ;
        RECT 2.265 1.165 2.4 1.485 ;
        RECT 1.505 1.24 1.64 1.485 ;
        RECT 0.99 1.115 1.06 1.485 ;
        RECT 0.195 1.24 0.33 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 5.13 0.085 ;
        RECT 4.99 -0.085 5.06 0.195 ;
        RECT 4.58 -0.085 4.715 0.18 ;
        RECT 4.2 -0.085 4.335 0.18 ;
        RECT 3.475 -0.085 3.61 0.48 ;
        RECT 2.475 -0.085 2.61 0.345 ;
        RECT 1.51 -0.085 1.645 0.345 ;
        RECT 0.96 -0.085 1.095 0.28 ;
        RECT 0.2 -0.085 0.335 0.465 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 2.91 1.18 3.445 1.25 ;
      RECT 3.375 0.985 3.445 1.25 ;
      RECT 2.91 0.83 2.98 1.25 ;
      RECT 3.375 0.985 5.015 1.055 ;
      RECT 4.945 0.26 5.015 1.055 ;
      RECT 2.26 0.83 2.98 0.965 ;
      RECT 3.69 0.26 3.76 0.495 ;
      RECT 3.69 0.26 5.015 0.33 ;
      RECT 3.375 0.85 4.745 0.92 ;
      RECT 4.675 0.525 4.745 0.92 ;
      RECT 4.295 0.415 4.365 0.92 ;
      RECT 3.825 0.415 4.365 0.485 ;
      RECT 3.045 1.045 3.31 1.115 ;
      RECT 3.24 0.695 3.31 1.115 ;
      RECT 3.24 0.695 4.23 0.765 ;
      RECT 4.095 0.56 4.23 0.765 ;
      RECT 3.205 0.415 3.275 0.76 ;
      RECT 3.045 0.415 3.275 0.485 ;
      RECT 1.355 1.105 1.425 1.25 ;
      RECT 1.355 1.105 1.855 1.175 ;
      RECT 1.785 0.76 1.855 1.175 ;
      RECT 3.07 0.845 3.175 0.98 ;
      RECT 3.07 0.56 3.14 0.98 ;
      RECT 1.785 0.76 2.05 0.83 ;
      RECT 1.98 0.425 2.05 0.83 ;
      RECT 2.285 0.56 3.14 0.63 ;
      RECT 1.98 0.425 2.075 0.575 ;
      RECT 2.285 0.155 2.355 0.63 ;
      RECT 1.355 0.425 2.075 0.495 ;
      RECT 1.75 0.155 1.82 0.495 ;
      RECT 1.355 0.36 1.425 0.495 ;
      RECT 1.75 0.155 2.355 0.225 ;
      RECT 1.925 0.895 1.995 1.25 ;
      RECT 1.925 0.895 2.195 0.965 ;
      RECT 2.125 0.695 2.195 0.965 ;
      RECT 2.125 0.695 2.825 0.765 ;
      RECT 2.15 0.29 2.22 0.765 ;
      RECT 1.895 0.29 2.22 0.36 ;
      RECT 2.485 1.03 2.555 1.25 ;
      RECT 2.115 1.03 2.185 1.25 ;
      RECT 2.115 1.03 2.555 1.1 ;
      RECT 1.195 0.87 1.265 1.25 ;
      RECT 1.195 0.87 1.705 0.94 ;
      RECT 1.635 0.56 1.705 0.94 ;
      RECT 1.635 0.625 1.915 0.695 ;
      RECT 1.195 0.56 1.705 0.63 ;
      RECT 1.195 0.315 1.265 0.63 ;
      RECT 0.585 1.18 0.9 1.25 ;
      RECT 0.83 0.35 0.9 1.25 ;
      RECT 0.83 0.705 1.57 0.775 ;
      RECT 0.585 0.35 0.9 0.42 ;
      RECT 0.045 1.045 0.115 1.25 ;
      RECT 0.045 1.045 0.765 1.115 ;
      RECT 0.695 0.535 0.765 1.115 ;
      RECT 0.045 0.535 0.765 0.605 ;
      RECT 0.045 0.38 0.115 0.605 ;
  END
END SDFFS_X2

MACRO SDFF_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFF_X1 0 0 ;
  SIZE 4.37 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.975 0.42 4.125 0.565 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.05 0.7 4.18 0.84 ;
        RECT 3.75 0.7 4.18 0.77 ;
        RECT 3.75 0.59 3.885 0.77 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.415 0.525 3.55 0.7 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.02 0.42 2.225 0.58 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.44 0.15 0.51 0.785 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.15 0.135 1.215 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 4.37 1.485 ;
        RECT 4.02 0.975 4.155 1.485 ;
        RECT 3.295 1.04 3.365 1.485 ;
        RECT 2.935 1.08 3.005 1.485 ;
        RECT 2.07 0.94 2.14 1.485 ;
        RECT 1.51 0.975 1.645 1.485 ;
        RECT 0.75 1.165 0.885 1.485 ;
        RECT 0.25 1.04 0.32 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 4.37 0.085 ;
        RECT 4.02 -0.085 4.155 0.16 ;
        RECT 3.295 -0.085 3.365 0.195 ;
        RECT 2.905 -0.085 3.04 0.19 ;
        RECT 2.04 -0.085 2.175 0.285 ;
        RECT 1.51 -0.085 1.645 0.285 ;
        RECT 0.75 -0.085 0.885 0.285 ;
        RECT 0.25 -0.085 0.32 0.425 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 4.245 0.15 4.315 1.215 ;
      RECT 3.615 0.45 3.685 0.84 ;
      RECT 3.615 0.45 3.88 0.52 ;
      RECT 3.81 0.28 3.88 0.52 ;
      RECT 3.81 0.28 4.315 0.35 ;
      RECT 3.67 0.905 3.74 1.215 ;
      RECT 3.28 0.905 3.74 0.975 ;
      RECT 3.28 0.285 3.35 0.975 ;
      RECT 2.9 0.695 3.35 0.83 ;
      RECT 3.28 0.285 3.74 0.355 ;
      RECT 3.67 0.15 3.74 0.355 ;
      RECT 3.125 0.92 3.195 1.215 ;
      RECT 2.205 1.14 2.835 1.21 ;
      RECT 2.765 0.545 2.835 1.21 ;
      RECT 2.205 0.815 2.275 1.21 ;
      RECT 2.765 0.92 3.195 0.99 ;
      RECT 2.765 0.545 3.215 0.615 ;
      RECT 3.145 0.15 3.215 0.615 ;
      RECT 2.53 0.975 2.7 1.045 ;
      RECT 2.63 0.215 2.7 1.045 ;
      RECT 2.63 0.325 3.08 0.46 ;
      RECT 2.53 0.215 2.7 0.285 ;
      RECT 1.885 0.2 1.955 1.09 ;
      RECT 2.37 0.68 2.44 0.95 ;
      RECT 1.885 0.68 2.565 0.75 ;
      RECT 2.495 0.35 2.565 0.75 ;
      RECT 1.26 0.65 1.955 0.72 ;
      RECT 1.73 0.84 1.8 1.215 ;
      RECT 1.125 0.84 1.8 0.91 ;
      RECT 1.125 0.475 1.195 0.91 ;
      RECT 1.125 0.475 1.8 0.545 ;
      RECT 1.73 0.32 1.8 0.545 ;
      RECT 0.99 1.15 1.265 1.22 ;
      RECT 0.99 0.23 1.06 1.22 ;
      RECT 0.73 0.525 1.06 0.66 ;
      RECT 0.99 0.23 1.265 0.3 ;
      RECT 0.595 0.15 0.665 1.215 ;
      RECT 0.2 0.885 0.665 0.955 ;
      RECT 0.2 0.51 0.27 0.955 ;
      RECT 0.595 0.73 0.925 0.865 ;
  END
END SDFF_X1

MACRO SDFF_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFF_X2 0 0 ;
  SIZE 4.56 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.165 0.42 4.33 0.56 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.95 0.7 4.355 0.84 ;
        RECT 3.95 0.595 4.02 0.84 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.48 0.42 3.58 0.56 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.225 0.42 2.41 0.58 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425 0.4 0.51 0.785 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.805 0.185 0.89 0.84 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 4.56 1.485 ;
        RECT 4.24 0.965 4.31 1.485 ;
        RECT 3.455 1.24 3.59 1.485 ;
        RECT 3.135 1.08 3.205 1.485 ;
        RECT 2.275 0.91 2.345 1.485 ;
        RECT 1.745 0.94 1.815 1.485 ;
        RECT 0.985 1.04 1.055 1.485 ;
        RECT 0.605 1.04 0.675 1.485 ;
        RECT 0.225 1.04 0.295 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 4.56 0.085 ;
        RECT 4.21 -0.085 4.345 0.16 ;
        RECT 3.485 -0.085 3.555 0.255 ;
        RECT 3.065 -0.085 3.2 0.165 ;
        RECT 2.275 -0.085 2.345 0.32 ;
        RECT 1.745 -0.085 1.815 0.32 ;
        RECT 0.985 -0.085 1.055 0.32 ;
        RECT 0.605 -0.085 0.675 0.195 ;
        RECT 0.225 -0.085 0.295 0.195 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 4.43 0.195 4.5 1.24 ;
      RECT 3.78 0.42 3.85 0.895 ;
      RECT 3.78 0.42 4.05 0.49 ;
      RECT 3.98 0.285 4.05 0.49 ;
      RECT 3.98 0.285 4.5 0.355 ;
      RECT 3.86 0.96 3.93 1.24 ;
      RECT 3.645 0.96 3.93 1.03 ;
      RECT 3.645 0.15 3.715 1.03 ;
      RECT 3.105 0.64 3.715 0.775 ;
      RECT 3.645 0.15 3.965 0.22 ;
      RECT 3.33 0.89 3.4 1.185 ;
      RECT 2.41 1.11 3.04 1.18 ;
      RECT 2.97 0.505 3.04 1.18 ;
      RECT 2.41 0.785 2.48 1.18 ;
      RECT 2.97 0.89 3.4 0.96 ;
      RECT 2.97 0.505 3.405 0.575 ;
      RECT 3.335 0.185 3.405 0.575 ;
      RECT 2.63 0.945 2.905 1.015 ;
      RECT 2.835 0.215 2.905 1.015 ;
      RECT 2.835 0.37 3.27 0.44 ;
      RECT 2.635 0.215 2.905 0.285 ;
      RECT 2.09 0.185 2.16 1.185 ;
      RECT 2.575 0.65 2.645 0.88 ;
      RECT 2.09 0.65 2.77 0.72 ;
      RECT 2.7 0.35 2.77 0.72 ;
      RECT 1.42 0.63 2.16 0.7 ;
      RECT 1.935 0.79 2.005 1.185 ;
      RECT 1.265 0.475 1.335 0.985 ;
      RECT 1.265 0.79 2.005 0.86 ;
      RECT 1.265 0.475 2.005 0.545 ;
      RECT 1.935 0.185 2.005 0.545 ;
      RECT 1.13 1.055 1.47 1.125 ;
      RECT 1.13 0.22 1.2 1.125 ;
      RECT 0.29 0.905 1.2 0.975 ;
      RECT 0.29 0.525 0.36 0.975 ;
      RECT 1.13 0.22 1.47 0.29 ;
      RECT 0.045 0.185 0.115 1.185 ;
      RECT 0.67 0.265 0.74 0.66 ;
      RECT 0.045 0.265 0.74 0.335 ;
  END
END SDFF_X2

MACRO TBUF_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUF_X1 0 0 ;
  SIZE 1.52 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.82 0.495 0.89 0.73 ;
        RECT 0.51 0.495 0.89 0.565 ;
        RECT 0.51 0.495 0.58 0.63 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.2 0.695 1.33 0.92 ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.035 0.97 0.14 1.245 ;
        RECT 0.035 0.15 0.14 0.425 ;
        RECT 0.035 0.15 0.105 1.245 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.52 1.485 ;
        RECT 1.19 1.24 1.325 1.485 ;
        RECT 0.69 1.145 0.76 1.485 ;
        RECT 0.225 1.145 0.36 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.52 0.085 ;
        RECT 1.15 -0.085 1.285 0.295 ;
        RECT 0.77 -0.085 0.905 0.295 ;
        RECT 0.225 -0.085 0.36 0.16 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.41 0.365 1.48 1.245 ;
      RECT 0.875 1.105 1.48 1.175 ;
      RECT 0.875 0.94 0.945 1.175 ;
      RECT 0.65 0.94 0.945 1.01 ;
      RECT 0.65 0.645 0.72 1.01 ;
      RECT 1.345 0.365 1.48 0.435 ;
      RECT 1.065 0.36 1.135 1.04 ;
      RECT 0.17 0.495 0.305 0.565 ;
      RECT 0.235 0.225 0.305 0.565 ;
      RECT 0.615 0.36 1.135 0.43 ;
      RECT 0.615 0.225 0.685 0.43 ;
      RECT 0.235 0.225 0.685 0.295 ;
      RECT 0.495 0.835 0.565 1.115 ;
      RECT 0.37 0.835 0.565 0.905 ;
      RECT 0.37 0.36 0.44 0.905 ;
      RECT 0.17 0.645 0.44 0.715 ;
      RECT 0.37 0.36 0.53 0.43 ;
  END
END TBUF_X1

MACRO TBUF_X16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUF_X16 0 0 ;
  SIZE 4.94 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.265 0.39 4.335 0.66 ;
        RECT 3.67 0.39 4.335 0.46 ;
        RECT 3.475 0.555 3.74 0.625 ;
        RECT 3.67 0.39 3.74 0.625 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.05 0.725 4.6 0.795 ;
        RECT 4.53 0.525 4.6 0.795 ;
        RECT 4.05 0.56 4.12 0.795 ;
        RECT 3.955 0.56 4.12 0.63 ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.895 0.36 3.03 1.005 ;
        RECT 0.36 0.56 3.03 0.7 ;
        RECT 2.515 0.36 2.65 1.005 ;
        RECT 2.14 0.56 2.275 1.005 ;
        RECT 2.135 0.36 2.27 0.7 ;
        RECT 1.76 0.36 1.895 0.7 ;
        RECT 1.755 0.56 1.89 1.005 ;
        RECT 1.38 0.56 1.515 1.005 ;
        RECT 1.375 0.36 1.51 0.7 ;
        RECT 1 0.36 1.135 0.7 ;
        RECT 0.995 0.56 1.13 1.005 ;
        RECT 0.62 0.36 0.755 1.005 ;
        RECT 0.24 0.86 0.43 0.93 ;
        RECT 0.36 0.36 0.43 0.93 ;
        RECT 0.24 0.36 0.43 0.43 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 4.94 1.485 ;
        RECT 4.605 1.24 4.74 1.485 ;
        RECT 3.845 1.24 3.98 1.485 ;
        RECT 3.465 1.24 3.6 1.485 ;
        RECT 3.085 1.24 3.22 1.485 ;
        RECT 2.705 1.24 2.84 1.485 ;
        RECT 2.325 1.24 2.46 1.485 ;
        RECT 1.945 1.24 2.08 1.485 ;
        RECT 1.565 1.24 1.7 1.485 ;
        RECT 1.185 1.24 1.32 1.485 ;
        RECT 0.805 1.24 0.94 1.485 ;
        RECT 0.425 1.24 0.56 1.485 ;
        RECT 0.05 1.24 0.185 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 4.94 0.085 ;
        RECT 4.605 -0.085 4.74 0.16 ;
        RECT 4.225 -0.085 4.36 0.16 ;
        RECT 3.845 -0.085 3.98 0.16 ;
        RECT 3.085 -0.085 3.22 0.16 ;
        RECT 2.705 -0.085 2.84 0.16 ;
        RECT 2.325 -0.085 2.46 0.16 ;
        RECT 1.945 -0.085 2.08 0.16 ;
        RECT 1.565 -0.085 1.7 0.16 ;
        RECT 1.185 -0.085 1.32 0.16 ;
        RECT 0.805 -0.085 0.94 0.16 ;
        RECT 0.425 -0.085 0.56 0.16 ;
        RECT 0.05 -0.085 0.185 0.16 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 4.825 0.26 4.895 1.25 ;
      RECT 3.86 0.995 4.895 1.065 ;
      RECT 3.86 0.83 3.93 1.065 ;
      RECT 3.23 0.83 3.93 0.9 ;
      RECT 3.805 0.525 3.875 0.9 ;
      RECT 3.23 0.525 3.3 0.9 ;
      RECT 4.23 0.86 4.735 0.93 ;
      RECT 4.665 0.225 4.735 0.93 ;
      RECT 0.105 0.495 0.29 0.565 ;
      RECT 0.105 0.225 0.175 0.565 ;
      RECT 0.105 0.225 4.735 0.295 ;
      RECT 0.105 1.085 3.79 1.155 ;
      RECT 3.095 0.36 3.165 1.155 ;
      RECT 0.105 0.65 0.175 1.155 ;
      RECT 0.105 0.65 0.295 0.72 ;
      RECT 3.095 0.36 3.6 0.43 ;
  END
END TBUF_X16

MACRO TBUF_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUF_X2 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.82 0.56 0.965 0.7 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.2 0.7 1.535 0.84 ;
        RECT 1.2 0.285 1.27 0.84 ;
        RECT 0.685 0.285 1.27 0.355 ;
        RECT 0.685 0.285 0.755 0.66 ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.06 0.8 0.335 0.87 ;
        RECT 0.06 0.35 0.33 0.42 ;
        RECT 0.06 0.35 0.13 0.87 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.71 1.485 ;
        RECT 1.39 1.065 1.46 1.485 ;
        RECT 0.975 1.065 1.045 1.485 ;
        RECT 0.415 1.135 0.485 1.485 ;
        RECT 0.04 0.995 0.11 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.71 0.085 ;
        RECT 1.405 -0.085 1.475 0.25 ;
        RECT 0.91 -0.085 0.98 0.2 ;
        RECT 0.415 -0.085 0.485 0.39 ;
        RECT 0.04 -0.085 0.11 0.25 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.6 0.15 1.67 1.25 ;
      RECT 1.335 0.56 1.67 0.63 ;
      RECT 0.4 0.925 1.27 0.995 ;
      RECT 1.065 0.43 1.135 0.995 ;
      RECT 0.4 0.65 0.47 0.995 ;
      RECT 0.235 0.65 0.47 0.72 ;
      RECT 1 0.43 1.135 0.5 ;
      RECT 0.55 0.725 0.705 0.795 ;
      RECT 0.55 0.15 0.62 0.795 ;
      RECT 0.235 0.495 0.62 0.565 ;
      RECT 0.55 0.15 0.825 0.22 ;
  END
END TBUF_X2

MACRO TBUF_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUF_X4 0 0 ;
  SIZE 2.09 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.35 0.525 1.46 0.7 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.75 0.525 1.84 0.7 ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235 1.065 0.745 1.135 ;
        RECT 0.235 0.33 0.745 0.4 ;
        RECT 0.235 0.33 0.32 1.135 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.09 1.485 ;
        RECT 1.745 0.86 1.815 1.485 ;
        RECT 1.21 1.205 1.28 1.485 ;
        RECT 0.83 1.205 0.9 1.485 ;
        RECT 0.45 1.205 0.52 1.485 ;
        RECT 0.075 1.205 0.145 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.09 0.085 ;
        RECT 1.74 -0.085 1.81 0.195 ;
        RECT 1.365 -0.085 1.435 0.195 ;
        RECT 0.83 -0.085 0.9 0.195 ;
        RECT 0.45 -0.085 0.52 0.195 ;
        RECT 0.075 -0.085 0.145 0.335 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.935 0.15 2.005 0.995 ;
      RECT 0.945 0.265 1.015 0.66 ;
      RECT 0.945 0.265 2.005 0.335 ;
      RECT 1.365 0.895 1.435 1.14 ;
      RECT 0.59 0.895 1.63 0.965 ;
      RECT 1.56 0.4 1.63 0.965 ;
      RECT 0.59 0.465 0.66 0.965 ;
      RECT 0.73 0.725 1.28 0.795 ;
      RECT 1.21 0.4 1.28 0.795 ;
      RECT 0.73 0.615 0.8 0.795 ;
  END
END TBUF_X4

MACRO TBUF_X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUF_X8 0 0 ;
  SIZE 3.42 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.72 0.39 2.79 0.66 ;
        RECT 2.14 0.39 2.79 0.46 ;
        RECT 1.95 0.56 2.21 0.63 ;
        RECT 2.14 0.39 2.21 0.63 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.465 0.725 3.08 0.795 ;
        RECT 3.01 0.525 3.08 0.795 ;
        RECT 2.465 0.525 2.6 0.795 ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.36 1.01 1.505 1.08 ;
        RECT 1.355 0.375 1.505 0.445 ;
        RECT 1.36 0.775 1.43 1.08 ;
        RECT 0.265 0.7 1.425 0.84 ;
        RECT 1.355 0.375 1.425 0.84 ;
        RECT 1.02 0.2 1.095 0.84 ;
        RECT 1.02 0.2 1.09 1.25 ;
        RECT 0.645 0.2 0.715 1.25 ;
        RECT 0.265 0.2 0.335 1.25 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 3.42 1.485 ;
        RECT 3.085 1.13 3.22 1.485 ;
        RECT 2.32 1.15 2.455 1.485 ;
        RECT 1.97 0.995 2.04 1.485 ;
        RECT 1.59 0.995 1.66 1.485 ;
        RECT 1.21 0.975 1.28 1.485 ;
        RECT 0.83 0.975 0.9 1.485 ;
        RECT 0.415 1.01 0.55 1.485 ;
        RECT 0.07 0.975 0.14 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 3.42 0.085 ;
        RECT 3.09 -0.085 3.225 0.16 ;
        RECT 2.7 -0.085 2.835 0.16 ;
        RECT 2.32 -0.085 2.455 0.16 ;
        RECT 1.56 -0.085 1.695 0.16 ;
        RECT 1.18 -0.085 1.315 0.16 ;
        RECT 0.8 -0.085 0.935 0.16 ;
        RECT 0.415 -0.085 0.55 0.375 ;
        RECT 0.07 -0.085 0.14 0.41 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 3.305 0.2 3.375 1.25 ;
      RECT 2.295 0.995 3.375 1.065 ;
      RECT 2.295 0.525 2.365 1.065 ;
      RECT 1.705 0.725 2.365 0.795 ;
      RECT 2.275 0.525 2.365 0.795 ;
      RECT 1.705 0.525 1.775 0.795 ;
      RECT 2.705 0.86 3.215 0.93 ;
      RECT 3.145 0.225 3.215 0.93 ;
      RECT 1.205 0.225 1.275 0.6 ;
      RECT 1.205 0.225 3.215 0.295 ;
      RECT 2.16 0.86 2.23 1.25 ;
      RECT 1.78 0.86 1.85 1.25 ;
      RECT 1.57 0.86 2.23 0.93 ;
      RECT 1.57 0.39 1.64 0.93 ;
      RECT 1.49 0.615 1.64 0.75 ;
      RECT 1.57 0.39 2.075 0.46 ;
  END
END TBUF_X8

MACRO TINV_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TINV_X1 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.45 0.65 0.585 0.72 ;
        RECT 0.175 0.84 0.52 0.98 ;
        RECT 0.45 0.65 0.52 0.98 ;
        RECT 0.175 0.625 0.245 0.98 ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.31 0.42 0.38 0.6 ;
        RECT 0.25 0.42 0.38 0.56 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.84 0.72 1.24 ;
        RECT 0.65 0.155 0.72 1.24 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 0.76 1.485 ;
        RECT 0.225 1.065 0.295 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 0.76 0.085 ;
        RECT 0.225 -0.085 0.295 0.195 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.04 0.195 0.11 1.24 ;
      RECT 0.45 0.495 0.585 0.565 ;
      RECT 0.45 0.275 0.52 0.565 ;
      RECT 0.04 0.275 0.52 0.345 ;
  END
END TINV_X1

MACRO TLAT_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLAT_X1 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.585 0.73 0.84 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.185 0.745 0.32 0.98 ;
    END
  END G
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.815 0.5 2.275 0.57 ;
        RECT 1.815 0.5 2.03 0.7 ;
    END
  END OE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.265 1.01 2.41 1.215 ;
        RECT 2.34 0.22 2.41 1.215 ;
        RECT 2.265 0.22 2.41 0.425 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 2.47 1.485 ;
        RECT 1.87 0.975 1.94 1.485 ;
        RECT 1.305 1.08 1.44 1.485 ;
        RECT 0.585 1.04 0.655 1.485 ;
        RECT 0.235 1.045 0.305 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 2.47 0.085 ;
        RECT 1.87 -0.085 1.94 0.32 ;
        RECT 1.335 -0.085 1.405 0.32 ;
        RECT 0.585 -0.085 0.655 0.46 ;
        RECT 0.235 -0.085 0.305 0.32 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.68 0.185 1.75 1.245 ;
      RECT 1.68 0.775 2.275 0.855 ;
      RECT 2.14 0.65 2.275 0.855 ;
      RECT 1.53 0.185 1.6 1.185 ;
      RECT 1.26 0.515 1.6 0.65 ;
      RECT 0.93 1.07 1.09 1.14 ;
      RECT 1.02 0.22 1.09 1.14 ;
      RECT 1.02 0.745 1.465 0.88 ;
      RECT 0.93 0.22 1.09 0.29 ;
      RECT 0.43 0.185 0.5 1.25 ;
      RECT 0.43 0.905 0.945 0.975 ;
      RECT 0.875 0.51 0.945 0.975 ;
      RECT 0.05 0.185 0.12 1.25 ;
      RECT 0.05 0.46 0.365 0.595 ;
  END
END TLAT_X1

MACRO XNOR2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2_X1 0 0 ;
  SIZE 1.14 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.65 0.555 0.81 0.625 ;
        RECT 0.65 0.39 0.72 0.625 ;
        RECT 0.185 0.39 0.72 0.46 ;
        RECT 0.185 0.39 0.32 0.56 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.35 0.84 0.965 0.91 ;
        RECT 0.895 0.525 0.965 0.91 ;
        RECT 0.35 0.84 0.51 0.98 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.98 1.1 1.05 ;
        RECT 1.03 0.295 1.1 1.05 ;
        RECT 0.785 0.295 1.1 0.365 ;
        RECT 0.63 0.98 0.7 1.25 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.14 1.485 ;
        RECT 1 1.115 1.07 1.485 ;
        RECT 0.43 1.115 0.5 1.485 ;
        RECT 0.05 1.115 0.12 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.14 0.085 ;
        RECT 0.395 -0.085 0.53 0.25 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.21 1.145 0.345 1.215 ;
      RECT 0.21 0.67 0.28 1.215 ;
      RECT 0.05 0.67 0.585 0.74 ;
      RECT 0.515 0.525 0.585 0.74 ;
      RECT 0.05 0.15 0.12 0.74 ;
      RECT 0.595 0.16 1.105 0.23 ;
  END
END XNOR2_X1

MACRO XNOR2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2_X2 0 0 ;
  SIZE 1.9 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.01 0.525 1.08 0.7 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.82 0.77 1.65 0.84 ;
        RECT 1.58 0.525 1.65 0.84 ;
        RECT 0.82 0.56 0.89 0.84 ;
        RECT 0.505 0.56 0.89 0.63 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.21 0.905 1.84 0.975 ;
        RECT 1.77 0.19 1.84 0.975 ;
        RECT 0.975 0.36 1.84 0.43 ;
        RECT 1.765 0.19 1.84 0.43 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.9 1.485 ;
        RECT 1.54 1.24 1.675 1.485 ;
        RECT 0.805 1.065 0.875 1.485 ;
        RECT 0.425 1.065 0.495 1.485 ;
        RECT 0.05 1.065 0.12 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.9 0.085 ;
        RECT 0.395 -0.085 0.53 0.16 ;
        RECT 0.05 -0.085 0.12 0.325 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.245 0.725 0.72 0.795 ;
      RECT 0.245 0.39 0.315 0.795 ;
      RECT 0.245 0.39 0.91 0.46 ;
      RECT 0.975 1.095 1.865 1.165 ;
      RECT 0.21 0.225 1.675 0.295 ;
  END
END XNOR2_X2

MACRO XOR2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2_X1 0 0 ;
  SIZE 1.14 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.63 0.525 0.755 0.66 ;
        RECT 0.175 0.73 0.7 0.8 ;
        RECT 0.63 0.525 0.7 0.8 ;
        RECT 0.175 0.665 0.245 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.82 0.525 0.945 0.66 ;
        RECT 0.305 0.875 0.89 0.945 ;
        RECT 0.82 0.525 0.89 0.945 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.775 1.04 1.08 1.11 ;
        RECT 1.01 0.35 1.08 1.11 ;
        RECT 0.62 0.35 1.08 0.42 ;
        RECT 0.62 0.15 0.69 0.42 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.14 1.485 ;
        RECT 0.42 1.15 0.49 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.14 0.085 ;
        RECT 0.99 -0.085 1.06 0.285 ;
        RECT 0.42 -0.085 0.49 0.285 ;
        RECT 0.04 -0.085 0.11 0.285 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.04 0.525 0.11 1.25 ;
      RECT 0.495 0.525 0.565 0.66 ;
      RECT 0.04 0.525 0.565 0.595 ;
      RECT 0.225 0.15 0.295 0.595 ;
      RECT 0.585 1.175 1.095 1.245 ;
  END
END XOR2_X1

MACRO XOR2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2_X2 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE FreePDK45_38x28_10R_NP_162NW_34O ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.255 0.395 1.325 0.66 ;
        RECT 0.745 0.395 1.325 0.465 ;
        RECT 0.745 0.285 0.82 0.66 ;
        RECT 0.06 0.285 0.82 0.355 ;
        RECT 0.06 0.285 0.165 0.7 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.365 0.77 1.125 0.84 ;
        RECT 0.99 0.56 1.125 0.84 ;
        RECT 0.365 0.56 0.5 0.84 ;
    END
  END B
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.8 0.905 1.465 0.975 ;
        RECT 1.39 0.26 1.465 0.975 ;
        RECT 0.885 0.26 1.465 0.33 ;
        RECT 0.885 0.15 0.955 0.33 ;
        RECT 0.61 0.15 0.955 0.22 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 1.315 1.71 1.485 ;
        RECT 1.585 1.205 1.655 1.485 ;
        RECT 0.445 1.205 0.515 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0 -0.085 1.71 0.085 ;
        RECT 1.585 -0.085 1.655 0.335 ;
        RECT 1.025 -0.085 1.095 0.195 ;
        RECT 0.445 -0.085 0.515 0.195 ;
        RECT 0.07 -0.085 0.14 0.21 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.04 1.04 1.6 1.11 ;
      RECT 1.53 0.525 1.6 1.11 ;
      RECT 0.23 0.425 0.3 1.11 ;
      RECT 0.575 0.425 0.645 0.66 ;
      RECT 0.23 0.425 0.645 0.495 ;
      RECT 0.61 1.175 1.5 1.245 ;
  END
END XOR2_X2

# END LIBRARY
#
# End of file
#
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_2048x39
  FOREIGN fakeram45_2048x39 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 206.910 BY 219.800 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.535 0.070 3.605 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.475 0.070 6.545 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.415 0.070 9.485 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.355 0.070 12.425 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.295 0.070 15.365 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.235 0.070 18.305 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.175 0.070 21.245 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.115 0.070 24.185 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.055 0.070 27.125 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.995 0.070 30.065 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.465 0.070 31.535 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.935 0.070 33.005 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.875 0.070 35.945 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.815 0.070 38.885 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.755 0.070 41.825 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.695 0.070 44.765 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.635 0.070 47.705 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.575 0.070 50.645 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.045 0.070 52.115 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.515 0.070 53.585 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.985 0.070 55.055 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.455 0.070 56.525 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END w_mask_in[38]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.595 0.070 63.665 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.065 0.070 65.135 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.535 0.070 66.605 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.475 0.070 69.545 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.945 0.070 71.015 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.415 0.070 72.485 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.355 0.070 75.425 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.825 0.070 76.895 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.295 0.070 78.365 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.235 0.070 81.305 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.705 0.070 82.775 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.175 0.070 84.245 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.115 0.070 87.185 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.585 0.070 88.655 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.055 0.070 90.125 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.525 0.070 91.595 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.995 0.070 93.065 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.465 0.070 94.535 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.935 0.070 96.005 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.405 0.070 97.475 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.875 0.070 98.945 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.345 0.070 100.415 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.815 0.070 101.885 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.285 0.070 103.355 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.755 0.070 104.825 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.225 0.070 106.295 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.695 0.070 107.765 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.165 0.070 109.235 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.635 0.070 110.705 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.105 0.070 112.175 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.575 0.070 113.645 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.045 0.070 115.115 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.515 0.070 116.585 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.985 0.070 118.055 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.455 0.070 119.525 ;
    END
  END rd_out[38]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.125 0.070 125.195 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.595 0.070 126.665 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.065 0.070 128.135 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.535 0.070 129.605 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.005 0.070 131.075 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.475 0.070 132.545 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.945 0.070 134.015 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.415 0.070 135.485 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.885 0.070 136.955 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.355 0.070 138.425 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.825 0.070 139.895 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.295 0.070 141.365 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.765 0.070 142.835 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.235 0.070 144.305 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.705 0.070 145.775 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.175 0.070 147.245 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.645 0.070 148.715 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.115 0.070 150.185 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.585 0.070 151.655 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.055 0.070 153.125 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.525 0.070 154.595 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.995 0.070 156.065 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.465 0.070 157.535 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.935 0.070 159.005 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.405 0.070 160.475 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.875 0.070 161.945 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.345 0.070 163.415 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.815 0.070 164.885 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.285 0.070 166.355 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.755 0.070 167.825 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.225 0.070 169.295 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.695 0.070 170.765 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.165 0.070 172.235 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.635 0.070 173.705 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.105 0.070 175.175 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.575 0.070 176.645 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.045 0.070 178.115 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.515 0.070 179.585 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.985 0.070 181.055 ;
    END
  END wd_in[38]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.655 0.070 186.725 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.125 0.070 188.195 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.595 0.070 189.665 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.065 0.070 191.135 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.535 0.070 192.605 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.005 0.070 194.075 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.475 0.070 195.545 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.945 0.070 197.015 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.415 0.070 198.485 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 199.885 0.070 199.955 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 201.355 0.070 201.425 ;
    END
  END addr_in[10]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 207.025 0.070 207.095 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 208.495 0.070 208.565 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 209.965 0.070 210.035 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 217.700 ;
      RECT 5.320 2.100 5.600 217.700 ;
      RECT 8.680 2.100 8.960 217.700 ;
      RECT 12.040 2.100 12.320 217.700 ;
      RECT 15.400 2.100 15.680 217.700 ;
      RECT 18.760 2.100 19.040 217.700 ;
      RECT 22.120 2.100 22.400 217.700 ;
      RECT 25.480 2.100 25.760 217.700 ;
      RECT 28.840 2.100 29.120 217.700 ;
      RECT 32.200 2.100 32.480 217.700 ;
      RECT 35.560 2.100 35.840 217.700 ;
      RECT 38.920 2.100 39.200 217.700 ;
      RECT 42.280 2.100 42.560 217.700 ;
      RECT 45.640 2.100 45.920 217.700 ;
      RECT 49.000 2.100 49.280 217.700 ;
      RECT 52.360 2.100 52.640 217.700 ;
      RECT 55.720 2.100 56.000 217.700 ;
      RECT 59.080 2.100 59.360 217.700 ;
      RECT 62.440 2.100 62.720 217.700 ;
      RECT 65.800 2.100 66.080 217.700 ;
      RECT 69.160 2.100 69.440 217.700 ;
      RECT 72.520 2.100 72.800 217.700 ;
      RECT 75.880 2.100 76.160 217.700 ;
      RECT 79.240 2.100 79.520 217.700 ;
      RECT 82.600 2.100 82.880 217.700 ;
      RECT 85.960 2.100 86.240 217.700 ;
      RECT 89.320 2.100 89.600 217.700 ;
      RECT 92.680 2.100 92.960 217.700 ;
      RECT 96.040 2.100 96.320 217.700 ;
      RECT 99.400 2.100 99.680 217.700 ;
      RECT 102.760 2.100 103.040 217.700 ;
      RECT 106.120 2.100 106.400 217.700 ;
      RECT 109.480 2.100 109.760 217.700 ;
      RECT 112.840 2.100 113.120 217.700 ;
      RECT 116.200 2.100 116.480 217.700 ;
      RECT 119.560 2.100 119.840 217.700 ;
      RECT 122.920 2.100 123.200 217.700 ;
      RECT 126.280 2.100 126.560 217.700 ;
      RECT 129.640 2.100 129.920 217.700 ;
      RECT 133.000 2.100 133.280 217.700 ;
      RECT 136.360 2.100 136.640 217.700 ;
      RECT 139.720 2.100 140.000 217.700 ;
      RECT 143.080 2.100 143.360 217.700 ;
      RECT 146.440 2.100 146.720 217.700 ;
      RECT 149.800 2.100 150.080 217.700 ;
      RECT 153.160 2.100 153.440 217.700 ;
      RECT 156.520 2.100 156.800 217.700 ;
      RECT 159.880 2.100 160.160 217.700 ;
      RECT 163.240 2.100 163.520 217.700 ;
      RECT 166.600 2.100 166.880 217.700 ;
      RECT 169.960 2.100 170.240 217.700 ;
      RECT 173.320 2.100 173.600 217.700 ;
      RECT 176.680 2.100 176.960 217.700 ;
      RECT 180.040 2.100 180.320 217.700 ;
      RECT 183.400 2.100 183.680 217.700 ;
      RECT 186.760 2.100 187.040 217.700 ;
      RECT 190.120 2.100 190.400 217.700 ;
      RECT 193.480 2.100 193.760 217.700 ;
      RECT 196.840 2.100 197.120 217.700 ;
      RECT 200.200 2.100 200.480 217.700 ;
      RECT 203.560 2.100 203.840 217.700 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 217.700 ;
      RECT 7.000 2.100 7.280 217.700 ;
      RECT 10.360 2.100 10.640 217.700 ;
      RECT 13.720 2.100 14.000 217.700 ;
      RECT 17.080 2.100 17.360 217.700 ;
      RECT 20.440 2.100 20.720 217.700 ;
      RECT 23.800 2.100 24.080 217.700 ;
      RECT 27.160 2.100 27.440 217.700 ;
      RECT 30.520 2.100 30.800 217.700 ;
      RECT 33.880 2.100 34.160 217.700 ;
      RECT 37.240 2.100 37.520 217.700 ;
      RECT 40.600 2.100 40.880 217.700 ;
      RECT 43.960 2.100 44.240 217.700 ;
      RECT 47.320 2.100 47.600 217.700 ;
      RECT 50.680 2.100 50.960 217.700 ;
      RECT 54.040 2.100 54.320 217.700 ;
      RECT 57.400 2.100 57.680 217.700 ;
      RECT 60.760 2.100 61.040 217.700 ;
      RECT 64.120 2.100 64.400 217.700 ;
      RECT 67.480 2.100 67.760 217.700 ;
      RECT 70.840 2.100 71.120 217.700 ;
      RECT 74.200 2.100 74.480 217.700 ;
      RECT 77.560 2.100 77.840 217.700 ;
      RECT 80.920 2.100 81.200 217.700 ;
      RECT 84.280 2.100 84.560 217.700 ;
      RECT 87.640 2.100 87.920 217.700 ;
      RECT 91.000 2.100 91.280 217.700 ;
      RECT 94.360 2.100 94.640 217.700 ;
      RECT 97.720 2.100 98.000 217.700 ;
      RECT 101.080 2.100 101.360 217.700 ;
      RECT 104.440 2.100 104.720 217.700 ;
      RECT 107.800 2.100 108.080 217.700 ;
      RECT 111.160 2.100 111.440 217.700 ;
      RECT 114.520 2.100 114.800 217.700 ;
      RECT 117.880 2.100 118.160 217.700 ;
      RECT 121.240 2.100 121.520 217.700 ;
      RECT 124.600 2.100 124.880 217.700 ;
      RECT 127.960 2.100 128.240 217.700 ;
      RECT 131.320 2.100 131.600 217.700 ;
      RECT 134.680 2.100 134.960 217.700 ;
      RECT 138.040 2.100 138.320 217.700 ;
      RECT 141.400 2.100 141.680 217.700 ;
      RECT 144.760 2.100 145.040 217.700 ;
      RECT 148.120 2.100 148.400 217.700 ;
      RECT 151.480 2.100 151.760 217.700 ;
      RECT 154.840 2.100 155.120 217.700 ;
      RECT 158.200 2.100 158.480 217.700 ;
      RECT 161.560 2.100 161.840 217.700 ;
      RECT 164.920 2.100 165.200 217.700 ;
      RECT 168.280 2.100 168.560 217.700 ;
      RECT 171.640 2.100 171.920 217.700 ;
      RECT 175.000 2.100 175.280 217.700 ;
      RECT 178.360 2.100 178.640 217.700 ;
      RECT 181.720 2.100 182.000 217.700 ;
      RECT 185.080 2.100 185.360 217.700 ;
      RECT 188.440 2.100 188.720 217.700 ;
      RECT 191.800 2.100 192.080 217.700 ;
      RECT 195.160 2.100 195.440 217.700 ;
      RECT 198.520 2.100 198.800 217.700 ;
      RECT 201.880 2.100 202.160 217.700 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 206.910 219.800 ;
    LAYER metal2 ;
    RECT 0 0 206.910 219.800 ;
    LAYER metal3 ;
    RECT 0.070 0 206.910 219.800 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 3.535 ;
    RECT 0 3.605 0.070 5.005 ;
    RECT 0 5.075 0.070 6.475 ;
    RECT 0 6.545 0.070 7.945 ;
    RECT 0 8.015 0.070 9.415 ;
    RECT 0 9.485 0.070 10.885 ;
    RECT 0 10.955 0.070 12.355 ;
    RECT 0 12.425 0.070 13.825 ;
    RECT 0 13.895 0.070 15.295 ;
    RECT 0 15.365 0.070 16.765 ;
    RECT 0 16.835 0.070 18.235 ;
    RECT 0 18.305 0.070 19.705 ;
    RECT 0 19.775 0.070 21.175 ;
    RECT 0 21.245 0.070 22.645 ;
    RECT 0 22.715 0.070 24.115 ;
    RECT 0 24.185 0.070 25.585 ;
    RECT 0 25.655 0.070 27.055 ;
    RECT 0 27.125 0.070 28.525 ;
    RECT 0 28.595 0.070 29.995 ;
    RECT 0 30.065 0.070 31.465 ;
    RECT 0 31.535 0.070 32.935 ;
    RECT 0 33.005 0.070 34.405 ;
    RECT 0 34.475 0.070 35.875 ;
    RECT 0 35.945 0.070 37.345 ;
    RECT 0 37.415 0.070 38.815 ;
    RECT 0 38.885 0.070 40.285 ;
    RECT 0 40.355 0.070 41.755 ;
    RECT 0 41.825 0.070 43.225 ;
    RECT 0 43.295 0.070 44.695 ;
    RECT 0 44.765 0.070 46.165 ;
    RECT 0 46.235 0.070 47.635 ;
    RECT 0 47.705 0.070 49.105 ;
    RECT 0 49.175 0.070 50.575 ;
    RECT 0 50.645 0.070 52.045 ;
    RECT 0 52.115 0.070 53.515 ;
    RECT 0 53.585 0.070 54.985 ;
    RECT 0 55.055 0.070 56.455 ;
    RECT 0 56.525 0.070 57.925 ;
    RECT 0 57.995 0.070 63.595 ;
    RECT 0 63.665 0.070 65.065 ;
    RECT 0 65.135 0.070 66.535 ;
    RECT 0 66.605 0.070 68.005 ;
    RECT 0 68.075 0.070 69.475 ;
    RECT 0 69.545 0.070 70.945 ;
    RECT 0 71.015 0.070 72.415 ;
    RECT 0 72.485 0.070 73.885 ;
    RECT 0 73.955 0.070 75.355 ;
    RECT 0 75.425 0.070 76.825 ;
    RECT 0 76.895 0.070 78.295 ;
    RECT 0 78.365 0.070 79.765 ;
    RECT 0 79.835 0.070 81.235 ;
    RECT 0 81.305 0.070 82.705 ;
    RECT 0 82.775 0.070 84.175 ;
    RECT 0 84.245 0.070 85.645 ;
    RECT 0 85.715 0.070 87.115 ;
    RECT 0 87.185 0.070 88.585 ;
    RECT 0 88.655 0.070 90.055 ;
    RECT 0 90.125 0.070 91.525 ;
    RECT 0 91.595 0.070 92.995 ;
    RECT 0 93.065 0.070 94.465 ;
    RECT 0 94.535 0.070 95.935 ;
    RECT 0 96.005 0.070 97.405 ;
    RECT 0 97.475 0.070 98.875 ;
    RECT 0 98.945 0.070 100.345 ;
    RECT 0 100.415 0.070 101.815 ;
    RECT 0 101.885 0.070 103.285 ;
    RECT 0 103.355 0.070 104.755 ;
    RECT 0 104.825 0.070 106.225 ;
    RECT 0 106.295 0.070 107.695 ;
    RECT 0 107.765 0.070 109.165 ;
    RECT 0 109.235 0.070 110.635 ;
    RECT 0 110.705 0.070 112.105 ;
    RECT 0 112.175 0.070 113.575 ;
    RECT 0 113.645 0.070 115.045 ;
    RECT 0 115.115 0.070 116.515 ;
    RECT 0 116.585 0.070 117.985 ;
    RECT 0 118.055 0.070 119.455 ;
    RECT 0 119.525 0.070 125.125 ;
    RECT 0 125.195 0.070 126.595 ;
    RECT 0 126.665 0.070 128.065 ;
    RECT 0 128.135 0.070 129.535 ;
    RECT 0 129.605 0.070 131.005 ;
    RECT 0 131.075 0.070 132.475 ;
    RECT 0 132.545 0.070 133.945 ;
    RECT 0 134.015 0.070 135.415 ;
    RECT 0 135.485 0.070 136.885 ;
    RECT 0 136.955 0.070 138.355 ;
    RECT 0 138.425 0.070 139.825 ;
    RECT 0 139.895 0.070 141.295 ;
    RECT 0 141.365 0.070 142.765 ;
    RECT 0 142.835 0.070 144.235 ;
    RECT 0 144.305 0.070 145.705 ;
    RECT 0 145.775 0.070 147.175 ;
    RECT 0 147.245 0.070 148.645 ;
    RECT 0 148.715 0.070 150.115 ;
    RECT 0 150.185 0.070 151.585 ;
    RECT 0 151.655 0.070 153.055 ;
    RECT 0 153.125 0.070 154.525 ;
    RECT 0 154.595 0.070 155.995 ;
    RECT 0 156.065 0.070 157.465 ;
    RECT 0 157.535 0.070 158.935 ;
    RECT 0 159.005 0.070 160.405 ;
    RECT 0 160.475 0.070 161.875 ;
    RECT 0 161.945 0.070 163.345 ;
    RECT 0 163.415 0.070 164.815 ;
    RECT 0 164.885 0.070 166.285 ;
    RECT 0 166.355 0.070 167.755 ;
    RECT 0 167.825 0.070 169.225 ;
    RECT 0 169.295 0.070 170.695 ;
    RECT 0 170.765 0.070 172.165 ;
    RECT 0 172.235 0.070 173.635 ;
    RECT 0 173.705 0.070 175.105 ;
    RECT 0 175.175 0.070 176.575 ;
    RECT 0 176.645 0.070 178.045 ;
    RECT 0 178.115 0.070 179.515 ;
    RECT 0 179.585 0.070 180.985 ;
    RECT 0 181.055 0.070 186.655 ;
    RECT 0 186.725 0.070 188.125 ;
    RECT 0 188.195 0.070 189.595 ;
    RECT 0 189.665 0.070 191.065 ;
    RECT 0 191.135 0.070 192.535 ;
    RECT 0 192.605 0.070 194.005 ;
    RECT 0 194.075 0.070 195.475 ;
    RECT 0 195.545 0.070 196.945 ;
    RECT 0 197.015 0.070 198.415 ;
    RECT 0 198.485 0.070 199.885 ;
    RECT 0 199.955 0.070 201.355 ;
    RECT 0 201.425 0.070 207.025 ;
    RECT 0 207.095 0.070 208.495 ;
    RECT 0 208.565 0.070 209.965 ;
    RECT 0 210.035 0.070 219.800 ;
    LAYER metal4 ;
    RECT 0 0 206.910 2.100 ;
    RECT 0 217.700 206.910 219.800 ;
    RECT 0.000 2.100 1.960 217.700 ;
    RECT 2.240 2.100 3.640 217.700 ;
    RECT 3.920 2.100 5.320 217.700 ;
    RECT 5.600 2.100 7.000 217.700 ;
    RECT 7.280 2.100 8.680 217.700 ;
    RECT 8.960 2.100 10.360 217.700 ;
    RECT 10.640 2.100 12.040 217.700 ;
    RECT 12.320 2.100 13.720 217.700 ;
    RECT 14.000 2.100 15.400 217.700 ;
    RECT 15.680 2.100 17.080 217.700 ;
    RECT 17.360 2.100 18.760 217.700 ;
    RECT 19.040 2.100 20.440 217.700 ;
    RECT 20.720 2.100 22.120 217.700 ;
    RECT 22.400 2.100 23.800 217.700 ;
    RECT 24.080 2.100 25.480 217.700 ;
    RECT 25.760 2.100 27.160 217.700 ;
    RECT 27.440 2.100 28.840 217.700 ;
    RECT 29.120 2.100 30.520 217.700 ;
    RECT 30.800 2.100 32.200 217.700 ;
    RECT 32.480 2.100 33.880 217.700 ;
    RECT 34.160 2.100 35.560 217.700 ;
    RECT 35.840 2.100 37.240 217.700 ;
    RECT 37.520 2.100 38.920 217.700 ;
    RECT 39.200 2.100 40.600 217.700 ;
    RECT 40.880 2.100 42.280 217.700 ;
    RECT 42.560 2.100 43.960 217.700 ;
    RECT 44.240 2.100 45.640 217.700 ;
    RECT 45.920 2.100 47.320 217.700 ;
    RECT 47.600 2.100 49.000 217.700 ;
    RECT 49.280 2.100 50.680 217.700 ;
    RECT 50.960 2.100 52.360 217.700 ;
    RECT 52.640 2.100 54.040 217.700 ;
    RECT 54.320 2.100 55.720 217.700 ;
    RECT 56.000 2.100 57.400 217.700 ;
    RECT 57.680 2.100 59.080 217.700 ;
    RECT 59.360 2.100 60.760 217.700 ;
    RECT 61.040 2.100 62.440 217.700 ;
    RECT 62.720 2.100 64.120 217.700 ;
    RECT 64.400 2.100 65.800 217.700 ;
    RECT 66.080 2.100 67.480 217.700 ;
    RECT 67.760 2.100 69.160 217.700 ;
    RECT 69.440 2.100 70.840 217.700 ;
    RECT 71.120 2.100 72.520 217.700 ;
    RECT 72.800 2.100 74.200 217.700 ;
    RECT 74.480 2.100 75.880 217.700 ;
    RECT 76.160 2.100 77.560 217.700 ;
    RECT 77.840 2.100 79.240 217.700 ;
    RECT 79.520 2.100 80.920 217.700 ;
    RECT 81.200 2.100 82.600 217.700 ;
    RECT 82.880 2.100 84.280 217.700 ;
    RECT 84.560 2.100 85.960 217.700 ;
    RECT 86.240 2.100 87.640 217.700 ;
    RECT 87.920 2.100 89.320 217.700 ;
    RECT 89.600 2.100 91.000 217.700 ;
    RECT 91.280 2.100 92.680 217.700 ;
    RECT 92.960 2.100 94.360 217.700 ;
    RECT 94.640 2.100 96.040 217.700 ;
    RECT 96.320 2.100 97.720 217.700 ;
    RECT 98.000 2.100 99.400 217.700 ;
    RECT 99.680 2.100 101.080 217.700 ;
    RECT 101.360 2.100 102.760 217.700 ;
    RECT 103.040 2.100 104.440 217.700 ;
    RECT 104.720 2.100 106.120 217.700 ;
    RECT 106.400 2.100 107.800 217.700 ;
    RECT 108.080 2.100 109.480 217.700 ;
    RECT 109.760 2.100 111.160 217.700 ;
    RECT 111.440 2.100 112.840 217.700 ;
    RECT 113.120 2.100 114.520 217.700 ;
    RECT 114.800 2.100 116.200 217.700 ;
    RECT 116.480 2.100 117.880 217.700 ;
    RECT 118.160 2.100 119.560 217.700 ;
    RECT 119.840 2.100 121.240 217.700 ;
    RECT 121.520 2.100 122.920 217.700 ;
    RECT 123.200 2.100 124.600 217.700 ;
    RECT 124.880 2.100 126.280 217.700 ;
    RECT 126.560 2.100 127.960 217.700 ;
    RECT 128.240 2.100 129.640 217.700 ;
    RECT 129.920 2.100 131.320 217.700 ;
    RECT 131.600 2.100 133.000 217.700 ;
    RECT 133.280 2.100 134.680 217.700 ;
    RECT 134.960 2.100 136.360 217.700 ;
    RECT 136.640 2.100 138.040 217.700 ;
    RECT 138.320 2.100 139.720 217.700 ;
    RECT 140.000 2.100 141.400 217.700 ;
    RECT 141.680 2.100 143.080 217.700 ;
    RECT 143.360 2.100 144.760 217.700 ;
    RECT 145.040 2.100 146.440 217.700 ;
    RECT 146.720 2.100 148.120 217.700 ;
    RECT 148.400 2.100 149.800 217.700 ;
    RECT 150.080 2.100 151.480 217.700 ;
    RECT 151.760 2.100 153.160 217.700 ;
    RECT 153.440 2.100 154.840 217.700 ;
    RECT 155.120 2.100 156.520 217.700 ;
    RECT 156.800 2.100 158.200 217.700 ;
    RECT 158.480 2.100 159.880 217.700 ;
    RECT 160.160 2.100 161.560 217.700 ;
    RECT 161.840 2.100 163.240 217.700 ;
    RECT 163.520 2.100 164.920 217.700 ;
    RECT 165.200 2.100 166.600 217.700 ;
    RECT 166.880 2.100 168.280 217.700 ;
    RECT 168.560 2.100 169.960 217.700 ;
    RECT 170.240 2.100 171.640 217.700 ;
    RECT 171.920 2.100 173.320 217.700 ;
    RECT 173.600 2.100 175.000 217.700 ;
    RECT 175.280 2.100 176.680 217.700 ;
    RECT 176.960 2.100 178.360 217.700 ;
    RECT 178.640 2.100 180.040 217.700 ;
    RECT 180.320 2.100 181.720 217.700 ;
    RECT 182.000 2.100 183.400 217.700 ;
    RECT 183.680 2.100 185.080 217.700 ;
    RECT 185.360 2.100 186.760 217.700 ;
    RECT 187.040 2.100 188.440 217.700 ;
    RECT 188.720 2.100 190.120 217.700 ;
    RECT 190.400 2.100 191.800 217.700 ;
    RECT 192.080 2.100 193.480 217.700 ;
    RECT 193.760 2.100 195.160 217.700 ;
    RECT 195.440 2.100 196.840 217.700 ;
    RECT 197.120 2.100 198.520 217.700 ;
    RECT 198.800 2.100 200.200 217.700 ;
    RECT 200.480 2.100 201.880 217.700 ;
    RECT 202.160 2.100 203.560 217.700 ;
    RECT 203.840 2.100 206.910 217.700 ;
    LAYER OVERLAP ;
    RECT 0 0 206.910 219.800 ;
  END
END fakeram45_2048x39

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_1024x32
  FOREIGN fakeram45_1024x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 152.190 BY 107.800 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.785 0.070 8.855 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.985 0.070 13.055 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.505 0.070 15.575 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.345 0.070 16.415 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.185 0.070 17.255 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.025 0.070 18.095 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.545 0.070 20.615 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.225 0.070 22.295 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.905 0.070 23.975 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.425 0.070 26.495 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.105 0.070 28.175 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.045 0.070 31.115 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.885 0.070 31.955 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.325 0.070 45.395 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.205 0.070 51.275 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.045 0.070 52.115 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.085 0.070 57.155 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.025 0.070 60.095 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.865 0.070 60.935 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.705 0.070 61.775 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.545 0.070 62.615 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.385 0.070 63.455 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.225 0.070 64.295 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.065 0.070 65.135 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.905 0.070 65.975 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.745 0.070 66.815 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.585 0.070 67.655 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.425 0.070 68.495 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.265 0.070 69.335 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.105 0.070 70.175 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.945 0.070 71.015 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.785 0.070 71.855 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.625 0.070 72.695 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.465 0.070 73.535 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.305 0.070 74.375 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.145 0.070 75.215 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.825 0.070 76.895 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.665 0.070 77.735 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.505 0.070 78.575 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.345 0.070 79.415 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.185 0.070 80.255 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.025 0.070 81.095 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.705 0.070 82.775 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.545 0.070 83.615 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.385 0.070 84.455 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.225 0.070 85.295 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.065 0.070 86.135 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.005 0.070 89.075 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.845 0.070 89.915 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.685 0.070 90.755 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.525 0.070 91.595 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.365 0.070 92.435 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.205 0.070 93.275 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.045 0.070 94.115 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.885 0.070 94.955 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.725 0.070 95.795 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.565 0.070 96.635 ;
    END
  END addr_in[9]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.505 0.070 99.575 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.345 0.070 100.415 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.185 0.070 101.255 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 105.700 ;
      RECT 5.320 2.100 5.600 105.700 ;
      RECT 8.680 2.100 8.960 105.700 ;
      RECT 12.040 2.100 12.320 105.700 ;
      RECT 15.400 2.100 15.680 105.700 ;
      RECT 18.760 2.100 19.040 105.700 ;
      RECT 22.120 2.100 22.400 105.700 ;
      RECT 25.480 2.100 25.760 105.700 ;
      RECT 28.840 2.100 29.120 105.700 ;
      RECT 32.200 2.100 32.480 105.700 ;
      RECT 35.560 2.100 35.840 105.700 ;
      RECT 38.920 2.100 39.200 105.700 ;
      RECT 42.280 2.100 42.560 105.700 ;
      RECT 45.640 2.100 45.920 105.700 ;
      RECT 49.000 2.100 49.280 105.700 ;
      RECT 52.360 2.100 52.640 105.700 ;
      RECT 55.720 2.100 56.000 105.700 ;
      RECT 59.080 2.100 59.360 105.700 ;
      RECT 62.440 2.100 62.720 105.700 ;
      RECT 65.800 2.100 66.080 105.700 ;
      RECT 69.160 2.100 69.440 105.700 ;
      RECT 72.520 2.100 72.800 105.700 ;
      RECT 75.880 2.100 76.160 105.700 ;
      RECT 79.240 2.100 79.520 105.700 ;
      RECT 82.600 2.100 82.880 105.700 ;
      RECT 85.960 2.100 86.240 105.700 ;
      RECT 89.320 2.100 89.600 105.700 ;
      RECT 92.680 2.100 92.960 105.700 ;
      RECT 96.040 2.100 96.320 105.700 ;
      RECT 99.400 2.100 99.680 105.700 ;
      RECT 102.760 2.100 103.040 105.700 ;
      RECT 106.120 2.100 106.400 105.700 ;
      RECT 109.480 2.100 109.760 105.700 ;
      RECT 112.840 2.100 113.120 105.700 ;
      RECT 116.200 2.100 116.480 105.700 ;
      RECT 119.560 2.100 119.840 105.700 ;
      RECT 122.920 2.100 123.200 105.700 ;
      RECT 126.280 2.100 126.560 105.700 ;
      RECT 129.640 2.100 129.920 105.700 ;
      RECT 133.000 2.100 133.280 105.700 ;
      RECT 136.360 2.100 136.640 105.700 ;
      RECT 139.720 2.100 140.000 105.700 ;
      RECT 143.080 2.100 143.360 105.700 ;
      RECT 146.440 2.100 146.720 105.700 ;
      RECT 149.800 2.100 150.080 105.700 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 105.700 ;
      RECT 7.000 2.100 7.280 105.700 ;
      RECT 10.360 2.100 10.640 105.700 ;
      RECT 13.720 2.100 14.000 105.700 ;
      RECT 17.080 2.100 17.360 105.700 ;
      RECT 20.440 2.100 20.720 105.700 ;
      RECT 23.800 2.100 24.080 105.700 ;
      RECT 27.160 2.100 27.440 105.700 ;
      RECT 30.520 2.100 30.800 105.700 ;
      RECT 33.880 2.100 34.160 105.700 ;
      RECT 37.240 2.100 37.520 105.700 ;
      RECT 40.600 2.100 40.880 105.700 ;
      RECT 43.960 2.100 44.240 105.700 ;
      RECT 47.320 2.100 47.600 105.700 ;
      RECT 50.680 2.100 50.960 105.700 ;
      RECT 54.040 2.100 54.320 105.700 ;
      RECT 57.400 2.100 57.680 105.700 ;
      RECT 60.760 2.100 61.040 105.700 ;
      RECT 64.120 2.100 64.400 105.700 ;
      RECT 67.480 2.100 67.760 105.700 ;
      RECT 70.840 2.100 71.120 105.700 ;
      RECT 74.200 2.100 74.480 105.700 ;
      RECT 77.560 2.100 77.840 105.700 ;
      RECT 80.920 2.100 81.200 105.700 ;
      RECT 84.280 2.100 84.560 105.700 ;
      RECT 87.640 2.100 87.920 105.700 ;
      RECT 91.000 2.100 91.280 105.700 ;
      RECT 94.360 2.100 94.640 105.700 ;
      RECT 97.720 2.100 98.000 105.700 ;
      RECT 101.080 2.100 101.360 105.700 ;
      RECT 104.440 2.100 104.720 105.700 ;
      RECT 107.800 2.100 108.080 105.700 ;
      RECT 111.160 2.100 111.440 105.700 ;
      RECT 114.520 2.100 114.800 105.700 ;
      RECT 117.880 2.100 118.160 105.700 ;
      RECT 121.240 2.100 121.520 105.700 ;
      RECT 124.600 2.100 124.880 105.700 ;
      RECT 127.960 2.100 128.240 105.700 ;
      RECT 131.320 2.100 131.600 105.700 ;
      RECT 134.680 2.100 134.960 105.700 ;
      RECT 138.040 2.100 138.320 105.700 ;
      RECT 141.400 2.100 141.680 105.700 ;
      RECT 144.760 2.100 145.040 105.700 ;
      RECT 148.120 2.100 148.400 105.700 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 152.190 107.800 ;
    LAYER metal2 ;
    RECT 0 0 152.190 107.800 ;
    LAYER metal3 ;
    RECT 0.070 0 152.190 107.800 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.905 ;
    RECT 0 2.975 0.070 3.745 ;
    RECT 0 3.815 0.070 4.585 ;
    RECT 0 4.655 0.070 5.425 ;
    RECT 0 5.495 0.070 6.265 ;
    RECT 0 6.335 0.070 7.105 ;
    RECT 0 7.175 0.070 7.945 ;
    RECT 0 8.015 0.070 8.785 ;
    RECT 0 8.855 0.070 9.625 ;
    RECT 0 9.695 0.070 10.465 ;
    RECT 0 10.535 0.070 11.305 ;
    RECT 0 11.375 0.070 12.145 ;
    RECT 0 12.215 0.070 12.985 ;
    RECT 0 13.055 0.070 13.825 ;
    RECT 0 13.895 0.070 14.665 ;
    RECT 0 14.735 0.070 15.505 ;
    RECT 0 15.575 0.070 16.345 ;
    RECT 0 16.415 0.070 17.185 ;
    RECT 0 17.255 0.070 18.025 ;
    RECT 0 18.095 0.070 18.865 ;
    RECT 0 18.935 0.070 19.705 ;
    RECT 0 19.775 0.070 20.545 ;
    RECT 0 20.615 0.070 21.385 ;
    RECT 0 21.455 0.070 22.225 ;
    RECT 0 22.295 0.070 23.065 ;
    RECT 0 23.135 0.070 23.905 ;
    RECT 0 23.975 0.070 24.745 ;
    RECT 0 24.815 0.070 25.585 ;
    RECT 0 25.655 0.070 26.425 ;
    RECT 0 26.495 0.070 27.265 ;
    RECT 0 27.335 0.070 28.105 ;
    RECT 0 28.175 0.070 31.045 ;
    RECT 0 31.115 0.070 31.885 ;
    RECT 0 31.955 0.070 32.725 ;
    RECT 0 32.795 0.070 33.565 ;
    RECT 0 33.635 0.070 34.405 ;
    RECT 0 34.475 0.070 35.245 ;
    RECT 0 35.315 0.070 36.085 ;
    RECT 0 36.155 0.070 36.925 ;
    RECT 0 36.995 0.070 37.765 ;
    RECT 0 37.835 0.070 38.605 ;
    RECT 0 38.675 0.070 39.445 ;
    RECT 0 39.515 0.070 40.285 ;
    RECT 0 40.355 0.070 41.125 ;
    RECT 0 41.195 0.070 41.965 ;
    RECT 0 42.035 0.070 42.805 ;
    RECT 0 42.875 0.070 43.645 ;
    RECT 0 43.715 0.070 44.485 ;
    RECT 0 44.555 0.070 45.325 ;
    RECT 0 45.395 0.070 46.165 ;
    RECT 0 46.235 0.070 47.005 ;
    RECT 0 47.075 0.070 47.845 ;
    RECT 0 47.915 0.070 48.685 ;
    RECT 0 48.755 0.070 49.525 ;
    RECT 0 49.595 0.070 50.365 ;
    RECT 0 50.435 0.070 51.205 ;
    RECT 0 51.275 0.070 52.045 ;
    RECT 0 52.115 0.070 52.885 ;
    RECT 0 52.955 0.070 53.725 ;
    RECT 0 53.795 0.070 54.565 ;
    RECT 0 54.635 0.070 55.405 ;
    RECT 0 55.475 0.070 56.245 ;
    RECT 0 56.315 0.070 57.085 ;
    RECT 0 57.155 0.070 60.025 ;
    RECT 0 60.095 0.070 60.865 ;
    RECT 0 60.935 0.070 61.705 ;
    RECT 0 61.775 0.070 62.545 ;
    RECT 0 62.615 0.070 63.385 ;
    RECT 0 63.455 0.070 64.225 ;
    RECT 0 64.295 0.070 65.065 ;
    RECT 0 65.135 0.070 65.905 ;
    RECT 0 65.975 0.070 66.745 ;
    RECT 0 66.815 0.070 67.585 ;
    RECT 0 67.655 0.070 68.425 ;
    RECT 0 68.495 0.070 69.265 ;
    RECT 0 69.335 0.070 70.105 ;
    RECT 0 70.175 0.070 70.945 ;
    RECT 0 71.015 0.070 71.785 ;
    RECT 0 71.855 0.070 72.625 ;
    RECT 0 72.695 0.070 73.465 ;
    RECT 0 73.535 0.070 74.305 ;
    RECT 0 74.375 0.070 75.145 ;
    RECT 0 75.215 0.070 75.985 ;
    RECT 0 76.055 0.070 76.825 ;
    RECT 0 76.895 0.070 77.665 ;
    RECT 0 77.735 0.070 78.505 ;
    RECT 0 78.575 0.070 79.345 ;
    RECT 0 79.415 0.070 80.185 ;
    RECT 0 80.255 0.070 81.025 ;
    RECT 0 81.095 0.070 81.865 ;
    RECT 0 81.935 0.070 82.705 ;
    RECT 0 82.775 0.070 83.545 ;
    RECT 0 83.615 0.070 84.385 ;
    RECT 0 84.455 0.070 85.225 ;
    RECT 0 85.295 0.070 86.065 ;
    RECT 0 86.135 0.070 89.005 ;
    RECT 0 89.075 0.070 89.845 ;
    RECT 0 89.915 0.070 90.685 ;
    RECT 0 90.755 0.070 91.525 ;
    RECT 0 91.595 0.070 92.365 ;
    RECT 0 92.435 0.070 93.205 ;
    RECT 0 93.275 0.070 94.045 ;
    RECT 0 94.115 0.070 94.885 ;
    RECT 0 94.955 0.070 95.725 ;
    RECT 0 95.795 0.070 96.565 ;
    RECT 0 96.635 0.070 99.505 ;
    RECT 0 99.575 0.070 100.345 ;
    RECT 0 100.415 0.070 101.185 ;
    RECT 0 101.255 0.070 107.800 ;
    LAYER metal4 ;
    RECT 0 0 152.190 2.100 ;
    RECT 0 105.700 152.190 107.800 ;
    RECT 0.000 2.100 1.960 105.700 ;
    RECT 2.240 2.100 3.640 105.700 ;
    RECT 3.920 2.100 5.320 105.700 ;
    RECT 5.600 2.100 7.000 105.700 ;
    RECT 7.280 2.100 8.680 105.700 ;
    RECT 8.960 2.100 10.360 105.700 ;
    RECT 10.640 2.100 12.040 105.700 ;
    RECT 12.320 2.100 13.720 105.700 ;
    RECT 14.000 2.100 15.400 105.700 ;
    RECT 15.680 2.100 17.080 105.700 ;
    RECT 17.360 2.100 18.760 105.700 ;
    RECT 19.040 2.100 20.440 105.700 ;
    RECT 20.720 2.100 22.120 105.700 ;
    RECT 22.400 2.100 23.800 105.700 ;
    RECT 24.080 2.100 25.480 105.700 ;
    RECT 25.760 2.100 27.160 105.700 ;
    RECT 27.440 2.100 28.840 105.700 ;
    RECT 29.120 2.100 30.520 105.700 ;
    RECT 30.800 2.100 32.200 105.700 ;
    RECT 32.480 2.100 33.880 105.700 ;
    RECT 34.160 2.100 35.560 105.700 ;
    RECT 35.840 2.100 37.240 105.700 ;
    RECT 37.520 2.100 38.920 105.700 ;
    RECT 39.200 2.100 40.600 105.700 ;
    RECT 40.880 2.100 42.280 105.700 ;
    RECT 42.560 2.100 43.960 105.700 ;
    RECT 44.240 2.100 45.640 105.700 ;
    RECT 45.920 2.100 47.320 105.700 ;
    RECT 47.600 2.100 49.000 105.700 ;
    RECT 49.280 2.100 50.680 105.700 ;
    RECT 50.960 2.100 52.360 105.700 ;
    RECT 52.640 2.100 54.040 105.700 ;
    RECT 54.320 2.100 55.720 105.700 ;
    RECT 56.000 2.100 57.400 105.700 ;
    RECT 57.680 2.100 59.080 105.700 ;
    RECT 59.360 2.100 60.760 105.700 ;
    RECT 61.040 2.100 62.440 105.700 ;
    RECT 62.720 2.100 64.120 105.700 ;
    RECT 64.400 2.100 65.800 105.700 ;
    RECT 66.080 2.100 67.480 105.700 ;
    RECT 67.760 2.100 69.160 105.700 ;
    RECT 69.440 2.100 70.840 105.700 ;
    RECT 71.120 2.100 72.520 105.700 ;
    RECT 72.800 2.100 74.200 105.700 ;
    RECT 74.480 2.100 75.880 105.700 ;
    RECT 76.160 2.100 77.560 105.700 ;
    RECT 77.840 2.100 79.240 105.700 ;
    RECT 79.520 2.100 80.920 105.700 ;
    RECT 81.200 2.100 82.600 105.700 ;
    RECT 82.880 2.100 84.280 105.700 ;
    RECT 84.560 2.100 85.960 105.700 ;
    RECT 86.240 2.100 87.640 105.700 ;
    RECT 87.920 2.100 89.320 105.700 ;
    RECT 89.600 2.100 91.000 105.700 ;
    RECT 91.280 2.100 92.680 105.700 ;
    RECT 92.960 2.100 94.360 105.700 ;
    RECT 94.640 2.100 96.040 105.700 ;
    RECT 96.320 2.100 97.720 105.700 ;
    RECT 98.000 2.100 99.400 105.700 ;
    RECT 99.680 2.100 101.080 105.700 ;
    RECT 101.360 2.100 102.760 105.700 ;
    RECT 103.040 2.100 104.440 105.700 ;
    RECT 104.720 2.100 106.120 105.700 ;
    RECT 106.400 2.100 107.800 105.700 ;
    RECT 108.080 2.100 109.480 105.700 ;
    RECT 109.760 2.100 111.160 105.700 ;
    RECT 111.440 2.100 112.840 105.700 ;
    RECT 113.120 2.100 114.520 105.700 ;
    RECT 114.800 2.100 116.200 105.700 ;
    RECT 116.480 2.100 117.880 105.700 ;
    RECT 118.160 2.100 119.560 105.700 ;
    RECT 119.840 2.100 121.240 105.700 ;
    RECT 121.520 2.100 122.920 105.700 ;
    RECT 123.200 2.100 124.600 105.700 ;
    RECT 124.880 2.100 126.280 105.700 ;
    RECT 126.560 2.100 127.960 105.700 ;
    RECT 128.240 2.100 129.640 105.700 ;
    RECT 129.920 2.100 131.320 105.700 ;
    RECT 131.600 2.100 133.000 105.700 ;
    RECT 133.280 2.100 134.680 105.700 ;
    RECT 134.960 2.100 136.360 105.700 ;
    RECT 136.640 2.100 138.040 105.700 ;
    RECT 138.320 2.100 139.720 105.700 ;
    RECT 140.000 2.100 141.400 105.700 ;
    RECT 141.680 2.100 143.080 105.700 ;
    RECT 143.360 2.100 144.760 105.700 ;
    RECT 145.040 2.100 146.440 105.700 ;
    RECT 146.720 2.100 148.120 105.700 ;
    RECT 148.400 2.100 149.800 105.700 ;
    RECT 150.080 2.100 152.190 105.700 ;
    LAYER OVERLAP ;
    RECT 0 0 152.190 107.800 ;
  END
END fakeram45_1024x32

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_512x64
  FOREIGN fakeram45_512x64 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 152.570 BY 113.400 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.785 0.070 8.855 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.985 0.070 13.055 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.505 0.070 15.575 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.345 0.070 16.415 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.185 0.070 17.255 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.605 0.070 17.675 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.025 0.070 18.095 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.545 0.070 20.615 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.225 0.070 22.295 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.905 0.070 23.975 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.425 0.070 26.495 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.685 0.070 27.755 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.105 0.070 28.175 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END w_mask_in[63]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.825 0.070 34.895 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.505 0.070 36.575 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.185 0.070 38.255 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.325 0.070 45.395 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.745 0.070 45.815 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.585 0.070 46.655 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.265 0.070 48.335 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.945 0.070 50.015 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.785 0.070 50.855 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.205 0.070 51.275 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.625 0.070 51.695 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.045 0.070 52.115 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.305 0.070 53.375 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.145 0.070 54.215 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.985 0.070 55.055 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.825 0.070 55.895 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.665 0.070 56.735 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.085 0.070 57.155 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.505 0.070 57.575 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.345 0.070 58.415 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.765 0.070 58.835 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.185 0.070 59.255 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.605 0.070 59.675 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.025 0.070 60.095 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.445 0.070 60.515 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.865 0.070 60.935 ;
    END
  END rd_out[63]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.745 0.070 66.815 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.165 0.070 67.235 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.585 0.070 67.655 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.425 0.070 68.495 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.845 0.070 68.915 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.265 0.070 69.335 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.685 0.070 69.755 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.105 0.070 70.175 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.945 0.070 71.015 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.785 0.070 71.855 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.205 0.070 72.275 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.625 0.070 72.695 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.465 0.070 73.535 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.305 0.070 74.375 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.725 0.070 74.795 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.145 0.070 75.215 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.405 0.070 76.475 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.825 0.070 76.895 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.245 0.070 77.315 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.665 0.070 77.735 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.085 0.070 78.155 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.505 0.070 78.575 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.925 0.070 78.995 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.345 0.070 79.415 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.185 0.070 80.255 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.605 0.070 80.675 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.025 0.070 81.095 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.445 0.070 81.515 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.285 0.070 82.355 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.705 0.070 82.775 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.125 0.070 83.195 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.545 0.070 83.615 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.965 0.070 84.035 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.385 0.070 84.455 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.225 0.070 85.295 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.065 0.070 86.135 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.485 0.070 86.555 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.905 0.070 86.975 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.325 0.070 87.395 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.745 0.070 87.815 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.165 0.070 88.235 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.585 0.070 88.655 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.005 0.070 89.075 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.425 0.070 89.495 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.845 0.070 89.915 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.265 0.070 90.335 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.685 0.070 90.755 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.105 0.070 91.175 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.525 0.070 91.595 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.945 0.070 92.015 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.365 0.070 92.435 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.785 0.070 92.855 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.205 0.070 93.275 ;
    END
  END wd_in[63]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.085 0.070 99.155 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.505 0.070 99.575 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.925 0.070 99.995 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.345 0.070 100.415 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.765 0.070 100.835 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.185 0.070 101.255 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.605 0.070 101.675 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.025 0.070 102.095 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.445 0.070 102.515 ;
    END
  END addr_in[8]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.325 0.070 108.395 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.745 0.070 108.815 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.165 0.070 109.235 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 111.300 ;
      RECT 5.320 2.100 5.600 111.300 ;
      RECT 8.680 2.100 8.960 111.300 ;
      RECT 12.040 2.100 12.320 111.300 ;
      RECT 15.400 2.100 15.680 111.300 ;
      RECT 18.760 2.100 19.040 111.300 ;
      RECT 22.120 2.100 22.400 111.300 ;
      RECT 25.480 2.100 25.760 111.300 ;
      RECT 28.840 2.100 29.120 111.300 ;
      RECT 32.200 2.100 32.480 111.300 ;
      RECT 35.560 2.100 35.840 111.300 ;
      RECT 38.920 2.100 39.200 111.300 ;
      RECT 42.280 2.100 42.560 111.300 ;
      RECT 45.640 2.100 45.920 111.300 ;
      RECT 49.000 2.100 49.280 111.300 ;
      RECT 52.360 2.100 52.640 111.300 ;
      RECT 55.720 2.100 56.000 111.300 ;
      RECT 59.080 2.100 59.360 111.300 ;
      RECT 62.440 2.100 62.720 111.300 ;
      RECT 65.800 2.100 66.080 111.300 ;
      RECT 69.160 2.100 69.440 111.300 ;
      RECT 72.520 2.100 72.800 111.300 ;
      RECT 75.880 2.100 76.160 111.300 ;
      RECT 79.240 2.100 79.520 111.300 ;
      RECT 82.600 2.100 82.880 111.300 ;
      RECT 85.960 2.100 86.240 111.300 ;
      RECT 89.320 2.100 89.600 111.300 ;
      RECT 92.680 2.100 92.960 111.300 ;
      RECT 96.040 2.100 96.320 111.300 ;
      RECT 99.400 2.100 99.680 111.300 ;
      RECT 102.760 2.100 103.040 111.300 ;
      RECT 106.120 2.100 106.400 111.300 ;
      RECT 109.480 2.100 109.760 111.300 ;
      RECT 112.840 2.100 113.120 111.300 ;
      RECT 116.200 2.100 116.480 111.300 ;
      RECT 119.560 2.100 119.840 111.300 ;
      RECT 122.920 2.100 123.200 111.300 ;
      RECT 126.280 2.100 126.560 111.300 ;
      RECT 129.640 2.100 129.920 111.300 ;
      RECT 133.000 2.100 133.280 111.300 ;
      RECT 136.360 2.100 136.640 111.300 ;
      RECT 139.720 2.100 140.000 111.300 ;
      RECT 143.080 2.100 143.360 111.300 ;
      RECT 146.440 2.100 146.720 111.300 ;
      RECT 149.800 2.100 150.080 111.300 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 111.300 ;
      RECT 7.000 2.100 7.280 111.300 ;
      RECT 10.360 2.100 10.640 111.300 ;
      RECT 13.720 2.100 14.000 111.300 ;
      RECT 17.080 2.100 17.360 111.300 ;
      RECT 20.440 2.100 20.720 111.300 ;
      RECT 23.800 2.100 24.080 111.300 ;
      RECT 27.160 2.100 27.440 111.300 ;
      RECT 30.520 2.100 30.800 111.300 ;
      RECT 33.880 2.100 34.160 111.300 ;
      RECT 37.240 2.100 37.520 111.300 ;
      RECT 40.600 2.100 40.880 111.300 ;
      RECT 43.960 2.100 44.240 111.300 ;
      RECT 47.320 2.100 47.600 111.300 ;
      RECT 50.680 2.100 50.960 111.300 ;
      RECT 54.040 2.100 54.320 111.300 ;
      RECT 57.400 2.100 57.680 111.300 ;
      RECT 60.760 2.100 61.040 111.300 ;
      RECT 64.120 2.100 64.400 111.300 ;
      RECT 67.480 2.100 67.760 111.300 ;
      RECT 70.840 2.100 71.120 111.300 ;
      RECT 74.200 2.100 74.480 111.300 ;
      RECT 77.560 2.100 77.840 111.300 ;
      RECT 80.920 2.100 81.200 111.300 ;
      RECT 84.280 2.100 84.560 111.300 ;
      RECT 87.640 2.100 87.920 111.300 ;
      RECT 91.000 2.100 91.280 111.300 ;
      RECT 94.360 2.100 94.640 111.300 ;
      RECT 97.720 2.100 98.000 111.300 ;
      RECT 101.080 2.100 101.360 111.300 ;
      RECT 104.440 2.100 104.720 111.300 ;
      RECT 107.800 2.100 108.080 111.300 ;
      RECT 111.160 2.100 111.440 111.300 ;
      RECT 114.520 2.100 114.800 111.300 ;
      RECT 117.880 2.100 118.160 111.300 ;
      RECT 121.240 2.100 121.520 111.300 ;
      RECT 124.600 2.100 124.880 111.300 ;
      RECT 127.960 2.100 128.240 111.300 ;
      RECT 131.320 2.100 131.600 111.300 ;
      RECT 134.680 2.100 134.960 111.300 ;
      RECT 138.040 2.100 138.320 111.300 ;
      RECT 141.400 2.100 141.680 111.300 ;
      RECT 144.760 2.100 145.040 111.300 ;
      RECT 148.120 2.100 148.400 111.300 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 152.570 113.400 ;
    LAYER metal2 ;
    RECT 0 0 152.570 113.400 ;
    LAYER metal3 ;
    RECT 0.070 0 152.570 113.400 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.485 ;
    RECT 0 2.555 0.070 2.905 ;
    RECT 0 2.975 0.070 3.325 ;
    RECT 0 3.395 0.070 3.745 ;
    RECT 0 3.815 0.070 4.165 ;
    RECT 0 4.235 0.070 4.585 ;
    RECT 0 4.655 0.070 5.005 ;
    RECT 0 5.075 0.070 5.425 ;
    RECT 0 5.495 0.070 5.845 ;
    RECT 0 5.915 0.070 6.265 ;
    RECT 0 6.335 0.070 6.685 ;
    RECT 0 6.755 0.070 7.105 ;
    RECT 0 7.175 0.070 7.525 ;
    RECT 0 7.595 0.070 7.945 ;
    RECT 0 8.015 0.070 8.365 ;
    RECT 0 8.435 0.070 8.785 ;
    RECT 0 8.855 0.070 9.205 ;
    RECT 0 9.275 0.070 9.625 ;
    RECT 0 9.695 0.070 10.045 ;
    RECT 0 10.115 0.070 10.465 ;
    RECT 0 10.535 0.070 10.885 ;
    RECT 0 10.955 0.070 11.305 ;
    RECT 0 11.375 0.070 11.725 ;
    RECT 0 11.795 0.070 12.145 ;
    RECT 0 12.215 0.070 12.565 ;
    RECT 0 12.635 0.070 12.985 ;
    RECT 0 13.055 0.070 13.405 ;
    RECT 0 13.475 0.070 13.825 ;
    RECT 0 13.895 0.070 14.245 ;
    RECT 0 14.315 0.070 14.665 ;
    RECT 0 14.735 0.070 15.085 ;
    RECT 0 15.155 0.070 15.505 ;
    RECT 0 15.575 0.070 15.925 ;
    RECT 0 15.995 0.070 16.345 ;
    RECT 0 16.415 0.070 16.765 ;
    RECT 0 16.835 0.070 17.185 ;
    RECT 0 17.255 0.070 17.605 ;
    RECT 0 17.675 0.070 18.025 ;
    RECT 0 18.095 0.070 18.445 ;
    RECT 0 18.515 0.070 18.865 ;
    RECT 0 18.935 0.070 19.285 ;
    RECT 0 19.355 0.070 19.705 ;
    RECT 0 19.775 0.070 20.125 ;
    RECT 0 20.195 0.070 20.545 ;
    RECT 0 20.615 0.070 20.965 ;
    RECT 0 21.035 0.070 21.385 ;
    RECT 0 21.455 0.070 21.805 ;
    RECT 0 21.875 0.070 22.225 ;
    RECT 0 22.295 0.070 22.645 ;
    RECT 0 22.715 0.070 23.065 ;
    RECT 0 23.135 0.070 23.485 ;
    RECT 0 23.555 0.070 23.905 ;
    RECT 0 23.975 0.070 24.325 ;
    RECT 0 24.395 0.070 24.745 ;
    RECT 0 24.815 0.070 25.165 ;
    RECT 0 25.235 0.070 25.585 ;
    RECT 0 25.655 0.070 26.005 ;
    RECT 0 26.075 0.070 26.425 ;
    RECT 0 26.495 0.070 26.845 ;
    RECT 0 26.915 0.070 27.265 ;
    RECT 0 27.335 0.070 27.685 ;
    RECT 0 27.755 0.070 28.105 ;
    RECT 0 28.175 0.070 28.525 ;
    RECT 0 28.595 0.070 34.405 ;
    RECT 0 34.475 0.070 34.825 ;
    RECT 0 34.895 0.070 35.245 ;
    RECT 0 35.315 0.070 35.665 ;
    RECT 0 35.735 0.070 36.085 ;
    RECT 0 36.155 0.070 36.505 ;
    RECT 0 36.575 0.070 36.925 ;
    RECT 0 36.995 0.070 37.345 ;
    RECT 0 37.415 0.070 37.765 ;
    RECT 0 37.835 0.070 38.185 ;
    RECT 0 38.255 0.070 38.605 ;
    RECT 0 38.675 0.070 39.025 ;
    RECT 0 39.095 0.070 39.445 ;
    RECT 0 39.515 0.070 39.865 ;
    RECT 0 39.935 0.070 40.285 ;
    RECT 0 40.355 0.070 40.705 ;
    RECT 0 40.775 0.070 41.125 ;
    RECT 0 41.195 0.070 41.545 ;
    RECT 0 41.615 0.070 41.965 ;
    RECT 0 42.035 0.070 42.385 ;
    RECT 0 42.455 0.070 42.805 ;
    RECT 0 42.875 0.070 43.225 ;
    RECT 0 43.295 0.070 43.645 ;
    RECT 0 43.715 0.070 44.065 ;
    RECT 0 44.135 0.070 44.485 ;
    RECT 0 44.555 0.070 44.905 ;
    RECT 0 44.975 0.070 45.325 ;
    RECT 0 45.395 0.070 45.745 ;
    RECT 0 45.815 0.070 46.165 ;
    RECT 0 46.235 0.070 46.585 ;
    RECT 0 46.655 0.070 47.005 ;
    RECT 0 47.075 0.070 47.425 ;
    RECT 0 47.495 0.070 47.845 ;
    RECT 0 47.915 0.070 48.265 ;
    RECT 0 48.335 0.070 48.685 ;
    RECT 0 48.755 0.070 49.105 ;
    RECT 0 49.175 0.070 49.525 ;
    RECT 0 49.595 0.070 49.945 ;
    RECT 0 50.015 0.070 50.365 ;
    RECT 0 50.435 0.070 50.785 ;
    RECT 0 50.855 0.070 51.205 ;
    RECT 0 51.275 0.070 51.625 ;
    RECT 0 51.695 0.070 52.045 ;
    RECT 0 52.115 0.070 52.465 ;
    RECT 0 52.535 0.070 52.885 ;
    RECT 0 52.955 0.070 53.305 ;
    RECT 0 53.375 0.070 53.725 ;
    RECT 0 53.795 0.070 54.145 ;
    RECT 0 54.215 0.070 54.565 ;
    RECT 0 54.635 0.070 54.985 ;
    RECT 0 55.055 0.070 55.405 ;
    RECT 0 55.475 0.070 55.825 ;
    RECT 0 55.895 0.070 56.245 ;
    RECT 0 56.315 0.070 56.665 ;
    RECT 0 56.735 0.070 57.085 ;
    RECT 0 57.155 0.070 57.505 ;
    RECT 0 57.575 0.070 57.925 ;
    RECT 0 57.995 0.070 58.345 ;
    RECT 0 58.415 0.070 58.765 ;
    RECT 0 58.835 0.070 59.185 ;
    RECT 0 59.255 0.070 59.605 ;
    RECT 0 59.675 0.070 60.025 ;
    RECT 0 60.095 0.070 60.445 ;
    RECT 0 60.515 0.070 60.865 ;
    RECT 0 60.935 0.070 66.745 ;
    RECT 0 66.815 0.070 67.165 ;
    RECT 0 67.235 0.070 67.585 ;
    RECT 0 67.655 0.070 68.005 ;
    RECT 0 68.075 0.070 68.425 ;
    RECT 0 68.495 0.070 68.845 ;
    RECT 0 68.915 0.070 69.265 ;
    RECT 0 69.335 0.070 69.685 ;
    RECT 0 69.755 0.070 70.105 ;
    RECT 0 70.175 0.070 70.525 ;
    RECT 0 70.595 0.070 70.945 ;
    RECT 0 71.015 0.070 71.365 ;
    RECT 0 71.435 0.070 71.785 ;
    RECT 0 71.855 0.070 72.205 ;
    RECT 0 72.275 0.070 72.625 ;
    RECT 0 72.695 0.070 73.045 ;
    RECT 0 73.115 0.070 73.465 ;
    RECT 0 73.535 0.070 73.885 ;
    RECT 0 73.955 0.070 74.305 ;
    RECT 0 74.375 0.070 74.725 ;
    RECT 0 74.795 0.070 75.145 ;
    RECT 0 75.215 0.070 75.565 ;
    RECT 0 75.635 0.070 75.985 ;
    RECT 0 76.055 0.070 76.405 ;
    RECT 0 76.475 0.070 76.825 ;
    RECT 0 76.895 0.070 77.245 ;
    RECT 0 77.315 0.070 77.665 ;
    RECT 0 77.735 0.070 78.085 ;
    RECT 0 78.155 0.070 78.505 ;
    RECT 0 78.575 0.070 78.925 ;
    RECT 0 78.995 0.070 79.345 ;
    RECT 0 79.415 0.070 79.765 ;
    RECT 0 79.835 0.070 80.185 ;
    RECT 0 80.255 0.070 80.605 ;
    RECT 0 80.675 0.070 81.025 ;
    RECT 0 81.095 0.070 81.445 ;
    RECT 0 81.515 0.070 81.865 ;
    RECT 0 81.935 0.070 82.285 ;
    RECT 0 82.355 0.070 82.705 ;
    RECT 0 82.775 0.070 83.125 ;
    RECT 0 83.195 0.070 83.545 ;
    RECT 0 83.615 0.070 83.965 ;
    RECT 0 84.035 0.070 84.385 ;
    RECT 0 84.455 0.070 84.805 ;
    RECT 0 84.875 0.070 85.225 ;
    RECT 0 85.295 0.070 85.645 ;
    RECT 0 85.715 0.070 86.065 ;
    RECT 0 86.135 0.070 86.485 ;
    RECT 0 86.555 0.070 86.905 ;
    RECT 0 86.975 0.070 87.325 ;
    RECT 0 87.395 0.070 87.745 ;
    RECT 0 87.815 0.070 88.165 ;
    RECT 0 88.235 0.070 88.585 ;
    RECT 0 88.655 0.070 89.005 ;
    RECT 0 89.075 0.070 89.425 ;
    RECT 0 89.495 0.070 89.845 ;
    RECT 0 89.915 0.070 90.265 ;
    RECT 0 90.335 0.070 90.685 ;
    RECT 0 90.755 0.070 91.105 ;
    RECT 0 91.175 0.070 91.525 ;
    RECT 0 91.595 0.070 91.945 ;
    RECT 0 92.015 0.070 92.365 ;
    RECT 0 92.435 0.070 92.785 ;
    RECT 0 92.855 0.070 93.205 ;
    RECT 0 93.275 0.070 99.085 ;
    RECT 0 99.155 0.070 99.505 ;
    RECT 0 99.575 0.070 99.925 ;
    RECT 0 99.995 0.070 100.345 ;
    RECT 0 100.415 0.070 100.765 ;
    RECT 0 100.835 0.070 101.185 ;
    RECT 0 101.255 0.070 101.605 ;
    RECT 0 101.675 0.070 102.025 ;
    RECT 0 102.095 0.070 102.445 ;
    RECT 0 102.515 0.070 108.325 ;
    RECT 0 108.395 0.070 108.745 ;
    RECT 0 108.815 0.070 109.165 ;
    RECT 0 109.235 0.070 113.400 ;
    LAYER metal4 ;
    RECT 0 0 152.570 2.100 ;
    RECT 0 111.300 152.570 113.400 ;
    RECT 0.000 2.100 1.960 111.300 ;
    RECT 2.240 2.100 3.640 111.300 ;
    RECT 3.920 2.100 5.320 111.300 ;
    RECT 5.600 2.100 7.000 111.300 ;
    RECT 7.280 2.100 8.680 111.300 ;
    RECT 8.960 2.100 10.360 111.300 ;
    RECT 10.640 2.100 12.040 111.300 ;
    RECT 12.320 2.100 13.720 111.300 ;
    RECT 14.000 2.100 15.400 111.300 ;
    RECT 15.680 2.100 17.080 111.300 ;
    RECT 17.360 2.100 18.760 111.300 ;
    RECT 19.040 2.100 20.440 111.300 ;
    RECT 20.720 2.100 22.120 111.300 ;
    RECT 22.400 2.100 23.800 111.300 ;
    RECT 24.080 2.100 25.480 111.300 ;
    RECT 25.760 2.100 27.160 111.300 ;
    RECT 27.440 2.100 28.840 111.300 ;
    RECT 29.120 2.100 30.520 111.300 ;
    RECT 30.800 2.100 32.200 111.300 ;
    RECT 32.480 2.100 33.880 111.300 ;
    RECT 34.160 2.100 35.560 111.300 ;
    RECT 35.840 2.100 37.240 111.300 ;
    RECT 37.520 2.100 38.920 111.300 ;
    RECT 39.200 2.100 40.600 111.300 ;
    RECT 40.880 2.100 42.280 111.300 ;
    RECT 42.560 2.100 43.960 111.300 ;
    RECT 44.240 2.100 45.640 111.300 ;
    RECT 45.920 2.100 47.320 111.300 ;
    RECT 47.600 2.100 49.000 111.300 ;
    RECT 49.280 2.100 50.680 111.300 ;
    RECT 50.960 2.100 52.360 111.300 ;
    RECT 52.640 2.100 54.040 111.300 ;
    RECT 54.320 2.100 55.720 111.300 ;
    RECT 56.000 2.100 57.400 111.300 ;
    RECT 57.680 2.100 59.080 111.300 ;
    RECT 59.360 2.100 60.760 111.300 ;
    RECT 61.040 2.100 62.440 111.300 ;
    RECT 62.720 2.100 64.120 111.300 ;
    RECT 64.400 2.100 65.800 111.300 ;
    RECT 66.080 2.100 67.480 111.300 ;
    RECT 67.760 2.100 69.160 111.300 ;
    RECT 69.440 2.100 70.840 111.300 ;
    RECT 71.120 2.100 72.520 111.300 ;
    RECT 72.800 2.100 74.200 111.300 ;
    RECT 74.480 2.100 75.880 111.300 ;
    RECT 76.160 2.100 77.560 111.300 ;
    RECT 77.840 2.100 79.240 111.300 ;
    RECT 79.520 2.100 80.920 111.300 ;
    RECT 81.200 2.100 82.600 111.300 ;
    RECT 82.880 2.100 84.280 111.300 ;
    RECT 84.560 2.100 85.960 111.300 ;
    RECT 86.240 2.100 87.640 111.300 ;
    RECT 87.920 2.100 89.320 111.300 ;
    RECT 89.600 2.100 91.000 111.300 ;
    RECT 91.280 2.100 92.680 111.300 ;
    RECT 92.960 2.100 94.360 111.300 ;
    RECT 94.640 2.100 96.040 111.300 ;
    RECT 96.320 2.100 97.720 111.300 ;
    RECT 98.000 2.100 99.400 111.300 ;
    RECT 99.680 2.100 101.080 111.300 ;
    RECT 101.360 2.100 102.760 111.300 ;
    RECT 103.040 2.100 104.440 111.300 ;
    RECT 104.720 2.100 106.120 111.300 ;
    RECT 106.400 2.100 107.800 111.300 ;
    RECT 108.080 2.100 109.480 111.300 ;
    RECT 109.760 2.100 111.160 111.300 ;
    RECT 111.440 2.100 112.840 111.300 ;
    RECT 113.120 2.100 114.520 111.300 ;
    RECT 114.800 2.100 116.200 111.300 ;
    RECT 116.480 2.100 117.880 111.300 ;
    RECT 118.160 2.100 119.560 111.300 ;
    RECT 119.840 2.100 121.240 111.300 ;
    RECT 121.520 2.100 122.920 111.300 ;
    RECT 123.200 2.100 124.600 111.300 ;
    RECT 124.880 2.100 126.280 111.300 ;
    RECT 126.560 2.100 127.960 111.300 ;
    RECT 128.240 2.100 129.640 111.300 ;
    RECT 129.920 2.100 131.320 111.300 ;
    RECT 131.600 2.100 133.000 111.300 ;
    RECT 133.280 2.100 134.680 111.300 ;
    RECT 134.960 2.100 136.360 111.300 ;
    RECT 136.640 2.100 138.040 111.300 ;
    RECT 138.320 2.100 139.720 111.300 ;
    RECT 140.000 2.100 141.400 111.300 ;
    RECT 141.680 2.100 143.080 111.300 ;
    RECT 143.360 2.100 144.760 111.300 ;
    RECT 145.040 2.100 146.440 111.300 ;
    RECT 146.720 2.100 148.120 111.300 ;
    RECT 148.400 2.100 149.800 111.300 ;
    RECT 150.080 2.100 152.570 111.300 ;
    LAYER OVERLAP ;
    RECT 0 0 152.570 113.400 ;
  END
END fakeram45_512x64

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_256x96
  FOREIGN fakeram45_256x96 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 115.140 BY 119.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.275 0.070 2.345 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.695 0.070 2.765 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.115 0.070 3.185 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.535 0.070 3.605 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.955 0.070 4.025 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.375 0.070 4.445 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.795 0.070 4.865 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.215 0.070 5.285 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.635 0.070 5.705 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.055 0.070 6.125 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.475 0.070 6.545 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.895 0.070 6.965 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.315 0.070 7.385 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.735 0.070 7.805 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.155 0.070 8.225 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.575 0.070 8.645 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.785 0.070 8.855 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.995 0.070 9.065 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.415 0.070 9.485 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.835 0.070 9.905 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.255 0.070 10.325 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.675 0.070 10.745 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.095 0.070 11.165 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.515 0.070 11.585 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.935 0.070 12.005 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.355 0.070 12.425 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.775 0.070 12.845 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.985 0.070 13.055 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.195 0.070 13.265 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.615 0.070 13.685 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.035 0.070 14.105 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.455 0.070 14.525 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.875 0.070 14.945 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.295 0.070 15.365 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.505 0.070 15.575 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.715 0.070 15.785 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.135 0.070 16.205 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.345 0.070 16.415 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.555 0.070 16.625 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.975 0.070 17.045 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.185 0.070 17.255 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.395 0.070 17.465 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.605 0.070 17.675 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.815 0.070 17.885 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.025 0.070 18.095 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.235 0.070 18.305 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.655 0.070 18.725 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.075 0.070 19.145 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.495 0.070 19.565 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.915 0.070 19.985 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.335 0.070 20.405 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.545 0.070 20.615 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.755 0.070 20.825 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.175 0.070 21.245 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.595 0.070 21.665 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.015 0.070 22.085 ;
    END
  END w_mask_in[95]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.825 0.070 34.895 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.035 0.070 35.105 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.455 0.070 35.525 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.875 0.070 35.945 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.295 0.070 36.365 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.505 0.070 36.575 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.715 0.070 36.785 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.135 0.070 37.205 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.555 0.070 37.625 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.975 0.070 38.045 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.185 0.070 38.255 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.395 0.070 38.465 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.815 0.070 38.885 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.235 0.070 39.305 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.655 0.070 39.725 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.075 0.070 40.145 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.495 0.070 40.565 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.915 0.070 40.985 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.335 0.070 41.405 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.755 0.070 41.825 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.175 0.070 42.245 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.595 0.070 42.665 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.015 0.070 43.085 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.435 0.070 43.505 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.855 0.070 43.925 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.275 0.070 44.345 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.695 0.070 44.765 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.115 0.070 45.185 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.325 0.070 45.395 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.535 0.070 45.605 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.745 0.070 45.815 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.955 0.070 46.025 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.375 0.070 46.445 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.585 0.070 46.655 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.795 0.070 46.865 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.215 0.070 47.285 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.635 0.070 47.705 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.055 0.070 48.125 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.265 0.070 48.335 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.475 0.070 48.545 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.895 0.070 48.965 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.315 0.070 49.385 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.735 0.070 49.805 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.945 0.070 50.015 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.155 0.070 50.225 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.575 0.070 50.645 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.785 0.070 50.855 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.995 0.070 51.065 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.205 0.070 51.275 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.415 0.070 51.485 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.625 0.070 51.695 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.835 0.070 51.905 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.045 0.070 52.115 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.255 0.070 52.325 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.675 0.070 52.745 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.095 0.070 53.165 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.305 0.070 53.375 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.515 0.070 53.585 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.935 0.070 54.005 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.145 0.070 54.215 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.355 0.070 54.425 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.775 0.070 54.845 ;
    END
  END rd_out[95]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.585 0.070 67.655 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.795 0.070 67.865 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.215 0.070 68.285 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.425 0.070 68.495 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.635 0.070 68.705 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.845 0.070 68.915 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.055 0.070 69.125 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.265 0.070 69.335 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.475 0.070 69.545 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.685 0.070 69.755 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.895 0.070 69.965 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.105 0.070 70.175 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.315 0.070 70.385 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.735 0.070 70.805 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.945 0.070 71.015 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.155 0.070 71.225 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.575 0.070 71.645 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.785 0.070 71.855 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.995 0.070 72.065 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.205 0.070 72.275 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.415 0.070 72.485 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.625 0.070 72.695 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.835 0.070 72.905 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.255 0.070 73.325 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.465 0.070 73.535 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.675 0.070 73.745 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.095 0.070 74.165 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.305 0.070 74.375 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.515 0.070 74.585 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.725 0.070 74.795 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.935 0.070 75.005 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.145 0.070 75.215 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.355 0.070 75.425 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.775 0.070 75.845 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.195 0.070 76.265 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.405 0.070 76.475 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.615 0.070 76.685 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.825 0.070 76.895 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.035 0.070 77.105 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.245 0.070 77.315 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.455 0.070 77.525 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.665 0.070 77.735 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.875 0.070 77.945 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.085 0.070 78.155 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.295 0.070 78.365 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.505 0.070 78.575 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.715 0.070 78.785 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.925 0.070 78.995 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.135 0.070 79.205 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.345 0.070 79.415 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.555 0.070 79.625 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.975 0.070 80.045 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.185 0.070 80.255 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.395 0.070 80.465 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.605 0.070 80.675 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.815 0.070 80.885 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.025 0.070 81.095 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.235 0.070 81.305 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.445 0.070 81.515 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.655 0.070 81.725 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.075 0.070 82.145 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.285 0.070 82.355 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.495 0.070 82.565 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.705 0.070 82.775 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.915 0.070 82.985 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.125 0.070 83.195 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.335 0.070 83.405 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.545 0.070 83.615 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.755 0.070 83.825 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.965 0.070 84.035 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.175 0.070 84.245 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.385 0.070 84.455 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.595 0.070 84.665 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.015 0.070 85.085 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.225 0.070 85.295 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.435 0.070 85.505 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.855 0.070 85.925 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.065 0.070 86.135 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.275 0.070 86.345 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.485 0.070 86.555 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.695 0.070 86.765 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.905 0.070 86.975 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.115 0.070 87.185 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.325 0.070 87.395 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.535 0.070 87.605 ;
    END
  END wd_in[95]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.345 0.070 100.415 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.555 0.070 100.625 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.765 0.070 100.835 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.975 0.070 101.045 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.185 0.070 101.255 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.395 0.070 101.465 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.605 0.070 101.675 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.815 0.070 101.885 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.625 0.070 114.695 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.835 0.070 114.905 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.045 0.070 115.115 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 116.900 ;
      RECT 5.320 2.100 5.600 116.900 ;
      RECT 8.680 2.100 8.960 116.900 ;
      RECT 12.040 2.100 12.320 116.900 ;
      RECT 15.400 2.100 15.680 116.900 ;
      RECT 18.760 2.100 19.040 116.900 ;
      RECT 22.120 2.100 22.400 116.900 ;
      RECT 25.480 2.100 25.760 116.900 ;
      RECT 28.840 2.100 29.120 116.900 ;
      RECT 32.200 2.100 32.480 116.900 ;
      RECT 35.560 2.100 35.840 116.900 ;
      RECT 38.920 2.100 39.200 116.900 ;
      RECT 42.280 2.100 42.560 116.900 ;
      RECT 45.640 2.100 45.920 116.900 ;
      RECT 49.000 2.100 49.280 116.900 ;
      RECT 52.360 2.100 52.640 116.900 ;
      RECT 55.720 2.100 56.000 116.900 ;
      RECT 59.080 2.100 59.360 116.900 ;
      RECT 62.440 2.100 62.720 116.900 ;
      RECT 65.800 2.100 66.080 116.900 ;
      RECT 69.160 2.100 69.440 116.900 ;
      RECT 72.520 2.100 72.800 116.900 ;
      RECT 75.880 2.100 76.160 116.900 ;
      RECT 79.240 2.100 79.520 116.900 ;
      RECT 82.600 2.100 82.880 116.900 ;
      RECT 85.960 2.100 86.240 116.900 ;
      RECT 89.320 2.100 89.600 116.900 ;
      RECT 92.680 2.100 92.960 116.900 ;
      RECT 96.040 2.100 96.320 116.900 ;
      RECT 99.400 2.100 99.680 116.900 ;
      RECT 102.760 2.100 103.040 116.900 ;
      RECT 106.120 2.100 106.400 116.900 ;
      RECT 109.480 2.100 109.760 116.900 ;
      RECT 112.840 2.100 113.120 116.900 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 116.900 ;
      RECT 7.000 2.100 7.280 116.900 ;
      RECT 10.360 2.100 10.640 116.900 ;
      RECT 13.720 2.100 14.000 116.900 ;
      RECT 17.080 2.100 17.360 116.900 ;
      RECT 20.440 2.100 20.720 116.900 ;
      RECT 23.800 2.100 24.080 116.900 ;
      RECT 27.160 2.100 27.440 116.900 ;
      RECT 30.520 2.100 30.800 116.900 ;
      RECT 33.880 2.100 34.160 116.900 ;
      RECT 37.240 2.100 37.520 116.900 ;
      RECT 40.600 2.100 40.880 116.900 ;
      RECT 43.960 2.100 44.240 116.900 ;
      RECT 47.320 2.100 47.600 116.900 ;
      RECT 50.680 2.100 50.960 116.900 ;
      RECT 54.040 2.100 54.320 116.900 ;
      RECT 57.400 2.100 57.680 116.900 ;
      RECT 60.760 2.100 61.040 116.900 ;
      RECT 64.120 2.100 64.400 116.900 ;
      RECT 67.480 2.100 67.760 116.900 ;
      RECT 70.840 2.100 71.120 116.900 ;
      RECT 74.200 2.100 74.480 116.900 ;
      RECT 77.560 2.100 77.840 116.900 ;
      RECT 80.920 2.100 81.200 116.900 ;
      RECT 84.280 2.100 84.560 116.900 ;
      RECT 87.640 2.100 87.920 116.900 ;
      RECT 91.000 2.100 91.280 116.900 ;
      RECT 94.360 2.100 94.640 116.900 ;
      RECT 97.720 2.100 98.000 116.900 ;
      RECT 101.080 2.100 101.360 116.900 ;
      RECT 104.440 2.100 104.720 116.900 ;
      RECT 107.800 2.100 108.080 116.900 ;
      RECT 111.160 2.100 111.440 116.900 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 115.140 119.000 ;
    LAYER metal2 ;
    RECT 0 0 115.140 119.000 ;
    LAYER metal3 ;
    RECT 0.070 0 115.140 119.000 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.275 ;
    RECT 0 2.345 0.070 2.485 ;
    RECT 0 2.555 0.070 2.695 ;
    RECT 0 2.765 0.070 2.905 ;
    RECT 0 2.975 0.070 3.115 ;
    RECT 0 3.185 0.070 3.325 ;
    RECT 0 3.395 0.070 3.535 ;
    RECT 0 3.605 0.070 3.745 ;
    RECT 0 3.815 0.070 3.955 ;
    RECT 0 4.025 0.070 4.165 ;
    RECT 0 4.235 0.070 4.375 ;
    RECT 0 4.445 0.070 4.585 ;
    RECT 0 4.655 0.070 4.795 ;
    RECT 0 4.865 0.070 5.005 ;
    RECT 0 5.075 0.070 5.215 ;
    RECT 0 5.285 0.070 5.425 ;
    RECT 0 5.495 0.070 5.635 ;
    RECT 0 5.705 0.070 5.845 ;
    RECT 0 5.915 0.070 6.055 ;
    RECT 0 6.125 0.070 6.265 ;
    RECT 0 6.335 0.070 6.475 ;
    RECT 0 6.545 0.070 6.685 ;
    RECT 0 6.755 0.070 6.895 ;
    RECT 0 6.965 0.070 7.105 ;
    RECT 0 7.175 0.070 7.315 ;
    RECT 0 7.385 0.070 7.525 ;
    RECT 0 7.595 0.070 7.735 ;
    RECT 0 7.805 0.070 7.945 ;
    RECT 0 8.015 0.070 8.155 ;
    RECT 0 8.225 0.070 8.365 ;
    RECT 0 8.435 0.070 8.575 ;
    RECT 0 8.645 0.070 8.785 ;
    RECT 0 8.855 0.070 8.995 ;
    RECT 0 9.065 0.070 9.205 ;
    RECT 0 9.275 0.070 9.415 ;
    RECT 0 9.485 0.070 9.625 ;
    RECT 0 9.695 0.070 9.835 ;
    RECT 0 9.905 0.070 10.045 ;
    RECT 0 10.115 0.070 10.255 ;
    RECT 0 10.325 0.070 10.465 ;
    RECT 0 10.535 0.070 10.675 ;
    RECT 0 10.745 0.070 10.885 ;
    RECT 0 10.955 0.070 11.095 ;
    RECT 0 11.165 0.070 11.305 ;
    RECT 0 11.375 0.070 11.515 ;
    RECT 0 11.585 0.070 11.725 ;
    RECT 0 11.795 0.070 11.935 ;
    RECT 0 12.005 0.070 12.145 ;
    RECT 0 12.215 0.070 12.355 ;
    RECT 0 12.425 0.070 12.565 ;
    RECT 0 12.635 0.070 12.775 ;
    RECT 0 12.845 0.070 12.985 ;
    RECT 0 13.055 0.070 13.195 ;
    RECT 0 13.265 0.070 13.405 ;
    RECT 0 13.475 0.070 13.615 ;
    RECT 0 13.685 0.070 13.825 ;
    RECT 0 13.895 0.070 14.035 ;
    RECT 0 14.105 0.070 14.245 ;
    RECT 0 14.315 0.070 14.455 ;
    RECT 0 14.525 0.070 14.665 ;
    RECT 0 14.735 0.070 14.875 ;
    RECT 0 14.945 0.070 15.085 ;
    RECT 0 15.155 0.070 15.295 ;
    RECT 0 15.365 0.070 15.505 ;
    RECT 0 15.575 0.070 15.715 ;
    RECT 0 15.785 0.070 15.925 ;
    RECT 0 15.995 0.070 16.135 ;
    RECT 0 16.205 0.070 16.345 ;
    RECT 0 16.415 0.070 16.555 ;
    RECT 0 16.625 0.070 16.765 ;
    RECT 0 16.835 0.070 16.975 ;
    RECT 0 17.045 0.070 17.185 ;
    RECT 0 17.255 0.070 17.395 ;
    RECT 0 17.465 0.070 17.605 ;
    RECT 0 17.675 0.070 17.815 ;
    RECT 0 17.885 0.070 18.025 ;
    RECT 0 18.095 0.070 18.235 ;
    RECT 0 18.305 0.070 18.445 ;
    RECT 0 18.515 0.070 18.655 ;
    RECT 0 18.725 0.070 18.865 ;
    RECT 0 18.935 0.070 19.075 ;
    RECT 0 19.145 0.070 19.285 ;
    RECT 0 19.355 0.070 19.495 ;
    RECT 0 19.565 0.070 19.705 ;
    RECT 0 19.775 0.070 19.915 ;
    RECT 0 19.985 0.070 20.125 ;
    RECT 0 20.195 0.070 20.335 ;
    RECT 0 20.405 0.070 20.545 ;
    RECT 0 20.615 0.070 20.755 ;
    RECT 0 20.825 0.070 20.965 ;
    RECT 0 21.035 0.070 21.175 ;
    RECT 0 21.245 0.070 21.385 ;
    RECT 0 21.455 0.070 21.595 ;
    RECT 0 21.665 0.070 21.805 ;
    RECT 0 21.875 0.070 22.015 ;
    RECT 0 22.085 0.070 34.825 ;
    RECT 0 34.895 0.070 35.035 ;
    RECT 0 35.105 0.070 35.245 ;
    RECT 0 35.315 0.070 35.455 ;
    RECT 0 35.525 0.070 35.665 ;
    RECT 0 35.735 0.070 35.875 ;
    RECT 0 35.945 0.070 36.085 ;
    RECT 0 36.155 0.070 36.295 ;
    RECT 0 36.365 0.070 36.505 ;
    RECT 0 36.575 0.070 36.715 ;
    RECT 0 36.785 0.070 36.925 ;
    RECT 0 36.995 0.070 37.135 ;
    RECT 0 37.205 0.070 37.345 ;
    RECT 0 37.415 0.070 37.555 ;
    RECT 0 37.625 0.070 37.765 ;
    RECT 0 37.835 0.070 37.975 ;
    RECT 0 38.045 0.070 38.185 ;
    RECT 0 38.255 0.070 38.395 ;
    RECT 0 38.465 0.070 38.605 ;
    RECT 0 38.675 0.070 38.815 ;
    RECT 0 38.885 0.070 39.025 ;
    RECT 0 39.095 0.070 39.235 ;
    RECT 0 39.305 0.070 39.445 ;
    RECT 0 39.515 0.070 39.655 ;
    RECT 0 39.725 0.070 39.865 ;
    RECT 0 39.935 0.070 40.075 ;
    RECT 0 40.145 0.070 40.285 ;
    RECT 0 40.355 0.070 40.495 ;
    RECT 0 40.565 0.070 40.705 ;
    RECT 0 40.775 0.070 40.915 ;
    RECT 0 40.985 0.070 41.125 ;
    RECT 0 41.195 0.070 41.335 ;
    RECT 0 41.405 0.070 41.545 ;
    RECT 0 41.615 0.070 41.755 ;
    RECT 0 41.825 0.070 41.965 ;
    RECT 0 42.035 0.070 42.175 ;
    RECT 0 42.245 0.070 42.385 ;
    RECT 0 42.455 0.070 42.595 ;
    RECT 0 42.665 0.070 42.805 ;
    RECT 0 42.875 0.070 43.015 ;
    RECT 0 43.085 0.070 43.225 ;
    RECT 0 43.295 0.070 43.435 ;
    RECT 0 43.505 0.070 43.645 ;
    RECT 0 43.715 0.070 43.855 ;
    RECT 0 43.925 0.070 44.065 ;
    RECT 0 44.135 0.070 44.275 ;
    RECT 0 44.345 0.070 44.485 ;
    RECT 0 44.555 0.070 44.695 ;
    RECT 0 44.765 0.070 44.905 ;
    RECT 0 44.975 0.070 45.115 ;
    RECT 0 45.185 0.070 45.325 ;
    RECT 0 45.395 0.070 45.535 ;
    RECT 0 45.605 0.070 45.745 ;
    RECT 0 45.815 0.070 45.955 ;
    RECT 0 46.025 0.070 46.165 ;
    RECT 0 46.235 0.070 46.375 ;
    RECT 0 46.445 0.070 46.585 ;
    RECT 0 46.655 0.070 46.795 ;
    RECT 0 46.865 0.070 47.005 ;
    RECT 0 47.075 0.070 47.215 ;
    RECT 0 47.285 0.070 47.425 ;
    RECT 0 47.495 0.070 47.635 ;
    RECT 0 47.705 0.070 47.845 ;
    RECT 0 47.915 0.070 48.055 ;
    RECT 0 48.125 0.070 48.265 ;
    RECT 0 48.335 0.070 48.475 ;
    RECT 0 48.545 0.070 48.685 ;
    RECT 0 48.755 0.070 48.895 ;
    RECT 0 48.965 0.070 49.105 ;
    RECT 0 49.175 0.070 49.315 ;
    RECT 0 49.385 0.070 49.525 ;
    RECT 0 49.595 0.070 49.735 ;
    RECT 0 49.805 0.070 49.945 ;
    RECT 0 50.015 0.070 50.155 ;
    RECT 0 50.225 0.070 50.365 ;
    RECT 0 50.435 0.070 50.575 ;
    RECT 0 50.645 0.070 50.785 ;
    RECT 0 50.855 0.070 50.995 ;
    RECT 0 51.065 0.070 51.205 ;
    RECT 0 51.275 0.070 51.415 ;
    RECT 0 51.485 0.070 51.625 ;
    RECT 0 51.695 0.070 51.835 ;
    RECT 0 51.905 0.070 52.045 ;
    RECT 0 52.115 0.070 52.255 ;
    RECT 0 52.325 0.070 52.465 ;
    RECT 0 52.535 0.070 52.675 ;
    RECT 0 52.745 0.070 52.885 ;
    RECT 0 52.955 0.070 53.095 ;
    RECT 0 53.165 0.070 53.305 ;
    RECT 0 53.375 0.070 53.515 ;
    RECT 0 53.585 0.070 53.725 ;
    RECT 0 53.795 0.070 53.935 ;
    RECT 0 54.005 0.070 54.145 ;
    RECT 0 54.215 0.070 54.355 ;
    RECT 0 54.425 0.070 54.565 ;
    RECT 0 54.635 0.070 54.775 ;
    RECT 0 54.845 0.070 67.585 ;
    RECT 0 67.655 0.070 67.795 ;
    RECT 0 67.865 0.070 68.005 ;
    RECT 0 68.075 0.070 68.215 ;
    RECT 0 68.285 0.070 68.425 ;
    RECT 0 68.495 0.070 68.635 ;
    RECT 0 68.705 0.070 68.845 ;
    RECT 0 68.915 0.070 69.055 ;
    RECT 0 69.125 0.070 69.265 ;
    RECT 0 69.335 0.070 69.475 ;
    RECT 0 69.545 0.070 69.685 ;
    RECT 0 69.755 0.070 69.895 ;
    RECT 0 69.965 0.070 70.105 ;
    RECT 0 70.175 0.070 70.315 ;
    RECT 0 70.385 0.070 70.525 ;
    RECT 0 70.595 0.070 70.735 ;
    RECT 0 70.805 0.070 70.945 ;
    RECT 0 71.015 0.070 71.155 ;
    RECT 0 71.225 0.070 71.365 ;
    RECT 0 71.435 0.070 71.575 ;
    RECT 0 71.645 0.070 71.785 ;
    RECT 0 71.855 0.070 71.995 ;
    RECT 0 72.065 0.070 72.205 ;
    RECT 0 72.275 0.070 72.415 ;
    RECT 0 72.485 0.070 72.625 ;
    RECT 0 72.695 0.070 72.835 ;
    RECT 0 72.905 0.070 73.045 ;
    RECT 0 73.115 0.070 73.255 ;
    RECT 0 73.325 0.070 73.465 ;
    RECT 0 73.535 0.070 73.675 ;
    RECT 0 73.745 0.070 73.885 ;
    RECT 0 73.955 0.070 74.095 ;
    RECT 0 74.165 0.070 74.305 ;
    RECT 0 74.375 0.070 74.515 ;
    RECT 0 74.585 0.070 74.725 ;
    RECT 0 74.795 0.070 74.935 ;
    RECT 0 75.005 0.070 75.145 ;
    RECT 0 75.215 0.070 75.355 ;
    RECT 0 75.425 0.070 75.565 ;
    RECT 0 75.635 0.070 75.775 ;
    RECT 0 75.845 0.070 75.985 ;
    RECT 0 76.055 0.070 76.195 ;
    RECT 0 76.265 0.070 76.405 ;
    RECT 0 76.475 0.070 76.615 ;
    RECT 0 76.685 0.070 76.825 ;
    RECT 0 76.895 0.070 77.035 ;
    RECT 0 77.105 0.070 77.245 ;
    RECT 0 77.315 0.070 77.455 ;
    RECT 0 77.525 0.070 77.665 ;
    RECT 0 77.735 0.070 77.875 ;
    RECT 0 77.945 0.070 78.085 ;
    RECT 0 78.155 0.070 78.295 ;
    RECT 0 78.365 0.070 78.505 ;
    RECT 0 78.575 0.070 78.715 ;
    RECT 0 78.785 0.070 78.925 ;
    RECT 0 78.995 0.070 79.135 ;
    RECT 0 79.205 0.070 79.345 ;
    RECT 0 79.415 0.070 79.555 ;
    RECT 0 79.625 0.070 79.765 ;
    RECT 0 79.835 0.070 79.975 ;
    RECT 0 80.045 0.070 80.185 ;
    RECT 0 80.255 0.070 80.395 ;
    RECT 0 80.465 0.070 80.605 ;
    RECT 0 80.675 0.070 80.815 ;
    RECT 0 80.885 0.070 81.025 ;
    RECT 0 81.095 0.070 81.235 ;
    RECT 0 81.305 0.070 81.445 ;
    RECT 0 81.515 0.070 81.655 ;
    RECT 0 81.725 0.070 81.865 ;
    RECT 0 81.935 0.070 82.075 ;
    RECT 0 82.145 0.070 82.285 ;
    RECT 0 82.355 0.070 82.495 ;
    RECT 0 82.565 0.070 82.705 ;
    RECT 0 82.775 0.070 82.915 ;
    RECT 0 82.985 0.070 83.125 ;
    RECT 0 83.195 0.070 83.335 ;
    RECT 0 83.405 0.070 83.545 ;
    RECT 0 83.615 0.070 83.755 ;
    RECT 0 83.825 0.070 83.965 ;
    RECT 0 84.035 0.070 84.175 ;
    RECT 0 84.245 0.070 84.385 ;
    RECT 0 84.455 0.070 84.595 ;
    RECT 0 84.665 0.070 84.805 ;
    RECT 0 84.875 0.070 85.015 ;
    RECT 0 85.085 0.070 85.225 ;
    RECT 0 85.295 0.070 85.435 ;
    RECT 0 85.505 0.070 85.645 ;
    RECT 0 85.715 0.070 85.855 ;
    RECT 0 85.925 0.070 86.065 ;
    RECT 0 86.135 0.070 86.275 ;
    RECT 0 86.345 0.070 86.485 ;
    RECT 0 86.555 0.070 86.695 ;
    RECT 0 86.765 0.070 86.905 ;
    RECT 0 86.975 0.070 87.115 ;
    RECT 0 87.185 0.070 87.325 ;
    RECT 0 87.395 0.070 87.535 ;
    RECT 0 87.605 0.070 100.345 ;
    RECT 0 100.415 0.070 100.555 ;
    RECT 0 100.625 0.070 100.765 ;
    RECT 0 100.835 0.070 100.975 ;
    RECT 0 101.045 0.070 101.185 ;
    RECT 0 101.255 0.070 101.395 ;
    RECT 0 101.465 0.070 101.605 ;
    RECT 0 101.675 0.070 101.815 ;
    RECT 0 101.885 0.070 114.625 ;
    RECT 0 114.695 0.070 114.835 ;
    RECT 0 114.905 0.070 115.045 ;
    RECT 0 115.115 0.070 119.000 ;
    LAYER metal4 ;
    RECT 0 0 115.140 2.100 ;
    RECT 0 116.900 115.140 119.000 ;
    RECT 0.000 2.100 1.960 116.900 ;
    RECT 2.240 2.100 3.640 116.900 ;
    RECT 3.920 2.100 5.320 116.900 ;
    RECT 5.600 2.100 7.000 116.900 ;
    RECT 7.280 2.100 8.680 116.900 ;
    RECT 8.960 2.100 10.360 116.900 ;
    RECT 10.640 2.100 12.040 116.900 ;
    RECT 12.320 2.100 13.720 116.900 ;
    RECT 14.000 2.100 15.400 116.900 ;
    RECT 15.680 2.100 17.080 116.900 ;
    RECT 17.360 2.100 18.760 116.900 ;
    RECT 19.040 2.100 20.440 116.900 ;
    RECT 20.720 2.100 22.120 116.900 ;
    RECT 22.400 2.100 23.800 116.900 ;
    RECT 24.080 2.100 25.480 116.900 ;
    RECT 25.760 2.100 27.160 116.900 ;
    RECT 27.440 2.100 28.840 116.900 ;
    RECT 29.120 2.100 30.520 116.900 ;
    RECT 30.800 2.100 32.200 116.900 ;
    RECT 32.480 2.100 33.880 116.900 ;
    RECT 34.160 2.100 35.560 116.900 ;
    RECT 35.840 2.100 37.240 116.900 ;
    RECT 37.520 2.100 38.920 116.900 ;
    RECT 39.200 2.100 40.600 116.900 ;
    RECT 40.880 2.100 42.280 116.900 ;
    RECT 42.560 2.100 43.960 116.900 ;
    RECT 44.240 2.100 45.640 116.900 ;
    RECT 45.920 2.100 47.320 116.900 ;
    RECT 47.600 2.100 49.000 116.900 ;
    RECT 49.280 2.100 50.680 116.900 ;
    RECT 50.960 2.100 52.360 116.900 ;
    RECT 52.640 2.100 54.040 116.900 ;
    RECT 54.320 2.100 55.720 116.900 ;
    RECT 56.000 2.100 57.400 116.900 ;
    RECT 57.680 2.100 59.080 116.900 ;
    RECT 59.360 2.100 60.760 116.900 ;
    RECT 61.040 2.100 62.440 116.900 ;
    RECT 62.720 2.100 64.120 116.900 ;
    RECT 64.400 2.100 65.800 116.900 ;
    RECT 66.080 2.100 67.480 116.900 ;
    RECT 67.760 2.100 69.160 116.900 ;
    RECT 69.440 2.100 70.840 116.900 ;
    RECT 71.120 2.100 72.520 116.900 ;
    RECT 72.800 2.100 74.200 116.900 ;
    RECT 74.480 2.100 75.880 116.900 ;
    RECT 76.160 2.100 77.560 116.900 ;
    RECT 77.840 2.100 79.240 116.900 ;
    RECT 79.520 2.100 80.920 116.900 ;
    RECT 81.200 2.100 82.600 116.900 ;
    RECT 82.880 2.100 84.280 116.900 ;
    RECT 84.560 2.100 85.960 116.900 ;
    RECT 86.240 2.100 87.640 116.900 ;
    RECT 87.920 2.100 89.320 116.900 ;
    RECT 89.600 2.100 91.000 116.900 ;
    RECT 91.280 2.100 92.680 116.900 ;
    RECT 92.960 2.100 94.360 116.900 ;
    RECT 94.640 2.100 96.040 116.900 ;
    RECT 96.320 2.100 97.720 116.900 ;
    RECT 98.000 2.100 99.400 116.900 ;
    RECT 99.680 2.100 101.080 116.900 ;
    RECT 101.360 2.100 102.760 116.900 ;
    RECT 103.040 2.100 104.440 116.900 ;
    RECT 104.720 2.100 106.120 116.900 ;
    RECT 106.400 2.100 107.800 116.900 ;
    RECT 108.080 2.100 109.480 116.900 ;
    RECT 109.760 2.100 111.160 116.900 ;
    RECT 111.440 2.100 112.840 116.900 ;
    RECT 113.120 2.100 115.140 116.900 ;
    LAYER OVERLAP ;
    RECT 0 0 115.140 119.000 ;
  END
END fakeram45_256x96

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_256x95
  FOREIGN fakeram45_256x95 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 115.140 BY 119.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.275 0.070 2.345 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.695 0.070 2.765 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.115 0.070 3.185 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.535 0.070 3.605 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.955 0.070 4.025 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.375 0.070 4.445 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.795 0.070 4.865 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.215 0.070 5.285 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.635 0.070 5.705 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.055 0.070 6.125 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.475 0.070 6.545 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.895 0.070 6.965 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.315 0.070 7.385 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.735 0.070 7.805 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.155 0.070 8.225 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.575 0.070 8.645 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.785 0.070 8.855 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.995 0.070 9.065 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.415 0.070 9.485 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.835 0.070 9.905 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.255 0.070 10.325 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.675 0.070 10.745 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.095 0.070 11.165 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.515 0.070 11.585 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.935 0.070 12.005 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.355 0.070 12.425 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.775 0.070 12.845 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.985 0.070 13.055 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.195 0.070 13.265 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.615 0.070 13.685 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.035 0.070 14.105 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.455 0.070 14.525 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.875 0.070 14.945 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.295 0.070 15.365 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.505 0.070 15.575 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.715 0.070 15.785 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.135 0.070 16.205 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.345 0.070 16.415 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.555 0.070 16.625 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.975 0.070 17.045 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.185 0.070 17.255 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.395 0.070 17.465 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.605 0.070 17.675 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.815 0.070 17.885 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.025 0.070 18.095 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.235 0.070 18.305 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.655 0.070 18.725 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.075 0.070 19.145 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.495 0.070 19.565 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.915 0.070 19.985 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.335 0.070 20.405 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.545 0.070 20.615 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.755 0.070 20.825 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.175 0.070 21.245 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.595 0.070 21.665 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END w_mask_in[94]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.825 0.070 34.895 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.035 0.070 35.105 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.455 0.070 35.525 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.875 0.070 35.945 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.295 0.070 36.365 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.505 0.070 36.575 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.715 0.070 36.785 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.135 0.070 37.205 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.555 0.070 37.625 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.975 0.070 38.045 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.185 0.070 38.255 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.395 0.070 38.465 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.815 0.070 38.885 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.235 0.070 39.305 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.655 0.070 39.725 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.075 0.070 40.145 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.495 0.070 40.565 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.915 0.070 40.985 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.335 0.070 41.405 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.755 0.070 41.825 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.175 0.070 42.245 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.595 0.070 42.665 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.015 0.070 43.085 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.435 0.070 43.505 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.855 0.070 43.925 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.275 0.070 44.345 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.695 0.070 44.765 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.115 0.070 45.185 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.325 0.070 45.395 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.535 0.070 45.605 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.745 0.070 45.815 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.955 0.070 46.025 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.375 0.070 46.445 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.585 0.070 46.655 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.795 0.070 46.865 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.215 0.070 47.285 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.635 0.070 47.705 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.055 0.070 48.125 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.265 0.070 48.335 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.475 0.070 48.545 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.895 0.070 48.965 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.315 0.070 49.385 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.735 0.070 49.805 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.945 0.070 50.015 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.155 0.070 50.225 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.575 0.070 50.645 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.785 0.070 50.855 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.995 0.070 51.065 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.205 0.070 51.275 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.415 0.070 51.485 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.625 0.070 51.695 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.835 0.070 51.905 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.045 0.070 52.115 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.255 0.070 52.325 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.675 0.070 52.745 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.095 0.070 53.165 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.305 0.070 53.375 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.515 0.070 53.585 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.935 0.070 54.005 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.145 0.070 54.215 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.355 0.070 54.425 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END rd_out[94]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.585 0.070 67.655 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.795 0.070 67.865 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.215 0.070 68.285 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.425 0.070 68.495 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.635 0.070 68.705 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.845 0.070 68.915 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.055 0.070 69.125 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.265 0.070 69.335 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.475 0.070 69.545 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.685 0.070 69.755 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.895 0.070 69.965 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.105 0.070 70.175 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.315 0.070 70.385 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.735 0.070 70.805 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.945 0.070 71.015 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.155 0.070 71.225 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.575 0.070 71.645 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.785 0.070 71.855 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.995 0.070 72.065 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.205 0.070 72.275 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.415 0.070 72.485 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.625 0.070 72.695 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.835 0.070 72.905 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.255 0.070 73.325 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.465 0.070 73.535 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.675 0.070 73.745 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.095 0.070 74.165 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.305 0.070 74.375 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.515 0.070 74.585 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.725 0.070 74.795 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.935 0.070 75.005 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.145 0.070 75.215 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.355 0.070 75.425 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.775 0.070 75.845 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.195 0.070 76.265 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.405 0.070 76.475 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.615 0.070 76.685 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.825 0.070 76.895 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.035 0.070 77.105 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.245 0.070 77.315 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.455 0.070 77.525 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.665 0.070 77.735 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.875 0.070 77.945 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.085 0.070 78.155 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.295 0.070 78.365 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.505 0.070 78.575 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.715 0.070 78.785 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.925 0.070 78.995 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.135 0.070 79.205 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.345 0.070 79.415 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.555 0.070 79.625 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.975 0.070 80.045 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.185 0.070 80.255 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.395 0.070 80.465 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.605 0.070 80.675 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.815 0.070 80.885 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.025 0.070 81.095 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.235 0.070 81.305 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.445 0.070 81.515 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.655 0.070 81.725 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.075 0.070 82.145 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.285 0.070 82.355 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.495 0.070 82.565 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.705 0.070 82.775 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.915 0.070 82.985 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.125 0.070 83.195 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.335 0.070 83.405 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.545 0.070 83.615 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.755 0.070 83.825 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.965 0.070 84.035 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.175 0.070 84.245 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.385 0.070 84.455 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.595 0.070 84.665 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.015 0.070 85.085 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.225 0.070 85.295 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.435 0.070 85.505 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.855 0.070 85.925 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.065 0.070 86.135 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.275 0.070 86.345 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.485 0.070 86.555 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.695 0.070 86.765 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.905 0.070 86.975 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.115 0.070 87.185 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.325 0.070 87.395 ;
    END
  END wd_in[94]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.345 0.070 100.415 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.555 0.070 100.625 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.765 0.070 100.835 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.975 0.070 101.045 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.185 0.070 101.255 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.395 0.070 101.465 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.605 0.070 101.675 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.815 0.070 101.885 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.835 0.070 114.905 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.045 0.070 115.115 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.255 0.070 115.325 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 116.900 ;
      RECT 5.320 2.100 5.600 116.900 ;
      RECT 8.680 2.100 8.960 116.900 ;
      RECT 12.040 2.100 12.320 116.900 ;
      RECT 15.400 2.100 15.680 116.900 ;
      RECT 18.760 2.100 19.040 116.900 ;
      RECT 22.120 2.100 22.400 116.900 ;
      RECT 25.480 2.100 25.760 116.900 ;
      RECT 28.840 2.100 29.120 116.900 ;
      RECT 32.200 2.100 32.480 116.900 ;
      RECT 35.560 2.100 35.840 116.900 ;
      RECT 38.920 2.100 39.200 116.900 ;
      RECT 42.280 2.100 42.560 116.900 ;
      RECT 45.640 2.100 45.920 116.900 ;
      RECT 49.000 2.100 49.280 116.900 ;
      RECT 52.360 2.100 52.640 116.900 ;
      RECT 55.720 2.100 56.000 116.900 ;
      RECT 59.080 2.100 59.360 116.900 ;
      RECT 62.440 2.100 62.720 116.900 ;
      RECT 65.800 2.100 66.080 116.900 ;
      RECT 69.160 2.100 69.440 116.900 ;
      RECT 72.520 2.100 72.800 116.900 ;
      RECT 75.880 2.100 76.160 116.900 ;
      RECT 79.240 2.100 79.520 116.900 ;
      RECT 82.600 2.100 82.880 116.900 ;
      RECT 85.960 2.100 86.240 116.900 ;
      RECT 89.320 2.100 89.600 116.900 ;
      RECT 92.680 2.100 92.960 116.900 ;
      RECT 96.040 2.100 96.320 116.900 ;
      RECT 99.400 2.100 99.680 116.900 ;
      RECT 102.760 2.100 103.040 116.900 ;
      RECT 106.120 2.100 106.400 116.900 ;
      RECT 109.480 2.100 109.760 116.900 ;
      RECT 112.840 2.100 113.120 116.900 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 116.900 ;
      RECT 7.000 2.100 7.280 116.900 ;
      RECT 10.360 2.100 10.640 116.900 ;
      RECT 13.720 2.100 14.000 116.900 ;
      RECT 17.080 2.100 17.360 116.900 ;
      RECT 20.440 2.100 20.720 116.900 ;
      RECT 23.800 2.100 24.080 116.900 ;
      RECT 27.160 2.100 27.440 116.900 ;
      RECT 30.520 2.100 30.800 116.900 ;
      RECT 33.880 2.100 34.160 116.900 ;
      RECT 37.240 2.100 37.520 116.900 ;
      RECT 40.600 2.100 40.880 116.900 ;
      RECT 43.960 2.100 44.240 116.900 ;
      RECT 47.320 2.100 47.600 116.900 ;
      RECT 50.680 2.100 50.960 116.900 ;
      RECT 54.040 2.100 54.320 116.900 ;
      RECT 57.400 2.100 57.680 116.900 ;
      RECT 60.760 2.100 61.040 116.900 ;
      RECT 64.120 2.100 64.400 116.900 ;
      RECT 67.480 2.100 67.760 116.900 ;
      RECT 70.840 2.100 71.120 116.900 ;
      RECT 74.200 2.100 74.480 116.900 ;
      RECT 77.560 2.100 77.840 116.900 ;
      RECT 80.920 2.100 81.200 116.900 ;
      RECT 84.280 2.100 84.560 116.900 ;
      RECT 87.640 2.100 87.920 116.900 ;
      RECT 91.000 2.100 91.280 116.900 ;
      RECT 94.360 2.100 94.640 116.900 ;
      RECT 97.720 2.100 98.000 116.900 ;
      RECT 101.080 2.100 101.360 116.900 ;
      RECT 104.440 2.100 104.720 116.900 ;
      RECT 107.800 2.100 108.080 116.900 ;
      RECT 111.160 2.100 111.440 116.900 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 115.140 119.000 ;
    LAYER metal2 ;
    RECT 0 0 115.140 119.000 ;
    LAYER metal3 ;
    RECT 0.070 0 115.140 119.000 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.275 ;
    RECT 0 2.345 0.070 2.485 ;
    RECT 0 2.555 0.070 2.695 ;
    RECT 0 2.765 0.070 2.905 ;
    RECT 0 2.975 0.070 3.115 ;
    RECT 0 3.185 0.070 3.325 ;
    RECT 0 3.395 0.070 3.535 ;
    RECT 0 3.605 0.070 3.745 ;
    RECT 0 3.815 0.070 3.955 ;
    RECT 0 4.025 0.070 4.165 ;
    RECT 0 4.235 0.070 4.375 ;
    RECT 0 4.445 0.070 4.585 ;
    RECT 0 4.655 0.070 4.795 ;
    RECT 0 4.865 0.070 5.005 ;
    RECT 0 5.075 0.070 5.215 ;
    RECT 0 5.285 0.070 5.425 ;
    RECT 0 5.495 0.070 5.635 ;
    RECT 0 5.705 0.070 5.845 ;
    RECT 0 5.915 0.070 6.055 ;
    RECT 0 6.125 0.070 6.265 ;
    RECT 0 6.335 0.070 6.475 ;
    RECT 0 6.545 0.070 6.685 ;
    RECT 0 6.755 0.070 6.895 ;
    RECT 0 6.965 0.070 7.105 ;
    RECT 0 7.175 0.070 7.315 ;
    RECT 0 7.385 0.070 7.525 ;
    RECT 0 7.595 0.070 7.735 ;
    RECT 0 7.805 0.070 7.945 ;
    RECT 0 8.015 0.070 8.155 ;
    RECT 0 8.225 0.070 8.365 ;
    RECT 0 8.435 0.070 8.575 ;
    RECT 0 8.645 0.070 8.785 ;
    RECT 0 8.855 0.070 8.995 ;
    RECT 0 9.065 0.070 9.205 ;
    RECT 0 9.275 0.070 9.415 ;
    RECT 0 9.485 0.070 9.625 ;
    RECT 0 9.695 0.070 9.835 ;
    RECT 0 9.905 0.070 10.045 ;
    RECT 0 10.115 0.070 10.255 ;
    RECT 0 10.325 0.070 10.465 ;
    RECT 0 10.535 0.070 10.675 ;
    RECT 0 10.745 0.070 10.885 ;
    RECT 0 10.955 0.070 11.095 ;
    RECT 0 11.165 0.070 11.305 ;
    RECT 0 11.375 0.070 11.515 ;
    RECT 0 11.585 0.070 11.725 ;
    RECT 0 11.795 0.070 11.935 ;
    RECT 0 12.005 0.070 12.145 ;
    RECT 0 12.215 0.070 12.355 ;
    RECT 0 12.425 0.070 12.565 ;
    RECT 0 12.635 0.070 12.775 ;
    RECT 0 12.845 0.070 12.985 ;
    RECT 0 13.055 0.070 13.195 ;
    RECT 0 13.265 0.070 13.405 ;
    RECT 0 13.475 0.070 13.615 ;
    RECT 0 13.685 0.070 13.825 ;
    RECT 0 13.895 0.070 14.035 ;
    RECT 0 14.105 0.070 14.245 ;
    RECT 0 14.315 0.070 14.455 ;
    RECT 0 14.525 0.070 14.665 ;
    RECT 0 14.735 0.070 14.875 ;
    RECT 0 14.945 0.070 15.085 ;
    RECT 0 15.155 0.070 15.295 ;
    RECT 0 15.365 0.070 15.505 ;
    RECT 0 15.575 0.070 15.715 ;
    RECT 0 15.785 0.070 15.925 ;
    RECT 0 15.995 0.070 16.135 ;
    RECT 0 16.205 0.070 16.345 ;
    RECT 0 16.415 0.070 16.555 ;
    RECT 0 16.625 0.070 16.765 ;
    RECT 0 16.835 0.070 16.975 ;
    RECT 0 17.045 0.070 17.185 ;
    RECT 0 17.255 0.070 17.395 ;
    RECT 0 17.465 0.070 17.605 ;
    RECT 0 17.675 0.070 17.815 ;
    RECT 0 17.885 0.070 18.025 ;
    RECT 0 18.095 0.070 18.235 ;
    RECT 0 18.305 0.070 18.445 ;
    RECT 0 18.515 0.070 18.655 ;
    RECT 0 18.725 0.070 18.865 ;
    RECT 0 18.935 0.070 19.075 ;
    RECT 0 19.145 0.070 19.285 ;
    RECT 0 19.355 0.070 19.495 ;
    RECT 0 19.565 0.070 19.705 ;
    RECT 0 19.775 0.070 19.915 ;
    RECT 0 19.985 0.070 20.125 ;
    RECT 0 20.195 0.070 20.335 ;
    RECT 0 20.405 0.070 20.545 ;
    RECT 0 20.615 0.070 20.755 ;
    RECT 0 20.825 0.070 20.965 ;
    RECT 0 21.035 0.070 21.175 ;
    RECT 0 21.245 0.070 21.385 ;
    RECT 0 21.455 0.070 21.595 ;
    RECT 0 21.665 0.070 21.805 ;
    RECT 0 21.875 0.070 34.825 ;
    RECT 0 34.895 0.070 35.035 ;
    RECT 0 35.105 0.070 35.245 ;
    RECT 0 35.315 0.070 35.455 ;
    RECT 0 35.525 0.070 35.665 ;
    RECT 0 35.735 0.070 35.875 ;
    RECT 0 35.945 0.070 36.085 ;
    RECT 0 36.155 0.070 36.295 ;
    RECT 0 36.365 0.070 36.505 ;
    RECT 0 36.575 0.070 36.715 ;
    RECT 0 36.785 0.070 36.925 ;
    RECT 0 36.995 0.070 37.135 ;
    RECT 0 37.205 0.070 37.345 ;
    RECT 0 37.415 0.070 37.555 ;
    RECT 0 37.625 0.070 37.765 ;
    RECT 0 37.835 0.070 37.975 ;
    RECT 0 38.045 0.070 38.185 ;
    RECT 0 38.255 0.070 38.395 ;
    RECT 0 38.465 0.070 38.605 ;
    RECT 0 38.675 0.070 38.815 ;
    RECT 0 38.885 0.070 39.025 ;
    RECT 0 39.095 0.070 39.235 ;
    RECT 0 39.305 0.070 39.445 ;
    RECT 0 39.515 0.070 39.655 ;
    RECT 0 39.725 0.070 39.865 ;
    RECT 0 39.935 0.070 40.075 ;
    RECT 0 40.145 0.070 40.285 ;
    RECT 0 40.355 0.070 40.495 ;
    RECT 0 40.565 0.070 40.705 ;
    RECT 0 40.775 0.070 40.915 ;
    RECT 0 40.985 0.070 41.125 ;
    RECT 0 41.195 0.070 41.335 ;
    RECT 0 41.405 0.070 41.545 ;
    RECT 0 41.615 0.070 41.755 ;
    RECT 0 41.825 0.070 41.965 ;
    RECT 0 42.035 0.070 42.175 ;
    RECT 0 42.245 0.070 42.385 ;
    RECT 0 42.455 0.070 42.595 ;
    RECT 0 42.665 0.070 42.805 ;
    RECT 0 42.875 0.070 43.015 ;
    RECT 0 43.085 0.070 43.225 ;
    RECT 0 43.295 0.070 43.435 ;
    RECT 0 43.505 0.070 43.645 ;
    RECT 0 43.715 0.070 43.855 ;
    RECT 0 43.925 0.070 44.065 ;
    RECT 0 44.135 0.070 44.275 ;
    RECT 0 44.345 0.070 44.485 ;
    RECT 0 44.555 0.070 44.695 ;
    RECT 0 44.765 0.070 44.905 ;
    RECT 0 44.975 0.070 45.115 ;
    RECT 0 45.185 0.070 45.325 ;
    RECT 0 45.395 0.070 45.535 ;
    RECT 0 45.605 0.070 45.745 ;
    RECT 0 45.815 0.070 45.955 ;
    RECT 0 46.025 0.070 46.165 ;
    RECT 0 46.235 0.070 46.375 ;
    RECT 0 46.445 0.070 46.585 ;
    RECT 0 46.655 0.070 46.795 ;
    RECT 0 46.865 0.070 47.005 ;
    RECT 0 47.075 0.070 47.215 ;
    RECT 0 47.285 0.070 47.425 ;
    RECT 0 47.495 0.070 47.635 ;
    RECT 0 47.705 0.070 47.845 ;
    RECT 0 47.915 0.070 48.055 ;
    RECT 0 48.125 0.070 48.265 ;
    RECT 0 48.335 0.070 48.475 ;
    RECT 0 48.545 0.070 48.685 ;
    RECT 0 48.755 0.070 48.895 ;
    RECT 0 48.965 0.070 49.105 ;
    RECT 0 49.175 0.070 49.315 ;
    RECT 0 49.385 0.070 49.525 ;
    RECT 0 49.595 0.070 49.735 ;
    RECT 0 49.805 0.070 49.945 ;
    RECT 0 50.015 0.070 50.155 ;
    RECT 0 50.225 0.070 50.365 ;
    RECT 0 50.435 0.070 50.575 ;
    RECT 0 50.645 0.070 50.785 ;
    RECT 0 50.855 0.070 50.995 ;
    RECT 0 51.065 0.070 51.205 ;
    RECT 0 51.275 0.070 51.415 ;
    RECT 0 51.485 0.070 51.625 ;
    RECT 0 51.695 0.070 51.835 ;
    RECT 0 51.905 0.070 52.045 ;
    RECT 0 52.115 0.070 52.255 ;
    RECT 0 52.325 0.070 52.465 ;
    RECT 0 52.535 0.070 52.675 ;
    RECT 0 52.745 0.070 52.885 ;
    RECT 0 52.955 0.070 53.095 ;
    RECT 0 53.165 0.070 53.305 ;
    RECT 0 53.375 0.070 53.515 ;
    RECT 0 53.585 0.070 53.725 ;
    RECT 0 53.795 0.070 53.935 ;
    RECT 0 54.005 0.070 54.145 ;
    RECT 0 54.215 0.070 54.355 ;
    RECT 0 54.425 0.070 54.565 ;
    RECT 0 54.635 0.070 67.585 ;
    RECT 0 67.655 0.070 67.795 ;
    RECT 0 67.865 0.070 68.005 ;
    RECT 0 68.075 0.070 68.215 ;
    RECT 0 68.285 0.070 68.425 ;
    RECT 0 68.495 0.070 68.635 ;
    RECT 0 68.705 0.070 68.845 ;
    RECT 0 68.915 0.070 69.055 ;
    RECT 0 69.125 0.070 69.265 ;
    RECT 0 69.335 0.070 69.475 ;
    RECT 0 69.545 0.070 69.685 ;
    RECT 0 69.755 0.070 69.895 ;
    RECT 0 69.965 0.070 70.105 ;
    RECT 0 70.175 0.070 70.315 ;
    RECT 0 70.385 0.070 70.525 ;
    RECT 0 70.595 0.070 70.735 ;
    RECT 0 70.805 0.070 70.945 ;
    RECT 0 71.015 0.070 71.155 ;
    RECT 0 71.225 0.070 71.365 ;
    RECT 0 71.435 0.070 71.575 ;
    RECT 0 71.645 0.070 71.785 ;
    RECT 0 71.855 0.070 71.995 ;
    RECT 0 72.065 0.070 72.205 ;
    RECT 0 72.275 0.070 72.415 ;
    RECT 0 72.485 0.070 72.625 ;
    RECT 0 72.695 0.070 72.835 ;
    RECT 0 72.905 0.070 73.045 ;
    RECT 0 73.115 0.070 73.255 ;
    RECT 0 73.325 0.070 73.465 ;
    RECT 0 73.535 0.070 73.675 ;
    RECT 0 73.745 0.070 73.885 ;
    RECT 0 73.955 0.070 74.095 ;
    RECT 0 74.165 0.070 74.305 ;
    RECT 0 74.375 0.070 74.515 ;
    RECT 0 74.585 0.070 74.725 ;
    RECT 0 74.795 0.070 74.935 ;
    RECT 0 75.005 0.070 75.145 ;
    RECT 0 75.215 0.070 75.355 ;
    RECT 0 75.425 0.070 75.565 ;
    RECT 0 75.635 0.070 75.775 ;
    RECT 0 75.845 0.070 75.985 ;
    RECT 0 76.055 0.070 76.195 ;
    RECT 0 76.265 0.070 76.405 ;
    RECT 0 76.475 0.070 76.615 ;
    RECT 0 76.685 0.070 76.825 ;
    RECT 0 76.895 0.070 77.035 ;
    RECT 0 77.105 0.070 77.245 ;
    RECT 0 77.315 0.070 77.455 ;
    RECT 0 77.525 0.070 77.665 ;
    RECT 0 77.735 0.070 77.875 ;
    RECT 0 77.945 0.070 78.085 ;
    RECT 0 78.155 0.070 78.295 ;
    RECT 0 78.365 0.070 78.505 ;
    RECT 0 78.575 0.070 78.715 ;
    RECT 0 78.785 0.070 78.925 ;
    RECT 0 78.995 0.070 79.135 ;
    RECT 0 79.205 0.070 79.345 ;
    RECT 0 79.415 0.070 79.555 ;
    RECT 0 79.625 0.070 79.765 ;
    RECT 0 79.835 0.070 79.975 ;
    RECT 0 80.045 0.070 80.185 ;
    RECT 0 80.255 0.070 80.395 ;
    RECT 0 80.465 0.070 80.605 ;
    RECT 0 80.675 0.070 80.815 ;
    RECT 0 80.885 0.070 81.025 ;
    RECT 0 81.095 0.070 81.235 ;
    RECT 0 81.305 0.070 81.445 ;
    RECT 0 81.515 0.070 81.655 ;
    RECT 0 81.725 0.070 81.865 ;
    RECT 0 81.935 0.070 82.075 ;
    RECT 0 82.145 0.070 82.285 ;
    RECT 0 82.355 0.070 82.495 ;
    RECT 0 82.565 0.070 82.705 ;
    RECT 0 82.775 0.070 82.915 ;
    RECT 0 82.985 0.070 83.125 ;
    RECT 0 83.195 0.070 83.335 ;
    RECT 0 83.405 0.070 83.545 ;
    RECT 0 83.615 0.070 83.755 ;
    RECT 0 83.825 0.070 83.965 ;
    RECT 0 84.035 0.070 84.175 ;
    RECT 0 84.245 0.070 84.385 ;
    RECT 0 84.455 0.070 84.595 ;
    RECT 0 84.665 0.070 84.805 ;
    RECT 0 84.875 0.070 85.015 ;
    RECT 0 85.085 0.070 85.225 ;
    RECT 0 85.295 0.070 85.435 ;
    RECT 0 85.505 0.070 85.645 ;
    RECT 0 85.715 0.070 85.855 ;
    RECT 0 85.925 0.070 86.065 ;
    RECT 0 86.135 0.070 86.275 ;
    RECT 0 86.345 0.070 86.485 ;
    RECT 0 86.555 0.070 86.695 ;
    RECT 0 86.765 0.070 86.905 ;
    RECT 0 86.975 0.070 87.115 ;
    RECT 0 87.185 0.070 87.325 ;
    RECT 0 87.395 0.070 100.345 ;
    RECT 0 100.415 0.070 100.555 ;
    RECT 0 100.625 0.070 100.765 ;
    RECT 0 100.835 0.070 100.975 ;
    RECT 0 101.045 0.070 101.185 ;
    RECT 0 101.255 0.070 101.395 ;
    RECT 0 101.465 0.070 101.605 ;
    RECT 0 101.675 0.070 101.815 ;
    RECT 0 101.885 0.070 114.835 ;
    RECT 0 114.905 0.070 115.045 ;
    RECT 0 115.115 0.070 115.255 ;
    RECT 0 115.325 0.070 119.000 ;
    LAYER metal4 ;
    RECT 0 0 115.140 2.100 ;
    RECT 0 116.900 115.140 119.000 ;
    RECT 0.000 2.100 1.960 116.900 ;
    RECT 2.240 2.100 3.640 116.900 ;
    RECT 3.920 2.100 5.320 116.900 ;
    RECT 5.600 2.100 7.000 116.900 ;
    RECT 7.280 2.100 8.680 116.900 ;
    RECT 8.960 2.100 10.360 116.900 ;
    RECT 10.640 2.100 12.040 116.900 ;
    RECT 12.320 2.100 13.720 116.900 ;
    RECT 14.000 2.100 15.400 116.900 ;
    RECT 15.680 2.100 17.080 116.900 ;
    RECT 17.360 2.100 18.760 116.900 ;
    RECT 19.040 2.100 20.440 116.900 ;
    RECT 20.720 2.100 22.120 116.900 ;
    RECT 22.400 2.100 23.800 116.900 ;
    RECT 24.080 2.100 25.480 116.900 ;
    RECT 25.760 2.100 27.160 116.900 ;
    RECT 27.440 2.100 28.840 116.900 ;
    RECT 29.120 2.100 30.520 116.900 ;
    RECT 30.800 2.100 32.200 116.900 ;
    RECT 32.480 2.100 33.880 116.900 ;
    RECT 34.160 2.100 35.560 116.900 ;
    RECT 35.840 2.100 37.240 116.900 ;
    RECT 37.520 2.100 38.920 116.900 ;
    RECT 39.200 2.100 40.600 116.900 ;
    RECT 40.880 2.100 42.280 116.900 ;
    RECT 42.560 2.100 43.960 116.900 ;
    RECT 44.240 2.100 45.640 116.900 ;
    RECT 45.920 2.100 47.320 116.900 ;
    RECT 47.600 2.100 49.000 116.900 ;
    RECT 49.280 2.100 50.680 116.900 ;
    RECT 50.960 2.100 52.360 116.900 ;
    RECT 52.640 2.100 54.040 116.900 ;
    RECT 54.320 2.100 55.720 116.900 ;
    RECT 56.000 2.100 57.400 116.900 ;
    RECT 57.680 2.100 59.080 116.900 ;
    RECT 59.360 2.100 60.760 116.900 ;
    RECT 61.040 2.100 62.440 116.900 ;
    RECT 62.720 2.100 64.120 116.900 ;
    RECT 64.400 2.100 65.800 116.900 ;
    RECT 66.080 2.100 67.480 116.900 ;
    RECT 67.760 2.100 69.160 116.900 ;
    RECT 69.440 2.100 70.840 116.900 ;
    RECT 71.120 2.100 72.520 116.900 ;
    RECT 72.800 2.100 74.200 116.900 ;
    RECT 74.480 2.100 75.880 116.900 ;
    RECT 76.160 2.100 77.560 116.900 ;
    RECT 77.840 2.100 79.240 116.900 ;
    RECT 79.520 2.100 80.920 116.900 ;
    RECT 81.200 2.100 82.600 116.900 ;
    RECT 82.880 2.100 84.280 116.900 ;
    RECT 84.560 2.100 85.960 116.900 ;
    RECT 86.240 2.100 87.640 116.900 ;
    RECT 87.920 2.100 89.320 116.900 ;
    RECT 89.600 2.100 91.000 116.900 ;
    RECT 91.280 2.100 92.680 116.900 ;
    RECT 92.960 2.100 94.360 116.900 ;
    RECT 94.640 2.100 96.040 116.900 ;
    RECT 96.320 2.100 97.720 116.900 ;
    RECT 98.000 2.100 99.400 116.900 ;
    RECT 99.680 2.100 101.080 116.900 ;
    RECT 101.360 2.100 102.760 116.900 ;
    RECT 103.040 2.100 104.440 116.900 ;
    RECT 104.720 2.100 106.120 116.900 ;
    RECT 106.400 2.100 107.800 116.900 ;
    RECT 108.080 2.100 109.480 116.900 ;
    RECT 109.760 2.100 111.160 116.900 ;
    RECT 111.440 2.100 112.840 116.900 ;
    RECT 113.120 2.100 115.140 116.900 ;
    LAYER OVERLAP ;
    RECT 0 0 115.140 119.000 ;
  END
END fakeram45_256x95

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_256x48
  FOREIGN fakeram45_256x48 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 64.030 BY 207.200 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.185 0.070 17.255 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.225 0.070 22.295 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.785 0.070 29.855 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.045 0.070 31.115 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.305 0.070 32.375 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.825 0.070 34.895 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.945 0.070 50.015 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.205 0.070 51.275 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.985 0.070 55.055 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.505 0.070 57.575 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.765 0.070 58.835 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.025 0.070 60.095 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.285 0.070 61.355 ;
    END
  END w_mask_in[47]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.175 0.070 63.245 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.435 0.070 64.505 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.695 0.070 65.765 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.955 0.070 67.025 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.215 0.070 68.285 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.475 0.070 69.545 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.735 0.070 70.805 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.995 0.070 72.065 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.255 0.070 73.325 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.515 0.070 74.585 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.775 0.070 75.845 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.035 0.070 77.105 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.295 0.070 78.365 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.555 0.070 79.625 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.815 0.070 80.885 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.075 0.070 82.145 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.335 0.070 83.405 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.595 0.070 84.665 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.855 0.070 85.925 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.115 0.070 87.185 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.375 0.070 88.445 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.635 0.070 89.705 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.895 0.070 90.965 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.155 0.070 92.225 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.415 0.070 93.485 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.675 0.070 94.745 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.935 0.070 96.005 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.195 0.070 97.265 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.455 0.070 98.525 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.715 0.070 99.785 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.975 0.070 101.045 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.235 0.070 102.305 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.495 0.070 103.565 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.755 0.070 104.825 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.015 0.070 106.085 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.275 0.070 107.345 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.535 0.070 108.605 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.795 0.070 109.865 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.055 0.070 111.125 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.315 0.070 112.385 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.575 0.070 113.645 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.835 0.070 114.905 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.095 0.070 116.165 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.355 0.070 117.425 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.615 0.070 118.685 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.875 0.070 119.945 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.135 0.070 121.205 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.395 0.070 122.465 ;
    END
  END rd_out[47]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.285 0.070 124.355 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.545 0.070 125.615 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.805 0.070 126.875 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 128.065 0.070 128.135 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.325 0.070 129.395 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.585 0.070 130.655 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 131.845 0.070 131.915 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.105 0.070 133.175 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 134.365 0.070 134.435 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.625 0.070 135.695 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.885 0.070 136.955 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.145 0.070 138.215 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.405 0.070 139.475 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 140.665 0.070 140.735 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.925 0.070 141.995 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 143.185 0.070 143.255 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.445 0.070 144.515 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.705 0.070 145.775 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.965 0.070 147.035 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.225 0.070 148.295 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.485 0.070 149.555 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.745 0.070 150.815 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.005 0.070 152.075 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.265 0.070 153.335 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.525 0.070 154.595 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.785 0.070 155.855 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.045 0.070 157.115 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.305 0.070 158.375 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.565 0.070 159.635 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.825 0.070 160.895 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.085 0.070 162.155 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.345 0.070 163.415 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.605 0.070 164.675 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.865 0.070 165.935 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.125 0.070 167.195 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.385 0.070 168.455 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.645 0.070 169.715 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.905 0.070 170.975 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.165 0.070 172.235 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.425 0.070 173.495 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.685 0.070 174.755 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.945 0.070 176.015 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.205 0.070 177.275 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.465 0.070 178.535 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.725 0.070 179.795 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.985 0.070 181.055 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.245 0.070 182.315 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.505 0.070 183.575 ;
    END
  END wd_in[47]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.395 0.070 185.465 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.655 0.070 186.725 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.915 0.070 187.985 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.175 0.070 189.245 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.435 0.070 190.505 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.695 0.070 191.765 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.955 0.070 193.025 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.215 0.070 194.285 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.105 0.070 196.175 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.365 0.070 197.435 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 198.625 0.070 198.695 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 205.100 ;
      RECT 5.320 2.100 5.600 205.100 ;
      RECT 8.680 2.100 8.960 205.100 ;
      RECT 12.040 2.100 12.320 205.100 ;
      RECT 15.400 2.100 15.680 205.100 ;
      RECT 18.760 2.100 19.040 205.100 ;
      RECT 22.120 2.100 22.400 205.100 ;
      RECT 25.480 2.100 25.760 205.100 ;
      RECT 28.840 2.100 29.120 205.100 ;
      RECT 32.200 2.100 32.480 205.100 ;
      RECT 35.560 2.100 35.840 205.100 ;
      RECT 38.920 2.100 39.200 205.100 ;
      RECT 42.280 2.100 42.560 205.100 ;
      RECT 45.640 2.100 45.920 205.100 ;
      RECT 49.000 2.100 49.280 205.100 ;
      RECT 52.360 2.100 52.640 205.100 ;
      RECT 55.720 2.100 56.000 205.100 ;
      RECT 59.080 2.100 59.360 205.100 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 205.100 ;
      RECT 7.000 2.100 7.280 205.100 ;
      RECT 10.360 2.100 10.640 205.100 ;
      RECT 13.720 2.100 14.000 205.100 ;
      RECT 17.080 2.100 17.360 205.100 ;
      RECT 20.440 2.100 20.720 205.100 ;
      RECT 23.800 2.100 24.080 205.100 ;
      RECT 27.160 2.100 27.440 205.100 ;
      RECT 30.520 2.100 30.800 205.100 ;
      RECT 33.880 2.100 34.160 205.100 ;
      RECT 37.240 2.100 37.520 205.100 ;
      RECT 40.600 2.100 40.880 205.100 ;
      RECT 43.960 2.100 44.240 205.100 ;
      RECT 47.320 2.100 47.600 205.100 ;
      RECT 50.680 2.100 50.960 205.100 ;
      RECT 54.040 2.100 54.320 205.100 ;
      RECT 57.400 2.100 57.680 205.100 ;
      RECT 60.760 2.100 61.040 205.100 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 64.030 207.200 ;
    LAYER metal2 ;
    RECT 0 0 64.030 207.200 ;
    LAYER metal3 ;
    RECT 0.070 0 64.030 207.200 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 3.325 ;
    RECT 0 3.395 0.070 4.585 ;
    RECT 0 4.655 0.070 5.845 ;
    RECT 0 5.915 0.070 7.105 ;
    RECT 0 7.175 0.070 8.365 ;
    RECT 0 8.435 0.070 9.625 ;
    RECT 0 9.695 0.070 10.885 ;
    RECT 0 10.955 0.070 12.145 ;
    RECT 0 12.215 0.070 13.405 ;
    RECT 0 13.475 0.070 14.665 ;
    RECT 0 14.735 0.070 15.925 ;
    RECT 0 15.995 0.070 17.185 ;
    RECT 0 17.255 0.070 18.445 ;
    RECT 0 18.515 0.070 19.705 ;
    RECT 0 19.775 0.070 20.965 ;
    RECT 0 21.035 0.070 22.225 ;
    RECT 0 22.295 0.070 23.485 ;
    RECT 0 23.555 0.070 24.745 ;
    RECT 0 24.815 0.070 26.005 ;
    RECT 0 26.075 0.070 27.265 ;
    RECT 0 27.335 0.070 28.525 ;
    RECT 0 28.595 0.070 29.785 ;
    RECT 0 29.855 0.070 31.045 ;
    RECT 0 31.115 0.070 32.305 ;
    RECT 0 32.375 0.070 33.565 ;
    RECT 0 33.635 0.070 34.825 ;
    RECT 0 34.895 0.070 36.085 ;
    RECT 0 36.155 0.070 37.345 ;
    RECT 0 37.415 0.070 38.605 ;
    RECT 0 38.675 0.070 39.865 ;
    RECT 0 39.935 0.070 41.125 ;
    RECT 0 41.195 0.070 42.385 ;
    RECT 0 42.455 0.070 43.645 ;
    RECT 0 43.715 0.070 44.905 ;
    RECT 0 44.975 0.070 46.165 ;
    RECT 0 46.235 0.070 47.425 ;
    RECT 0 47.495 0.070 48.685 ;
    RECT 0 48.755 0.070 49.945 ;
    RECT 0 50.015 0.070 51.205 ;
    RECT 0 51.275 0.070 52.465 ;
    RECT 0 52.535 0.070 53.725 ;
    RECT 0 53.795 0.070 54.985 ;
    RECT 0 55.055 0.070 56.245 ;
    RECT 0 56.315 0.070 57.505 ;
    RECT 0 57.575 0.070 58.765 ;
    RECT 0 58.835 0.070 60.025 ;
    RECT 0 60.095 0.070 61.285 ;
    RECT 0 61.355 0.070 63.175 ;
    RECT 0 63.245 0.070 64.435 ;
    RECT 0 64.505 0.070 65.695 ;
    RECT 0 65.765 0.070 66.955 ;
    RECT 0 67.025 0.070 68.215 ;
    RECT 0 68.285 0.070 69.475 ;
    RECT 0 69.545 0.070 70.735 ;
    RECT 0 70.805 0.070 71.995 ;
    RECT 0 72.065 0.070 73.255 ;
    RECT 0 73.325 0.070 74.515 ;
    RECT 0 74.585 0.070 75.775 ;
    RECT 0 75.845 0.070 77.035 ;
    RECT 0 77.105 0.070 78.295 ;
    RECT 0 78.365 0.070 79.555 ;
    RECT 0 79.625 0.070 80.815 ;
    RECT 0 80.885 0.070 82.075 ;
    RECT 0 82.145 0.070 83.335 ;
    RECT 0 83.405 0.070 84.595 ;
    RECT 0 84.665 0.070 85.855 ;
    RECT 0 85.925 0.070 87.115 ;
    RECT 0 87.185 0.070 88.375 ;
    RECT 0 88.445 0.070 89.635 ;
    RECT 0 89.705 0.070 90.895 ;
    RECT 0 90.965 0.070 92.155 ;
    RECT 0 92.225 0.070 93.415 ;
    RECT 0 93.485 0.070 94.675 ;
    RECT 0 94.745 0.070 95.935 ;
    RECT 0 96.005 0.070 97.195 ;
    RECT 0 97.265 0.070 98.455 ;
    RECT 0 98.525 0.070 99.715 ;
    RECT 0 99.785 0.070 100.975 ;
    RECT 0 101.045 0.070 102.235 ;
    RECT 0 102.305 0.070 103.495 ;
    RECT 0 103.565 0.070 104.755 ;
    RECT 0 104.825 0.070 106.015 ;
    RECT 0 106.085 0.070 107.275 ;
    RECT 0 107.345 0.070 108.535 ;
    RECT 0 108.605 0.070 109.795 ;
    RECT 0 109.865 0.070 111.055 ;
    RECT 0 111.125 0.070 112.315 ;
    RECT 0 112.385 0.070 113.575 ;
    RECT 0 113.645 0.070 114.835 ;
    RECT 0 114.905 0.070 116.095 ;
    RECT 0 116.165 0.070 117.355 ;
    RECT 0 117.425 0.070 118.615 ;
    RECT 0 118.685 0.070 119.875 ;
    RECT 0 119.945 0.070 121.135 ;
    RECT 0 121.205 0.070 122.395 ;
    RECT 0 122.465 0.070 124.285 ;
    RECT 0 124.355 0.070 125.545 ;
    RECT 0 125.615 0.070 126.805 ;
    RECT 0 126.875 0.070 128.065 ;
    RECT 0 128.135 0.070 129.325 ;
    RECT 0 129.395 0.070 130.585 ;
    RECT 0 130.655 0.070 131.845 ;
    RECT 0 131.915 0.070 133.105 ;
    RECT 0 133.175 0.070 134.365 ;
    RECT 0 134.435 0.070 135.625 ;
    RECT 0 135.695 0.070 136.885 ;
    RECT 0 136.955 0.070 138.145 ;
    RECT 0 138.215 0.070 139.405 ;
    RECT 0 139.475 0.070 140.665 ;
    RECT 0 140.735 0.070 141.925 ;
    RECT 0 141.995 0.070 143.185 ;
    RECT 0 143.255 0.070 144.445 ;
    RECT 0 144.515 0.070 145.705 ;
    RECT 0 145.775 0.070 146.965 ;
    RECT 0 147.035 0.070 148.225 ;
    RECT 0 148.295 0.070 149.485 ;
    RECT 0 149.555 0.070 150.745 ;
    RECT 0 150.815 0.070 152.005 ;
    RECT 0 152.075 0.070 153.265 ;
    RECT 0 153.335 0.070 154.525 ;
    RECT 0 154.595 0.070 155.785 ;
    RECT 0 155.855 0.070 157.045 ;
    RECT 0 157.115 0.070 158.305 ;
    RECT 0 158.375 0.070 159.565 ;
    RECT 0 159.635 0.070 160.825 ;
    RECT 0 160.895 0.070 162.085 ;
    RECT 0 162.155 0.070 163.345 ;
    RECT 0 163.415 0.070 164.605 ;
    RECT 0 164.675 0.070 165.865 ;
    RECT 0 165.935 0.070 167.125 ;
    RECT 0 167.195 0.070 168.385 ;
    RECT 0 168.455 0.070 169.645 ;
    RECT 0 169.715 0.070 170.905 ;
    RECT 0 170.975 0.070 172.165 ;
    RECT 0 172.235 0.070 173.425 ;
    RECT 0 173.495 0.070 174.685 ;
    RECT 0 174.755 0.070 175.945 ;
    RECT 0 176.015 0.070 177.205 ;
    RECT 0 177.275 0.070 178.465 ;
    RECT 0 178.535 0.070 179.725 ;
    RECT 0 179.795 0.070 180.985 ;
    RECT 0 181.055 0.070 182.245 ;
    RECT 0 182.315 0.070 183.505 ;
    RECT 0 183.575 0.070 185.395 ;
    RECT 0 185.465 0.070 186.655 ;
    RECT 0 186.725 0.070 187.915 ;
    RECT 0 187.985 0.070 189.175 ;
    RECT 0 189.245 0.070 190.435 ;
    RECT 0 190.505 0.070 191.695 ;
    RECT 0 191.765 0.070 192.955 ;
    RECT 0 193.025 0.070 194.215 ;
    RECT 0 194.285 0.070 196.105 ;
    RECT 0 196.175 0.070 197.365 ;
    RECT 0 197.435 0.070 198.625 ;
    RECT 0 198.695 0.070 207.200 ;
    LAYER metal4 ;
    RECT 0 0 64.030 2.100 ;
    RECT 0 205.100 64.030 207.200 ;
    RECT 0.000 2.100 1.960 205.100 ;
    RECT 2.240 2.100 3.640 205.100 ;
    RECT 3.920 2.100 5.320 205.100 ;
    RECT 5.600 2.100 7.000 205.100 ;
    RECT 7.280 2.100 8.680 205.100 ;
    RECT 8.960 2.100 10.360 205.100 ;
    RECT 10.640 2.100 12.040 205.100 ;
    RECT 12.320 2.100 13.720 205.100 ;
    RECT 14.000 2.100 15.400 205.100 ;
    RECT 15.680 2.100 17.080 205.100 ;
    RECT 17.360 2.100 18.760 205.100 ;
    RECT 19.040 2.100 20.440 205.100 ;
    RECT 20.720 2.100 22.120 205.100 ;
    RECT 22.400 2.100 23.800 205.100 ;
    RECT 24.080 2.100 25.480 205.100 ;
    RECT 25.760 2.100 27.160 205.100 ;
    RECT 27.440 2.100 28.840 205.100 ;
    RECT 29.120 2.100 30.520 205.100 ;
    RECT 30.800 2.100 32.200 205.100 ;
    RECT 32.480 2.100 33.880 205.100 ;
    RECT 34.160 2.100 35.560 205.100 ;
    RECT 35.840 2.100 37.240 205.100 ;
    RECT 37.520 2.100 38.920 205.100 ;
    RECT 39.200 2.100 40.600 205.100 ;
    RECT 40.880 2.100 42.280 205.100 ;
    RECT 42.560 2.100 43.960 205.100 ;
    RECT 44.240 2.100 45.640 205.100 ;
    RECT 45.920 2.100 47.320 205.100 ;
    RECT 47.600 2.100 49.000 205.100 ;
    RECT 49.280 2.100 50.680 205.100 ;
    RECT 50.960 2.100 52.360 205.100 ;
    RECT 52.640 2.100 54.040 205.100 ;
    RECT 54.320 2.100 55.720 205.100 ;
    RECT 56.000 2.100 57.400 205.100 ;
    RECT 57.680 2.100 59.080 205.100 ;
    RECT 59.360 2.100 60.760 205.100 ;
    RECT 61.040 2.100 64.030 205.100 ;
    LAYER OVERLAP ;
    RECT 0 0 64.030 207.200 ;
  END
END fakeram45_256x48

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_256x34
  FOREIGN fakeram45_256x34 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 98.420 BY 65.800 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.785 0.070 8.855 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.985 0.070 13.055 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.505 0.070 15.575 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[33]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.545 0.070 20.615 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.225 0.070 22.295 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.905 0.070 23.975 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.425 0.070 26.495 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.685 0.070 27.755 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.105 0.070 28.175 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.945 0.070 29.015 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.785 0.070 29.855 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.205 0.070 30.275 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.625 0.070 30.695 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.045 0.070 31.115 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.465 0.070 31.535 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.885 0.070 31.955 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.305 0.070 32.375 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.145 0.070 33.215 ;
    END
  END rd_out[33]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.505 0.070 36.575 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.185 0.070 38.255 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.325 0.070 45.395 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.745 0.070 45.815 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.585 0.070 46.655 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.265 0.070 48.335 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.945 0.070 50.015 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END wd_in[33]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.145 0.070 54.215 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.985 0.070 55.055 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.825 0.070 55.895 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.665 0.070 56.735 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.025 0.070 60.095 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.445 0.070 60.515 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.865 0.070 60.935 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 63.700 ;
      RECT 5.320 2.100 5.600 63.700 ;
      RECT 8.680 2.100 8.960 63.700 ;
      RECT 12.040 2.100 12.320 63.700 ;
      RECT 15.400 2.100 15.680 63.700 ;
      RECT 18.760 2.100 19.040 63.700 ;
      RECT 22.120 2.100 22.400 63.700 ;
      RECT 25.480 2.100 25.760 63.700 ;
      RECT 28.840 2.100 29.120 63.700 ;
      RECT 32.200 2.100 32.480 63.700 ;
      RECT 35.560 2.100 35.840 63.700 ;
      RECT 38.920 2.100 39.200 63.700 ;
      RECT 42.280 2.100 42.560 63.700 ;
      RECT 45.640 2.100 45.920 63.700 ;
      RECT 49.000 2.100 49.280 63.700 ;
      RECT 52.360 2.100 52.640 63.700 ;
      RECT 55.720 2.100 56.000 63.700 ;
      RECT 59.080 2.100 59.360 63.700 ;
      RECT 62.440 2.100 62.720 63.700 ;
      RECT 65.800 2.100 66.080 63.700 ;
      RECT 69.160 2.100 69.440 63.700 ;
      RECT 72.520 2.100 72.800 63.700 ;
      RECT 75.880 2.100 76.160 63.700 ;
      RECT 79.240 2.100 79.520 63.700 ;
      RECT 82.600 2.100 82.880 63.700 ;
      RECT 85.960 2.100 86.240 63.700 ;
      RECT 89.320 2.100 89.600 63.700 ;
      RECT 92.680 2.100 92.960 63.700 ;
      RECT 96.040 2.100 96.320 63.700 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 63.700 ;
      RECT 7.000 2.100 7.280 63.700 ;
      RECT 10.360 2.100 10.640 63.700 ;
      RECT 13.720 2.100 14.000 63.700 ;
      RECT 17.080 2.100 17.360 63.700 ;
      RECT 20.440 2.100 20.720 63.700 ;
      RECT 23.800 2.100 24.080 63.700 ;
      RECT 27.160 2.100 27.440 63.700 ;
      RECT 30.520 2.100 30.800 63.700 ;
      RECT 33.880 2.100 34.160 63.700 ;
      RECT 37.240 2.100 37.520 63.700 ;
      RECT 40.600 2.100 40.880 63.700 ;
      RECT 43.960 2.100 44.240 63.700 ;
      RECT 47.320 2.100 47.600 63.700 ;
      RECT 50.680 2.100 50.960 63.700 ;
      RECT 54.040 2.100 54.320 63.700 ;
      RECT 57.400 2.100 57.680 63.700 ;
      RECT 60.760 2.100 61.040 63.700 ;
      RECT 64.120 2.100 64.400 63.700 ;
      RECT 67.480 2.100 67.760 63.700 ;
      RECT 70.840 2.100 71.120 63.700 ;
      RECT 74.200 2.100 74.480 63.700 ;
      RECT 77.560 2.100 77.840 63.700 ;
      RECT 80.920 2.100 81.200 63.700 ;
      RECT 84.280 2.100 84.560 63.700 ;
      RECT 87.640 2.100 87.920 63.700 ;
      RECT 91.000 2.100 91.280 63.700 ;
      RECT 94.360 2.100 94.640 63.700 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 98.420 65.800 ;
    LAYER metal2 ;
    RECT 0 0 98.420 65.800 ;
    LAYER metal3 ;
    RECT 0.070 0 98.420 65.800 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.485 ;
    RECT 0 2.555 0.070 2.905 ;
    RECT 0 2.975 0.070 3.325 ;
    RECT 0 3.395 0.070 3.745 ;
    RECT 0 3.815 0.070 4.165 ;
    RECT 0 4.235 0.070 4.585 ;
    RECT 0 4.655 0.070 5.005 ;
    RECT 0 5.075 0.070 5.425 ;
    RECT 0 5.495 0.070 5.845 ;
    RECT 0 5.915 0.070 6.265 ;
    RECT 0 6.335 0.070 6.685 ;
    RECT 0 6.755 0.070 7.105 ;
    RECT 0 7.175 0.070 7.525 ;
    RECT 0 7.595 0.070 7.945 ;
    RECT 0 8.015 0.070 8.365 ;
    RECT 0 8.435 0.070 8.785 ;
    RECT 0 8.855 0.070 9.205 ;
    RECT 0 9.275 0.070 9.625 ;
    RECT 0 9.695 0.070 10.045 ;
    RECT 0 10.115 0.070 10.465 ;
    RECT 0 10.535 0.070 10.885 ;
    RECT 0 10.955 0.070 11.305 ;
    RECT 0 11.375 0.070 11.725 ;
    RECT 0 11.795 0.070 12.145 ;
    RECT 0 12.215 0.070 12.565 ;
    RECT 0 12.635 0.070 12.985 ;
    RECT 0 13.055 0.070 13.405 ;
    RECT 0 13.475 0.070 13.825 ;
    RECT 0 13.895 0.070 14.245 ;
    RECT 0 14.315 0.070 14.665 ;
    RECT 0 14.735 0.070 15.085 ;
    RECT 0 15.155 0.070 15.505 ;
    RECT 0 15.575 0.070 15.925 ;
    RECT 0 15.995 0.070 19.285 ;
    RECT 0 19.355 0.070 19.705 ;
    RECT 0 19.775 0.070 20.125 ;
    RECT 0 20.195 0.070 20.545 ;
    RECT 0 20.615 0.070 20.965 ;
    RECT 0 21.035 0.070 21.385 ;
    RECT 0 21.455 0.070 21.805 ;
    RECT 0 21.875 0.070 22.225 ;
    RECT 0 22.295 0.070 22.645 ;
    RECT 0 22.715 0.070 23.065 ;
    RECT 0 23.135 0.070 23.485 ;
    RECT 0 23.555 0.070 23.905 ;
    RECT 0 23.975 0.070 24.325 ;
    RECT 0 24.395 0.070 24.745 ;
    RECT 0 24.815 0.070 25.165 ;
    RECT 0 25.235 0.070 25.585 ;
    RECT 0 25.655 0.070 26.005 ;
    RECT 0 26.075 0.070 26.425 ;
    RECT 0 26.495 0.070 26.845 ;
    RECT 0 26.915 0.070 27.265 ;
    RECT 0 27.335 0.070 27.685 ;
    RECT 0 27.755 0.070 28.105 ;
    RECT 0 28.175 0.070 28.525 ;
    RECT 0 28.595 0.070 28.945 ;
    RECT 0 29.015 0.070 29.365 ;
    RECT 0 29.435 0.070 29.785 ;
    RECT 0 29.855 0.070 30.205 ;
    RECT 0 30.275 0.070 30.625 ;
    RECT 0 30.695 0.070 31.045 ;
    RECT 0 31.115 0.070 31.465 ;
    RECT 0 31.535 0.070 31.885 ;
    RECT 0 31.955 0.070 32.305 ;
    RECT 0 32.375 0.070 32.725 ;
    RECT 0 32.795 0.070 33.145 ;
    RECT 0 33.215 0.070 36.505 ;
    RECT 0 36.575 0.070 36.925 ;
    RECT 0 36.995 0.070 37.345 ;
    RECT 0 37.415 0.070 37.765 ;
    RECT 0 37.835 0.070 38.185 ;
    RECT 0 38.255 0.070 38.605 ;
    RECT 0 38.675 0.070 39.025 ;
    RECT 0 39.095 0.070 39.445 ;
    RECT 0 39.515 0.070 39.865 ;
    RECT 0 39.935 0.070 40.285 ;
    RECT 0 40.355 0.070 40.705 ;
    RECT 0 40.775 0.070 41.125 ;
    RECT 0 41.195 0.070 41.545 ;
    RECT 0 41.615 0.070 41.965 ;
    RECT 0 42.035 0.070 42.385 ;
    RECT 0 42.455 0.070 42.805 ;
    RECT 0 42.875 0.070 43.225 ;
    RECT 0 43.295 0.070 43.645 ;
    RECT 0 43.715 0.070 44.065 ;
    RECT 0 44.135 0.070 44.485 ;
    RECT 0 44.555 0.070 44.905 ;
    RECT 0 44.975 0.070 45.325 ;
    RECT 0 45.395 0.070 45.745 ;
    RECT 0 45.815 0.070 46.165 ;
    RECT 0 46.235 0.070 46.585 ;
    RECT 0 46.655 0.070 47.005 ;
    RECT 0 47.075 0.070 47.425 ;
    RECT 0 47.495 0.070 47.845 ;
    RECT 0 47.915 0.070 48.265 ;
    RECT 0 48.335 0.070 48.685 ;
    RECT 0 48.755 0.070 49.105 ;
    RECT 0 49.175 0.070 49.525 ;
    RECT 0 49.595 0.070 49.945 ;
    RECT 0 50.015 0.070 50.365 ;
    RECT 0 50.435 0.070 53.725 ;
    RECT 0 53.795 0.070 54.145 ;
    RECT 0 54.215 0.070 54.565 ;
    RECT 0 54.635 0.070 54.985 ;
    RECT 0 55.055 0.070 55.405 ;
    RECT 0 55.475 0.070 55.825 ;
    RECT 0 55.895 0.070 56.245 ;
    RECT 0 56.315 0.070 56.665 ;
    RECT 0 56.735 0.070 60.025 ;
    RECT 0 60.095 0.070 60.445 ;
    RECT 0 60.515 0.070 60.865 ;
    RECT 0 60.935 0.070 65.800 ;
    LAYER metal4 ;
    RECT 0 0 98.420 2.100 ;
    RECT 0 63.700 98.420 65.800 ;
    RECT 0.000 2.100 1.960 63.700 ;
    RECT 2.240 2.100 3.640 63.700 ;
    RECT 3.920 2.100 5.320 63.700 ;
    RECT 5.600 2.100 7.000 63.700 ;
    RECT 7.280 2.100 8.680 63.700 ;
    RECT 8.960 2.100 10.360 63.700 ;
    RECT 10.640 2.100 12.040 63.700 ;
    RECT 12.320 2.100 13.720 63.700 ;
    RECT 14.000 2.100 15.400 63.700 ;
    RECT 15.680 2.100 17.080 63.700 ;
    RECT 17.360 2.100 18.760 63.700 ;
    RECT 19.040 2.100 20.440 63.700 ;
    RECT 20.720 2.100 22.120 63.700 ;
    RECT 22.400 2.100 23.800 63.700 ;
    RECT 24.080 2.100 25.480 63.700 ;
    RECT 25.760 2.100 27.160 63.700 ;
    RECT 27.440 2.100 28.840 63.700 ;
    RECT 29.120 2.100 30.520 63.700 ;
    RECT 30.800 2.100 32.200 63.700 ;
    RECT 32.480 2.100 33.880 63.700 ;
    RECT 34.160 2.100 35.560 63.700 ;
    RECT 35.840 2.100 37.240 63.700 ;
    RECT 37.520 2.100 38.920 63.700 ;
    RECT 39.200 2.100 40.600 63.700 ;
    RECT 40.880 2.100 42.280 63.700 ;
    RECT 42.560 2.100 43.960 63.700 ;
    RECT 44.240 2.100 45.640 63.700 ;
    RECT 45.920 2.100 47.320 63.700 ;
    RECT 47.600 2.100 49.000 63.700 ;
    RECT 49.280 2.100 50.680 63.700 ;
    RECT 50.960 2.100 52.360 63.700 ;
    RECT 52.640 2.100 54.040 63.700 ;
    RECT 54.320 2.100 55.720 63.700 ;
    RECT 56.000 2.100 57.400 63.700 ;
    RECT 57.680 2.100 59.080 63.700 ;
    RECT 59.360 2.100 60.760 63.700 ;
    RECT 61.040 2.100 62.440 63.700 ;
    RECT 62.720 2.100 64.120 63.700 ;
    RECT 64.400 2.100 65.800 63.700 ;
    RECT 66.080 2.100 67.480 63.700 ;
    RECT 67.760 2.100 69.160 63.700 ;
    RECT 69.440 2.100 70.840 63.700 ;
    RECT 71.120 2.100 72.520 63.700 ;
    RECT 72.800 2.100 74.200 63.700 ;
    RECT 74.480 2.100 75.880 63.700 ;
    RECT 76.160 2.100 77.560 63.700 ;
    RECT 77.840 2.100 79.240 63.700 ;
    RECT 79.520 2.100 80.920 63.700 ;
    RECT 81.200 2.100 82.600 63.700 ;
    RECT 82.880 2.100 84.280 63.700 ;
    RECT 84.560 2.100 85.960 63.700 ;
    RECT 86.240 2.100 87.640 63.700 ;
    RECT 87.920 2.100 89.320 63.700 ;
    RECT 89.600 2.100 91.000 63.700 ;
    RECT 91.280 2.100 92.680 63.700 ;
    RECT 92.960 2.100 94.360 63.700 ;
    RECT 94.640 2.100 96.040 63.700 ;
    RECT 96.320 2.100 98.420 63.700 ;
    LAYER OVERLAP ;
    RECT 0 0 98.420 65.800 ;
  END
END fakeram45_256x34

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_256x32
  FOREIGN fakeram45_256x32 0 0 ;
  SYMMETRY X Y ;
  SIZE 60.610 BY 169.400 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.535 0.070 3.605 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.475 0.070 6.545 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.415 0.070 9.485 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.355 0.070 12.425 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.295 0.070 15.365 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.235 0.070 18.305 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.175 0.070 21.245 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.115 0.070 24.185 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.055 0.070 27.125 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.995 0.070 30.065 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.465 0.070 31.535 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.935 0.070 33.005 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.875 0.070 35.945 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.815 0.070 38.885 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.755 0.070 41.825 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.695 0.070 44.765 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.635 0.070 47.705 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.995 0.070 51.065 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.935 0.070 54.005 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.875 0.070 56.945 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.345 0.070 58.415 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.815 0.070 59.885 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.285 0.070 61.355 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.755 0.070 62.825 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.225 0.070 64.295 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.695 0.070 65.765 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.165 0.070 67.235 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.635 0.070 68.705 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.105 0.070 70.175 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.575 0.070 71.645 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.515 0.070 74.585 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.455 0.070 77.525 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.925 0.070 78.995 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.395 0.070 80.465 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.335 0.070 83.405 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.275 0.070 86.345 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.745 0.070 87.815 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.215 0.070 89.285 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.685 0.070 90.755 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.155 0.070 92.225 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.625 0.070 93.695 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.095 0.070 95.165 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.985 0.070 97.055 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.455 0.070 98.525 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.925 0.070 99.995 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.395 0.070 101.465 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.865 0.070 102.935 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.335 0.070 104.405 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.805 0.070 105.875 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.275 0.070 107.345 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.745 0.070 108.815 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.215 0.070 110.285 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.685 0.070 111.755 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.155 0.070 113.225 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.625 0.070 114.695 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.095 0.070 116.165 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.565 0.070 117.635 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.035 0.070 119.105 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.505 0.070 120.575 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.975 0.070 122.045 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.445 0.070 123.515 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.915 0.070 124.985 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.385 0.070 126.455 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.855 0.070 127.925 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.325 0.070 129.395 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.795 0.070 130.865 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.265 0.070 132.335 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.735 0.070 133.805 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.205 0.070 135.275 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.675 0.070 136.745 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.145 0.070 138.215 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.615 0.070 139.685 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.085 0.070 141.155 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.555 0.070 142.625 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.445 0.070 144.515 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.915 0.070 145.985 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.385 0.070 147.455 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.855 0.070 148.925 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.325 0.070 150.395 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.795 0.070 151.865 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.265 0.070 153.335 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.735 0.070 154.805 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.625 0.070 156.695 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.095 0.070 158.165 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.565 0.070 159.635 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 167.300 ;
      RECT 5.320 2.100 5.600 167.300 ;
      RECT 8.680 2.100 8.960 167.300 ;
      RECT 12.040 2.100 12.320 167.300 ;
      RECT 15.400 2.100 15.680 167.300 ;
      RECT 18.760 2.100 19.040 167.300 ;
      RECT 22.120 2.100 22.400 167.300 ;
      RECT 25.480 2.100 25.760 167.300 ;
      RECT 28.840 2.100 29.120 167.300 ;
      RECT 32.200 2.100 32.480 167.300 ;
      RECT 35.560 2.100 35.840 167.300 ;
      RECT 38.920 2.100 39.200 167.300 ;
      RECT 42.280 2.100 42.560 167.300 ;
      RECT 45.640 2.100 45.920 167.300 ;
      RECT 49.000 2.100 49.280 167.300 ;
      RECT 52.360 2.100 52.640 167.300 ;
      RECT 55.720 2.100 56.000 167.300 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 167.300 ;
      RECT 7.000 2.100 7.280 167.300 ;
      RECT 10.360 2.100 10.640 167.300 ;
      RECT 13.720 2.100 14.000 167.300 ;
      RECT 17.080 2.100 17.360 167.300 ;
      RECT 20.440 2.100 20.720 167.300 ;
      RECT 23.800 2.100 24.080 167.300 ;
      RECT 27.160 2.100 27.440 167.300 ;
      RECT 30.520 2.100 30.800 167.300 ;
      RECT 33.880 2.100 34.160 167.300 ;
      RECT 37.240 2.100 37.520 167.300 ;
      RECT 40.600 2.100 40.880 167.300 ;
      RECT 43.960 2.100 44.240 167.300 ;
      RECT 47.320 2.100 47.600 167.300 ;
      RECT 50.680 2.100 50.960 167.300 ;
      RECT 54.040 2.100 54.320 167.300 ;
      RECT 57.400 2.100 57.680 167.300 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 60.610 169.400 ;
    LAYER metal2 ;
    RECT 0 0 60.610 169.400 ;
    LAYER metal3 ;
    RECT 0.070 0 60.610 169.400 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 3.535 ;
    RECT 0 3.605 0.070 5.005 ;
    RECT 0 5.075 0.070 6.475 ;
    RECT 0 6.545 0.070 7.945 ;
    RECT 0 8.015 0.070 9.415 ;
    RECT 0 9.485 0.070 10.885 ;
    RECT 0 10.955 0.070 12.355 ;
    RECT 0 12.425 0.070 13.825 ;
    RECT 0 13.895 0.070 15.295 ;
    RECT 0 15.365 0.070 16.765 ;
    RECT 0 16.835 0.070 18.235 ;
    RECT 0 18.305 0.070 19.705 ;
    RECT 0 19.775 0.070 21.175 ;
    RECT 0 21.245 0.070 22.645 ;
    RECT 0 22.715 0.070 24.115 ;
    RECT 0 24.185 0.070 25.585 ;
    RECT 0 25.655 0.070 27.055 ;
    RECT 0 27.125 0.070 28.525 ;
    RECT 0 28.595 0.070 29.995 ;
    RECT 0 30.065 0.070 31.465 ;
    RECT 0 31.535 0.070 32.935 ;
    RECT 0 33.005 0.070 34.405 ;
    RECT 0 34.475 0.070 35.875 ;
    RECT 0 35.945 0.070 37.345 ;
    RECT 0 37.415 0.070 38.815 ;
    RECT 0 38.885 0.070 40.285 ;
    RECT 0 40.355 0.070 41.755 ;
    RECT 0 41.825 0.070 43.225 ;
    RECT 0 43.295 0.070 44.695 ;
    RECT 0 44.765 0.070 46.165 ;
    RECT 0 46.235 0.070 47.635 ;
    RECT 0 47.705 0.070 49.525 ;
    RECT 0 49.595 0.070 50.995 ;
    RECT 0 51.065 0.070 52.465 ;
    RECT 0 52.535 0.070 53.935 ;
    RECT 0 54.005 0.070 55.405 ;
    RECT 0 55.475 0.070 56.875 ;
    RECT 0 56.945 0.070 58.345 ;
    RECT 0 58.415 0.070 59.815 ;
    RECT 0 59.885 0.070 61.285 ;
    RECT 0 61.355 0.070 62.755 ;
    RECT 0 62.825 0.070 64.225 ;
    RECT 0 64.295 0.070 65.695 ;
    RECT 0 65.765 0.070 67.165 ;
    RECT 0 67.235 0.070 68.635 ;
    RECT 0 68.705 0.070 70.105 ;
    RECT 0 70.175 0.070 71.575 ;
    RECT 0 71.645 0.070 73.045 ;
    RECT 0 73.115 0.070 74.515 ;
    RECT 0 74.585 0.070 75.985 ;
    RECT 0 76.055 0.070 77.455 ;
    RECT 0 77.525 0.070 78.925 ;
    RECT 0 78.995 0.070 80.395 ;
    RECT 0 80.465 0.070 81.865 ;
    RECT 0 81.935 0.070 83.335 ;
    RECT 0 83.405 0.070 84.805 ;
    RECT 0 84.875 0.070 86.275 ;
    RECT 0 86.345 0.070 87.745 ;
    RECT 0 87.815 0.070 89.215 ;
    RECT 0 89.285 0.070 90.685 ;
    RECT 0 90.755 0.070 92.155 ;
    RECT 0 92.225 0.070 93.625 ;
    RECT 0 93.695 0.070 95.095 ;
    RECT 0 95.165 0.070 96.985 ;
    RECT 0 97.055 0.070 98.455 ;
    RECT 0 98.525 0.070 99.925 ;
    RECT 0 99.995 0.070 101.395 ;
    RECT 0 101.465 0.070 102.865 ;
    RECT 0 102.935 0.070 104.335 ;
    RECT 0 104.405 0.070 105.805 ;
    RECT 0 105.875 0.070 107.275 ;
    RECT 0 107.345 0.070 108.745 ;
    RECT 0 108.815 0.070 110.215 ;
    RECT 0 110.285 0.070 111.685 ;
    RECT 0 111.755 0.070 113.155 ;
    RECT 0 113.225 0.070 114.625 ;
    RECT 0 114.695 0.070 116.095 ;
    RECT 0 116.165 0.070 117.565 ;
    RECT 0 117.635 0.070 119.035 ;
    RECT 0 119.105 0.070 120.505 ;
    RECT 0 120.575 0.070 121.975 ;
    RECT 0 122.045 0.070 123.445 ;
    RECT 0 123.515 0.070 124.915 ;
    RECT 0 124.985 0.070 126.385 ;
    RECT 0 126.455 0.070 127.855 ;
    RECT 0 127.925 0.070 129.325 ;
    RECT 0 129.395 0.070 130.795 ;
    RECT 0 130.865 0.070 132.265 ;
    RECT 0 132.335 0.070 133.735 ;
    RECT 0 133.805 0.070 135.205 ;
    RECT 0 135.275 0.070 136.675 ;
    RECT 0 136.745 0.070 138.145 ;
    RECT 0 138.215 0.070 139.615 ;
    RECT 0 139.685 0.070 141.085 ;
    RECT 0 141.155 0.070 142.555 ;
    RECT 0 142.625 0.070 144.445 ;
    RECT 0 144.515 0.070 145.915 ;
    RECT 0 145.985 0.070 147.385 ;
    RECT 0 147.455 0.070 148.855 ;
    RECT 0 148.925 0.070 150.325 ;
    RECT 0 150.395 0.070 151.795 ;
    RECT 0 151.865 0.070 153.265 ;
    RECT 0 153.335 0.070 154.735 ;
    RECT 0 154.805 0.070 156.625 ;
    RECT 0 156.695 0.070 158.095 ;
    RECT 0 158.165 0.070 159.565 ;
    RECT 0 159.635 0.070 169.400 ;
    LAYER metal4 ;
    RECT 0 0 60.610 2.100 ;
    RECT 0 167.300 60.610 169.400 ;
    RECT 0.000 2.100 1.960 167.300 ;
    RECT 2.240 2.100 3.640 167.300 ;
    RECT 3.920 2.100 5.320 167.300 ;
    RECT 5.600 2.100 7.000 167.300 ;
    RECT 7.280 2.100 8.680 167.300 ;
    RECT 8.960 2.100 10.360 167.300 ;
    RECT 10.640 2.100 12.040 167.300 ;
    RECT 12.320 2.100 13.720 167.300 ;
    RECT 14.000 2.100 15.400 167.300 ;
    RECT 15.680 2.100 17.080 167.300 ;
    RECT 17.360 2.100 18.760 167.300 ;
    RECT 19.040 2.100 20.440 167.300 ;
    RECT 20.720 2.100 22.120 167.300 ;
    RECT 22.400 2.100 23.800 167.300 ;
    RECT 24.080 2.100 25.480 167.300 ;
    RECT 25.760 2.100 27.160 167.300 ;
    RECT 27.440 2.100 28.840 167.300 ;
    RECT 29.120 2.100 30.520 167.300 ;
    RECT 30.800 2.100 32.200 167.300 ;
    RECT 32.480 2.100 33.880 167.300 ;
    RECT 34.160 2.100 35.560 167.300 ;
    RECT 35.840 2.100 37.240 167.300 ;
    RECT 37.520 2.100 38.920 167.300 ;
    RECT 39.200 2.100 40.600 167.300 ;
    RECT 40.880 2.100 42.280 167.300 ;
    RECT 42.560 2.100 43.960 167.300 ;
    RECT 44.240 2.100 45.640 167.300 ;
    RECT 45.920 2.100 47.320 167.300 ;
    RECT 47.600 2.100 49.000 167.300 ;
    RECT 49.280 2.100 50.680 167.300 ;
    RECT 50.960 2.100 52.360 167.300 ;
    RECT 52.640 2.100 54.040 167.300 ;
    RECT 54.320 2.100 55.720 167.300 ;
    RECT 56.000 2.100 57.400 167.300 ;
    RECT 57.680 2.100 60.610 167.300 ;
    LAYER OVERLAP ;
    RECT 0 0 60.610 169.400 ;
  END
END fakeram45_256x32

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_256x16
  FOREIGN fakeram45_256x16 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 77.710 BY 40.600 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[15]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.095 0.070 11.165 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.515 0.070 11.585 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.935 0.070 12.005 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.355 0.070 12.425 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.775 0.070 12.845 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.195 0.070 13.265 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.615 0.070 13.685 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.035 0.070 14.105 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.455 0.070 14.525 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.875 0.070 14.945 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.295 0.070 15.365 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.715 0.070 15.785 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.135 0.070 16.205 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.555 0.070 16.625 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.975 0.070 17.045 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.395 0.070 17.465 ;
    END
  END rd_out[15]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.545 0.070 20.615 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.225 0.070 22.295 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.905 0.070 23.975 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.425 0.070 26.495 ;
    END
  END wd_in[15]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.155 0.070 29.225 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.575 0.070 29.645 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.995 0.070 30.065 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.415 0.070 30.485 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.835 0.070 30.905 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.255 0.070 31.325 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.675 0.070 31.745 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.095 0.070 32.165 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.825 0.070 34.895 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 38.500 ;
      RECT 5.320 2.100 5.600 38.500 ;
      RECT 8.680 2.100 8.960 38.500 ;
      RECT 12.040 2.100 12.320 38.500 ;
      RECT 15.400 2.100 15.680 38.500 ;
      RECT 18.760 2.100 19.040 38.500 ;
      RECT 22.120 2.100 22.400 38.500 ;
      RECT 25.480 2.100 25.760 38.500 ;
      RECT 28.840 2.100 29.120 38.500 ;
      RECT 32.200 2.100 32.480 38.500 ;
      RECT 35.560 2.100 35.840 38.500 ;
      RECT 38.920 2.100 39.200 38.500 ;
      RECT 42.280 2.100 42.560 38.500 ;
      RECT 45.640 2.100 45.920 38.500 ;
      RECT 49.000 2.100 49.280 38.500 ;
      RECT 52.360 2.100 52.640 38.500 ;
      RECT 55.720 2.100 56.000 38.500 ;
      RECT 59.080 2.100 59.360 38.500 ;
      RECT 62.440 2.100 62.720 38.500 ;
      RECT 65.800 2.100 66.080 38.500 ;
      RECT 69.160 2.100 69.440 38.500 ;
      RECT 72.520 2.100 72.800 38.500 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 38.500 ;
      RECT 7.000 2.100 7.280 38.500 ;
      RECT 10.360 2.100 10.640 38.500 ;
      RECT 13.720 2.100 14.000 38.500 ;
      RECT 17.080 2.100 17.360 38.500 ;
      RECT 20.440 2.100 20.720 38.500 ;
      RECT 23.800 2.100 24.080 38.500 ;
      RECT 27.160 2.100 27.440 38.500 ;
      RECT 30.520 2.100 30.800 38.500 ;
      RECT 33.880 2.100 34.160 38.500 ;
      RECT 37.240 2.100 37.520 38.500 ;
      RECT 40.600 2.100 40.880 38.500 ;
      RECT 43.960 2.100 44.240 38.500 ;
      RECT 47.320 2.100 47.600 38.500 ;
      RECT 50.680 2.100 50.960 38.500 ;
      RECT 54.040 2.100 54.320 38.500 ;
      RECT 57.400 2.100 57.680 38.500 ;
      RECT 60.760 2.100 61.040 38.500 ;
      RECT 64.120 2.100 64.400 38.500 ;
      RECT 67.480 2.100 67.760 38.500 ;
      RECT 70.840 2.100 71.120 38.500 ;
      RECT 74.200 2.100 74.480 38.500 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 77.710 40.600 ;
    LAYER metal2 ;
    RECT 0 0 77.710 40.600 ;
    LAYER metal3 ;
    RECT 0.070 0 77.710 40.600 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.485 ;
    RECT 0 2.555 0.070 2.905 ;
    RECT 0 2.975 0.070 3.325 ;
    RECT 0 3.395 0.070 3.745 ;
    RECT 0 3.815 0.070 4.165 ;
    RECT 0 4.235 0.070 4.585 ;
    RECT 0 4.655 0.070 5.005 ;
    RECT 0 5.075 0.070 5.425 ;
    RECT 0 5.495 0.070 5.845 ;
    RECT 0 5.915 0.070 6.265 ;
    RECT 0 6.335 0.070 6.685 ;
    RECT 0 6.755 0.070 7.105 ;
    RECT 0 7.175 0.070 7.525 ;
    RECT 0 7.595 0.070 7.945 ;
    RECT 0 8.015 0.070 8.365 ;
    RECT 0 8.435 0.070 11.095 ;
    RECT 0 11.165 0.070 11.515 ;
    RECT 0 11.585 0.070 11.935 ;
    RECT 0 12.005 0.070 12.355 ;
    RECT 0 12.425 0.070 12.775 ;
    RECT 0 12.845 0.070 13.195 ;
    RECT 0 13.265 0.070 13.615 ;
    RECT 0 13.685 0.070 14.035 ;
    RECT 0 14.105 0.070 14.455 ;
    RECT 0 14.525 0.070 14.875 ;
    RECT 0 14.945 0.070 15.295 ;
    RECT 0 15.365 0.070 15.715 ;
    RECT 0 15.785 0.070 16.135 ;
    RECT 0 16.205 0.070 16.555 ;
    RECT 0 16.625 0.070 16.975 ;
    RECT 0 17.045 0.070 17.395 ;
    RECT 0 17.465 0.070 20.125 ;
    RECT 0 20.195 0.070 20.545 ;
    RECT 0 20.615 0.070 20.965 ;
    RECT 0 21.035 0.070 21.385 ;
    RECT 0 21.455 0.070 21.805 ;
    RECT 0 21.875 0.070 22.225 ;
    RECT 0 22.295 0.070 22.645 ;
    RECT 0 22.715 0.070 23.065 ;
    RECT 0 23.135 0.070 23.485 ;
    RECT 0 23.555 0.070 23.905 ;
    RECT 0 23.975 0.070 24.325 ;
    RECT 0 24.395 0.070 24.745 ;
    RECT 0 24.815 0.070 25.165 ;
    RECT 0 25.235 0.070 25.585 ;
    RECT 0 25.655 0.070 26.005 ;
    RECT 0 26.075 0.070 26.425 ;
    RECT 0 26.495 0.070 29.155 ;
    RECT 0 29.225 0.070 29.575 ;
    RECT 0 29.645 0.070 29.995 ;
    RECT 0 30.065 0.070 30.415 ;
    RECT 0 30.485 0.070 30.835 ;
    RECT 0 30.905 0.070 31.255 ;
    RECT 0 31.325 0.070 31.675 ;
    RECT 0 31.745 0.070 32.095 ;
    RECT 0 32.165 0.070 34.825 ;
    RECT 0 34.895 0.070 35.245 ;
    RECT 0 35.315 0.070 35.665 ;
    RECT 0 35.735 0.070 40.600 ;
    LAYER metal4 ;
    RECT 0 0 77.710 2.100 ;
    RECT 0 38.500 77.710 40.600 ;
    RECT 0.000 2.100 1.960 38.500 ;
    RECT 2.240 2.100 3.640 38.500 ;
    RECT 3.920 2.100 5.320 38.500 ;
    RECT 5.600 2.100 7.000 38.500 ;
    RECT 7.280 2.100 8.680 38.500 ;
    RECT 8.960 2.100 10.360 38.500 ;
    RECT 10.640 2.100 12.040 38.500 ;
    RECT 12.320 2.100 13.720 38.500 ;
    RECT 14.000 2.100 15.400 38.500 ;
    RECT 15.680 2.100 17.080 38.500 ;
    RECT 17.360 2.100 18.760 38.500 ;
    RECT 19.040 2.100 20.440 38.500 ;
    RECT 20.720 2.100 22.120 38.500 ;
    RECT 22.400 2.100 23.800 38.500 ;
    RECT 24.080 2.100 25.480 38.500 ;
    RECT 25.760 2.100 27.160 38.500 ;
    RECT 27.440 2.100 28.840 38.500 ;
    RECT 29.120 2.100 30.520 38.500 ;
    RECT 30.800 2.100 32.200 38.500 ;
    RECT 32.480 2.100 33.880 38.500 ;
    RECT 34.160 2.100 35.560 38.500 ;
    RECT 35.840 2.100 37.240 38.500 ;
    RECT 37.520 2.100 38.920 38.500 ;
    RECT 39.200 2.100 40.600 38.500 ;
    RECT 40.880 2.100 42.280 38.500 ;
    RECT 42.560 2.100 43.960 38.500 ;
    RECT 44.240 2.100 45.640 38.500 ;
    RECT 45.920 2.100 47.320 38.500 ;
    RECT 47.600 2.100 49.000 38.500 ;
    RECT 49.280 2.100 50.680 38.500 ;
    RECT 50.960 2.100 52.360 38.500 ;
    RECT 52.640 2.100 54.040 38.500 ;
    RECT 54.320 2.100 55.720 38.500 ;
    RECT 56.000 2.100 57.400 38.500 ;
    RECT 57.680 2.100 59.080 38.500 ;
    RECT 59.360 2.100 60.760 38.500 ;
    RECT 61.040 2.100 62.440 38.500 ;
    RECT 62.720 2.100 64.120 38.500 ;
    RECT 64.400 2.100 65.800 38.500 ;
    RECT 66.080 2.100 67.480 38.500 ;
    RECT 67.760 2.100 69.160 38.500 ;
    RECT 69.440 2.100 70.840 38.500 ;
    RECT 71.120 2.100 72.520 38.500 ;
    RECT 72.800 2.100 74.200 38.500 ;
    RECT 74.480 2.100 77.710 38.500 ;
    LAYER OVERLAP ;
    RECT 0 0 77.710 40.600 ;
  END
END fakeram45_256x16

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_128x256
  FOREIGN fakeram45_128x256 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 153.710 BY 238.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.275 0.070 2.345 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.695 0.070 2.765 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.115 0.070 3.185 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.535 0.070 3.605 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.955 0.070 4.025 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.375 0.070 4.445 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.795 0.070 4.865 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.215 0.070 5.285 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.635 0.070 5.705 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.055 0.070 6.125 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.475 0.070 6.545 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.895 0.070 6.965 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.315 0.070 7.385 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.735 0.070 7.805 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.155 0.070 8.225 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.575 0.070 8.645 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.785 0.070 8.855 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.995 0.070 9.065 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.415 0.070 9.485 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.835 0.070 9.905 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.255 0.070 10.325 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.675 0.070 10.745 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.095 0.070 11.165 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.515 0.070 11.585 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.935 0.070 12.005 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.355 0.070 12.425 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.775 0.070 12.845 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.985 0.070 13.055 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.195 0.070 13.265 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.615 0.070 13.685 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.035 0.070 14.105 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.455 0.070 14.525 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.875 0.070 14.945 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.295 0.070 15.365 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.505 0.070 15.575 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.715 0.070 15.785 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.135 0.070 16.205 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.345 0.070 16.415 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.555 0.070 16.625 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.975 0.070 17.045 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.185 0.070 17.255 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.395 0.070 17.465 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.605 0.070 17.675 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.815 0.070 17.885 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.025 0.070 18.095 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.235 0.070 18.305 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.655 0.070 18.725 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.075 0.070 19.145 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.495 0.070 19.565 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.915 0.070 19.985 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.335 0.070 20.405 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.545 0.070 20.615 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.755 0.070 20.825 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.175 0.070 21.245 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.595 0.070 21.665 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.015 0.070 22.085 ;
    END
  END w_mask_in[95]
  PIN w_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.225 0.070 22.295 ;
    END
  END w_mask_in[96]
  PIN w_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.435 0.070 22.505 ;
    END
  END w_mask_in[97]
  PIN w_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END w_mask_in[98]
  PIN w_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.855 0.070 22.925 ;
    END
  END w_mask_in[99]
  PIN w_mask_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END w_mask_in[100]
  PIN w_mask_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.275 0.070 23.345 ;
    END
  END w_mask_in[101]
  PIN w_mask_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END w_mask_in[102]
  PIN w_mask_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.695 0.070 23.765 ;
    END
  END w_mask_in[103]
  PIN w_mask_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.905 0.070 23.975 ;
    END
  END w_mask_in[104]
  PIN w_mask_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.115 0.070 24.185 ;
    END
  END w_mask_in[105]
  PIN w_mask_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END w_mask_in[106]
  PIN w_mask_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.535 0.070 24.605 ;
    END
  END w_mask_in[107]
  PIN w_mask_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END w_mask_in[108]
  PIN w_mask_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.955 0.070 25.025 ;
    END
  END w_mask_in[109]
  PIN w_mask_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END w_mask_in[110]
  PIN w_mask_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.375 0.070 25.445 ;
    END
  END w_mask_in[111]
  PIN w_mask_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END w_mask_in[112]
  PIN w_mask_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.795 0.070 25.865 ;
    END
  END w_mask_in[113]
  PIN w_mask_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END w_mask_in[114]
  PIN w_mask_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.215 0.070 26.285 ;
    END
  END w_mask_in[115]
  PIN w_mask_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.425 0.070 26.495 ;
    END
  END w_mask_in[116]
  PIN w_mask_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.635 0.070 26.705 ;
    END
  END w_mask_in[117]
  PIN w_mask_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END w_mask_in[118]
  PIN w_mask_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.055 0.070 27.125 ;
    END
  END w_mask_in[119]
  PIN w_mask_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END w_mask_in[120]
  PIN w_mask_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.475 0.070 27.545 ;
    END
  END w_mask_in[121]
  PIN w_mask_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.685 0.070 27.755 ;
    END
  END w_mask_in[122]
  PIN w_mask_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.895 0.070 27.965 ;
    END
  END w_mask_in[123]
  PIN w_mask_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.105 0.070 28.175 ;
    END
  END w_mask_in[124]
  PIN w_mask_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.315 0.070 28.385 ;
    END
  END w_mask_in[125]
  PIN w_mask_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END w_mask_in[126]
  PIN w_mask_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.735 0.070 28.805 ;
    END
  END w_mask_in[127]
  PIN w_mask_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.945 0.070 29.015 ;
    END
  END w_mask_in[128]
  PIN w_mask_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.155 0.070 29.225 ;
    END
  END w_mask_in[129]
  PIN w_mask_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END w_mask_in[130]
  PIN w_mask_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.575 0.070 29.645 ;
    END
  END w_mask_in[131]
  PIN w_mask_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.785 0.070 29.855 ;
    END
  END w_mask_in[132]
  PIN w_mask_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.995 0.070 30.065 ;
    END
  END w_mask_in[133]
  PIN w_mask_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.205 0.070 30.275 ;
    END
  END w_mask_in[134]
  PIN w_mask_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.415 0.070 30.485 ;
    END
  END w_mask_in[135]
  PIN w_mask_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.625 0.070 30.695 ;
    END
  END w_mask_in[136]
  PIN w_mask_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.835 0.070 30.905 ;
    END
  END w_mask_in[137]
  PIN w_mask_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.045 0.070 31.115 ;
    END
  END w_mask_in[138]
  PIN w_mask_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.255 0.070 31.325 ;
    END
  END w_mask_in[139]
  PIN w_mask_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.465 0.070 31.535 ;
    END
  END w_mask_in[140]
  PIN w_mask_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.675 0.070 31.745 ;
    END
  END w_mask_in[141]
  PIN w_mask_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.885 0.070 31.955 ;
    END
  END w_mask_in[142]
  PIN w_mask_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.095 0.070 32.165 ;
    END
  END w_mask_in[143]
  PIN w_mask_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.305 0.070 32.375 ;
    END
  END w_mask_in[144]
  PIN w_mask_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.515 0.070 32.585 ;
    END
  END w_mask_in[145]
  PIN w_mask_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END w_mask_in[146]
  PIN w_mask_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.935 0.070 33.005 ;
    END
  END w_mask_in[147]
  PIN w_mask_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.145 0.070 33.215 ;
    END
  END w_mask_in[148]
  PIN w_mask_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.355 0.070 33.425 ;
    END
  END w_mask_in[149]
  PIN w_mask_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END w_mask_in[150]
  PIN w_mask_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.775 0.070 33.845 ;
    END
  END w_mask_in[151]
  PIN w_mask_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.985 0.070 34.055 ;
    END
  END w_mask_in[152]
  PIN w_mask_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.195 0.070 34.265 ;
    END
  END w_mask_in[153]
  PIN w_mask_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END w_mask_in[154]
  PIN w_mask_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.615 0.070 34.685 ;
    END
  END w_mask_in[155]
  PIN w_mask_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.825 0.070 34.895 ;
    END
  END w_mask_in[156]
  PIN w_mask_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.035 0.070 35.105 ;
    END
  END w_mask_in[157]
  PIN w_mask_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END w_mask_in[158]
  PIN w_mask_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.455 0.070 35.525 ;
    END
  END w_mask_in[159]
  PIN w_mask_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END w_mask_in[160]
  PIN w_mask_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.875 0.070 35.945 ;
    END
  END w_mask_in[161]
  PIN w_mask_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END w_mask_in[162]
  PIN w_mask_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.295 0.070 36.365 ;
    END
  END w_mask_in[163]
  PIN w_mask_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.505 0.070 36.575 ;
    END
  END w_mask_in[164]
  PIN w_mask_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.715 0.070 36.785 ;
    END
  END w_mask_in[165]
  PIN w_mask_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END w_mask_in[166]
  PIN w_mask_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.135 0.070 37.205 ;
    END
  END w_mask_in[167]
  PIN w_mask_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END w_mask_in[168]
  PIN w_mask_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.555 0.070 37.625 ;
    END
  END w_mask_in[169]
  PIN w_mask_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END w_mask_in[170]
  PIN w_mask_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.975 0.070 38.045 ;
    END
  END w_mask_in[171]
  PIN w_mask_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.185 0.070 38.255 ;
    END
  END w_mask_in[172]
  PIN w_mask_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.395 0.070 38.465 ;
    END
  END w_mask_in[173]
  PIN w_mask_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END w_mask_in[174]
  PIN w_mask_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.815 0.070 38.885 ;
    END
  END w_mask_in[175]
  PIN w_mask_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END w_mask_in[176]
  PIN w_mask_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.235 0.070 39.305 ;
    END
  END w_mask_in[177]
  PIN w_mask_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END w_mask_in[178]
  PIN w_mask_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.655 0.070 39.725 ;
    END
  END w_mask_in[179]
  PIN w_mask_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END w_mask_in[180]
  PIN w_mask_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.075 0.070 40.145 ;
    END
  END w_mask_in[181]
  PIN w_mask_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END w_mask_in[182]
  PIN w_mask_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.495 0.070 40.565 ;
    END
  END w_mask_in[183]
  PIN w_mask_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END w_mask_in[184]
  PIN w_mask_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.915 0.070 40.985 ;
    END
  END w_mask_in[185]
  PIN w_mask_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END w_mask_in[186]
  PIN w_mask_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.335 0.070 41.405 ;
    END
  END w_mask_in[187]
  PIN w_mask_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END w_mask_in[188]
  PIN w_mask_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.755 0.070 41.825 ;
    END
  END w_mask_in[189]
  PIN w_mask_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END w_mask_in[190]
  PIN w_mask_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.175 0.070 42.245 ;
    END
  END w_mask_in[191]
  PIN w_mask_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END w_mask_in[192]
  PIN w_mask_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.595 0.070 42.665 ;
    END
  END w_mask_in[193]
  PIN w_mask_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END w_mask_in[194]
  PIN w_mask_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.015 0.070 43.085 ;
    END
  END w_mask_in[195]
  PIN w_mask_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END w_mask_in[196]
  PIN w_mask_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.435 0.070 43.505 ;
    END
  END w_mask_in[197]
  PIN w_mask_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END w_mask_in[198]
  PIN w_mask_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.855 0.070 43.925 ;
    END
  END w_mask_in[199]
  PIN w_mask_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END w_mask_in[200]
  PIN w_mask_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.275 0.070 44.345 ;
    END
  END w_mask_in[201]
  PIN w_mask_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END w_mask_in[202]
  PIN w_mask_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.695 0.070 44.765 ;
    END
  END w_mask_in[203]
  PIN w_mask_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END w_mask_in[204]
  PIN w_mask_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.115 0.070 45.185 ;
    END
  END w_mask_in[205]
  PIN w_mask_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.325 0.070 45.395 ;
    END
  END w_mask_in[206]
  PIN w_mask_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.535 0.070 45.605 ;
    END
  END w_mask_in[207]
  PIN w_mask_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.745 0.070 45.815 ;
    END
  END w_mask_in[208]
  PIN w_mask_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.955 0.070 46.025 ;
    END
  END w_mask_in[209]
  PIN w_mask_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END w_mask_in[210]
  PIN w_mask_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.375 0.070 46.445 ;
    END
  END w_mask_in[211]
  PIN w_mask_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.585 0.070 46.655 ;
    END
  END w_mask_in[212]
  PIN w_mask_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.795 0.070 46.865 ;
    END
  END w_mask_in[213]
  PIN w_mask_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END w_mask_in[214]
  PIN w_mask_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.215 0.070 47.285 ;
    END
  END w_mask_in[215]
  PIN w_mask_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END w_mask_in[216]
  PIN w_mask_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.635 0.070 47.705 ;
    END
  END w_mask_in[217]
  PIN w_mask_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END w_mask_in[218]
  PIN w_mask_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.055 0.070 48.125 ;
    END
  END w_mask_in[219]
  PIN w_mask_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.265 0.070 48.335 ;
    END
  END w_mask_in[220]
  PIN w_mask_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.475 0.070 48.545 ;
    END
  END w_mask_in[221]
  PIN w_mask_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END w_mask_in[222]
  PIN w_mask_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.895 0.070 48.965 ;
    END
  END w_mask_in[223]
  PIN w_mask_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END w_mask_in[224]
  PIN w_mask_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.315 0.070 49.385 ;
    END
  END w_mask_in[225]
  PIN w_mask_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END w_mask_in[226]
  PIN w_mask_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.735 0.070 49.805 ;
    END
  END w_mask_in[227]
  PIN w_mask_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.945 0.070 50.015 ;
    END
  END w_mask_in[228]
  PIN w_mask_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.155 0.070 50.225 ;
    END
  END w_mask_in[229]
  PIN w_mask_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END w_mask_in[230]
  PIN w_mask_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.575 0.070 50.645 ;
    END
  END w_mask_in[231]
  PIN w_mask_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.785 0.070 50.855 ;
    END
  END w_mask_in[232]
  PIN w_mask_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.995 0.070 51.065 ;
    END
  END w_mask_in[233]
  PIN w_mask_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.205 0.070 51.275 ;
    END
  END w_mask_in[234]
  PIN w_mask_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.415 0.070 51.485 ;
    END
  END w_mask_in[235]
  PIN w_mask_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.625 0.070 51.695 ;
    END
  END w_mask_in[236]
  PIN w_mask_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.835 0.070 51.905 ;
    END
  END w_mask_in[237]
  PIN w_mask_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.045 0.070 52.115 ;
    END
  END w_mask_in[238]
  PIN w_mask_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.255 0.070 52.325 ;
    END
  END w_mask_in[239]
  PIN w_mask_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END w_mask_in[240]
  PIN w_mask_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.675 0.070 52.745 ;
    END
  END w_mask_in[241]
  PIN w_mask_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END w_mask_in[242]
  PIN w_mask_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.095 0.070 53.165 ;
    END
  END w_mask_in[243]
  PIN w_mask_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.305 0.070 53.375 ;
    END
  END w_mask_in[244]
  PIN w_mask_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.515 0.070 53.585 ;
    END
  END w_mask_in[245]
  PIN w_mask_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END w_mask_in[246]
  PIN w_mask_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.935 0.070 54.005 ;
    END
  END w_mask_in[247]
  PIN w_mask_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.145 0.070 54.215 ;
    END
  END w_mask_in[248]
  PIN w_mask_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.355 0.070 54.425 ;
    END
  END w_mask_in[249]
  PIN w_mask_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END w_mask_in[250]
  PIN w_mask_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.775 0.070 54.845 ;
    END
  END w_mask_in[251]
  PIN w_mask_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.985 0.070 55.055 ;
    END
  END w_mask_in[252]
  PIN w_mask_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.195 0.070 55.265 ;
    END
  END w_mask_in[253]
  PIN w_mask_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END w_mask_in[254]
  PIN w_mask_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.615 0.070 55.685 ;
    END
  END w_mask_in[255]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.255 0.070 73.325 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.465 0.070 73.535 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.675 0.070 73.745 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.095 0.070 74.165 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.305 0.070 74.375 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.515 0.070 74.585 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.725 0.070 74.795 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.935 0.070 75.005 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.145 0.070 75.215 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.355 0.070 75.425 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.775 0.070 75.845 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.195 0.070 76.265 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.405 0.070 76.475 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.615 0.070 76.685 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.825 0.070 76.895 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.035 0.070 77.105 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.245 0.070 77.315 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.455 0.070 77.525 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.665 0.070 77.735 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.875 0.070 77.945 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.085 0.070 78.155 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.295 0.070 78.365 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.505 0.070 78.575 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.715 0.070 78.785 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.925 0.070 78.995 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.135 0.070 79.205 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.345 0.070 79.415 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.555 0.070 79.625 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.975 0.070 80.045 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.185 0.070 80.255 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.395 0.070 80.465 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.605 0.070 80.675 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.815 0.070 80.885 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.025 0.070 81.095 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.235 0.070 81.305 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.445 0.070 81.515 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.655 0.070 81.725 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.075 0.070 82.145 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.285 0.070 82.355 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.495 0.070 82.565 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.705 0.070 82.775 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.915 0.070 82.985 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.125 0.070 83.195 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.335 0.070 83.405 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.545 0.070 83.615 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.755 0.070 83.825 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.965 0.070 84.035 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.175 0.070 84.245 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.385 0.070 84.455 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.595 0.070 84.665 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.015 0.070 85.085 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.225 0.070 85.295 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.435 0.070 85.505 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.855 0.070 85.925 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.065 0.070 86.135 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.275 0.070 86.345 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.485 0.070 86.555 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.695 0.070 86.765 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.905 0.070 86.975 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.115 0.070 87.185 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.325 0.070 87.395 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.535 0.070 87.605 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.745 0.070 87.815 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.955 0.070 88.025 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.165 0.070 88.235 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.375 0.070 88.445 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.585 0.070 88.655 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.795 0.070 88.865 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.005 0.070 89.075 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.215 0.070 89.285 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.425 0.070 89.495 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.635 0.070 89.705 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.845 0.070 89.915 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.055 0.070 90.125 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.265 0.070 90.335 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.475 0.070 90.545 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.685 0.070 90.755 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.895 0.070 90.965 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.105 0.070 91.175 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.315 0.070 91.385 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.525 0.070 91.595 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.735 0.070 91.805 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.945 0.070 92.015 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.155 0.070 92.225 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.365 0.070 92.435 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.575 0.070 92.645 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.785 0.070 92.855 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.995 0.070 93.065 ;
    END
  END rd_out[95]
  PIN rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.205 0.070 93.275 ;
    END
  END rd_out[96]
  PIN rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.415 0.070 93.485 ;
    END
  END rd_out[97]
  PIN rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.625 0.070 93.695 ;
    END
  END rd_out[98]
  PIN rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.835 0.070 93.905 ;
    END
  END rd_out[99]
  PIN rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.045 0.070 94.115 ;
    END
  END rd_out[100]
  PIN rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.255 0.070 94.325 ;
    END
  END rd_out[101]
  PIN rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.465 0.070 94.535 ;
    END
  END rd_out[102]
  PIN rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.675 0.070 94.745 ;
    END
  END rd_out[103]
  PIN rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.885 0.070 94.955 ;
    END
  END rd_out[104]
  PIN rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.095 0.070 95.165 ;
    END
  END rd_out[105]
  PIN rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.305 0.070 95.375 ;
    END
  END rd_out[106]
  PIN rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.515 0.070 95.585 ;
    END
  END rd_out[107]
  PIN rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.725 0.070 95.795 ;
    END
  END rd_out[108]
  PIN rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.935 0.070 96.005 ;
    END
  END rd_out[109]
  PIN rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.145 0.070 96.215 ;
    END
  END rd_out[110]
  PIN rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.355 0.070 96.425 ;
    END
  END rd_out[111]
  PIN rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.565 0.070 96.635 ;
    END
  END rd_out[112]
  PIN rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.775 0.070 96.845 ;
    END
  END rd_out[113]
  PIN rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.985 0.070 97.055 ;
    END
  END rd_out[114]
  PIN rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.195 0.070 97.265 ;
    END
  END rd_out[115]
  PIN rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.405 0.070 97.475 ;
    END
  END rd_out[116]
  PIN rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.615 0.070 97.685 ;
    END
  END rd_out[117]
  PIN rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.825 0.070 97.895 ;
    END
  END rd_out[118]
  PIN rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.035 0.070 98.105 ;
    END
  END rd_out[119]
  PIN rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.245 0.070 98.315 ;
    END
  END rd_out[120]
  PIN rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.455 0.070 98.525 ;
    END
  END rd_out[121]
  PIN rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.665 0.070 98.735 ;
    END
  END rd_out[122]
  PIN rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.875 0.070 98.945 ;
    END
  END rd_out[123]
  PIN rd_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.085 0.070 99.155 ;
    END
  END rd_out[124]
  PIN rd_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.295 0.070 99.365 ;
    END
  END rd_out[125]
  PIN rd_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.505 0.070 99.575 ;
    END
  END rd_out[126]
  PIN rd_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.715 0.070 99.785 ;
    END
  END rd_out[127]
  PIN rd_out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.925 0.070 99.995 ;
    END
  END rd_out[128]
  PIN rd_out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.135 0.070 100.205 ;
    END
  END rd_out[129]
  PIN rd_out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.345 0.070 100.415 ;
    END
  END rd_out[130]
  PIN rd_out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.555 0.070 100.625 ;
    END
  END rd_out[131]
  PIN rd_out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.765 0.070 100.835 ;
    END
  END rd_out[132]
  PIN rd_out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.975 0.070 101.045 ;
    END
  END rd_out[133]
  PIN rd_out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.185 0.070 101.255 ;
    END
  END rd_out[134]
  PIN rd_out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.395 0.070 101.465 ;
    END
  END rd_out[135]
  PIN rd_out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.605 0.070 101.675 ;
    END
  END rd_out[136]
  PIN rd_out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.815 0.070 101.885 ;
    END
  END rd_out[137]
  PIN rd_out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.025 0.070 102.095 ;
    END
  END rd_out[138]
  PIN rd_out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.235 0.070 102.305 ;
    END
  END rd_out[139]
  PIN rd_out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.445 0.070 102.515 ;
    END
  END rd_out[140]
  PIN rd_out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.655 0.070 102.725 ;
    END
  END rd_out[141]
  PIN rd_out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.865 0.070 102.935 ;
    END
  END rd_out[142]
  PIN rd_out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.075 0.070 103.145 ;
    END
  END rd_out[143]
  PIN rd_out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.285 0.070 103.355 ;
    END
  END rd_out[144]
  PIN rd_out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.495 0.070 103.565 ;
    END
  END rd_out[145]
  PIN rd_out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.705 0.070 103.775 ;
    END
  END rd_out[146]
  PIN rd_out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.915 0.070 103.985 ;
    END
  END rd_out[147]
  PIN rd_out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.125 0.070 104.195 ;
    END
  END rd_out[148]
  PIN rd_out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.335 0.070 104.405 ;
    END
  END rd_out[149]
  PIN rd_out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.545 0.070 104.615 ;
    END
  END rd_out[150]
  PIN rd_out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.755 0.070 104.825 ;
    END
  END rd_out[151]
  PIN rd_out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.965 0.070 105.035 ;
    END
  END rd_out[152]
  PIN rd_out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.175 0.070 105.245 ;
    END
  END rd_out[153]
  PIN rd_out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.385 0.070 105.455 ;
    END
  END rd_out[154]
  PIN rd_out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.595 0.070 105.665 ;
    END
  END rd_out[155]
  PIN rd_out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.805 0.070 105.875 ;
    END
  END rd_out[156]
  PIN rd_out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.015 0.070 106.085 ;
    END
  END rd_out[157]
  PIN rd_out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.225 0.070 106.295 ;
    END
  END rd_out[158]
  PIN rd_out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.435 0.070 106.505 ;
    END
  END rd_out[159]
  PIN rd_out[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.645 0.070 106.715 ;
    END
  END rd_out[160]
  PIN rd_out[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.855 0.070 106.925 ;
    END
  END rd_out[161]
  PIN rd_out[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.065 0.070 107.135 ;
    END
  END rd_out[162]
  PIN rd_out[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.275 0.070 107.345 ;
    END
  END rd_out[163]
  PIN rd_out[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.485 0.070 107.555 ;
    END
  END rd_out[164]
  PIN rd_out[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.695 0.070 107.765 ;
    END
  END rd_out[165]
  PIN rd_out[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.905 0.070 107.975 ;
    END
  END rd_out[166]
  PIN rd_out[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.115 0.070 108.185 ;
    END
  END rd_out[167]
  PIN rd_out[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.325 0.070 108.395 ;
    END
  END rd_out[168]
  PIN rd_out[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.535 0.070 108.605 ;
    END
  END rd_out[169]
  PIN rd_out[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.745 0.070 108.815 ;
    END
  END rd_out[170]
  PIN rd_out[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.955 0.070 109.025 ;
    END
  END rd_out[171]
  PIN rd_out[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.165 0.070 109.235 ;
    END
  END rd_out[172]
  PIN rd_out[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.375 0.070 109.445 ;
    END
  END rd_out[173]
  PIN rd_out[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.585 0.070 109.655 ;
    END
  END rd_out[174]
  PIN rd_out[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.795 0.070 109.865 ;
    END
  END rd_out[175]
  PIN rd_out[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.005 0.070 110.075 ;
    END
  END rd_out[176]
  PIN rd_out[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.215 0.070 110.285 ;
    END
  END rd_out[177]
  PIN rd_out[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.425 0.070 110.495 ;
    END
  END rd_out[178]
  PIN rd_out[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.635 0.070 110.705 ;
    END
  END rd_out[179]
  PIN rd_out[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.845 0.070 110.915 ;
    END
  END rd_out[180]
  PIN rd_out[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.055 0.070 111.125 ;
    END
  END rd_out[181]
  PIN rd_out[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.265 0.070 111.335 ;
    END
  END rd_out[182]
  PIN rd_out[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.475 0.070 111.545 ;
    END
  END rd_out[183]
  PIN rd_out[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.685 0.070 111.755 ;
    END
  END rd_out[184]
  PIN rd_out[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.895 0.070 111.965 ;
    END
  END rd_out[185]
  PIN rd_out[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.105 0.070 112.175 ;
    END
  END rd_out[186]
  PIN rd_out[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.315 0.070 112.385 ;
    END
  END rd_out[187]
  PIN rd_out[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.525 0.070 112.595 ;
    END
  END rd_out[188]
  PIN rd_out[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.735 0.070 112.805 ;
    END
  END rd_out[189]
  PIN rd_out[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 112.945 0.070 113.015 ;
    END
  END rd_out[190]
  PIN rd_out[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.155 0.070 113.225 ;
    END
  END rd_out[191]
  PIN rd_out[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.365 0.070 113.435 ;
    END
  END rd_out[192]
  PIN rd_out[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.575 0.070 113.645 ;
    END
  END rd_out[193]
  PIN rd_out[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.785 0.070 113.855 ;
    END
  END rd_out[194]
  PIN rd_out[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.995 0.070 114.065 ;
    END
  END rd_out[195]
  PIN rd_out[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.205 0.070 114.275 ;
    END
  END rd_out[196]
  PIN rd_out[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.415 0.070 114.485 ;
    END
  END rd_out[197]
  PIN rd_out[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.625 0.070 114.695 ;
    END
  END rd_out[198]
  PIN rd_out[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.835 0.070 114.905 ;
    END
  END rd_out[199]
  PIN rd_out[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.045 0.070 115.115 ;
    END
  END rd_out[200]
  PIN rd_out[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.255 0.070 115.325 ;
    END
  END rd_out[201]
  PIN rd_out[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.465 0.070 115.535 ;
    END
  END rd_out[202]
  PIN rd_out[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.675 0.070 115.745 ;
    END
  END rd_out[203]
  PIN rd_out[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.885 0.070 115.955 ;
    END
  END rd_out[204]
  PIN rd_out[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.095 0.070 116.165 ;
    END
  END rd_out[205]
  PIN rd_out[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.305 0.070 116.375 ;
    END
  END rd_out[206]
  PIN rd_out[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.515 0.070 116.585 ;
    END
  END rd_out[207]
  PIN rd_out[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.725 0.070 116.795 ;
    END
  END rd_out[208]
  PIN rd_out[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.935 0.070 117.005 ;
    END
  END rd_out[209]
  PIN rd_out[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.145 0.070 117.215 ;
    END
  END rd_out[210]
  PIN rd_out[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.355 0.070 117.425 ;
    END
  END rd_out[211]
  PIN rd_out[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.565 0.070 117.635 ;
    END
  END rd_out[212]
  PIN rd_out[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.775 0.070 117.845 ;
    END
  END rd_out[213]
  PIN rd_out[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.985 0.070 118.055 ;
    END
  END rd_out[214]
  PIN rd_out[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.195 0.070 118.265 ;
    END
  END rd_out[215]
  PIN rd_out[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.405 0.070 118.475 ;
    END
  END rd_out[216]
  PIN rd_out[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.615 0.070 118.685 ;
    END
  END rd_out[217]
  PIN rd_out[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 118.825 0.070 118.895 ;
    END
  END rd_out[218]
  PIN rd_out[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.035 0.070 119.105 ;
    END
  END rd_out[219]
  PIN rd_out[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.245 0.070 119.315 ;
    END
  END rd_out[220]
  PIN rd_out[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.455 0.070 119.525 ;
    END
  END rd_out[221]
  PIN rd_out[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.665 0.070 119.735 ;
    END
  END rd_out[222]
  PIN rd_out[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.875 0.070 119.945 ;
    END
  END rd_out[223]
  PIN rd_out[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.085 0.070 120.155 ;
    END
  END rd_out[224]
  PIN rd_out[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.295 0.070 120.365 ;
    END
  END rd_out[225]
  PIN rd_out[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.505 0.070 120.575 ;
    END
  END rd_out[226]
  PIN rd_out[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.715 0.070 120.785 ;
    END
  END rd_out[227]
  PIN rd_out[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.925 0.070 120.995 ;
    END
  END rd_out[228]
  PIN rd_out[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.135 0.070 121.205 ;
    END
  END rd_out[229]
  PIN rd_out[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.345 0.070 121.415 ;
    END
  END rd_out[230]
  PIN rd_out[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.555 0.070 121.625 ;
    END
  END rd_out[231]
  PIN rd_out[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.765 0.070 121.835 ;
    END
  END rd_out[232]
  PIN rd_out[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.975 0.070 122.045 ;
    END
  END rd_out[233]
  PIN rd_out[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.185 0.070 122.255 ;
    END
  END rd_out[234]
  PIN rd_out[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.395 0.070 122.465 ;
    END
  END rd_out[235]
  PIN rd_out[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.605 0.070 122.675 ;
    END
  END rd_out[236]
  PIN rd_out[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 122.815 0.070 122.885 ;
    END
  END rd_out[237]
  PIN rd_out[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.025 0.070 123.095 ;
    END
  END rd_out[238]
  PIN rd_out[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.235 0.070 123.305 ;
    END
  END rd_out[239]
  PIN rd_out[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.445 0.070 123.515 ;
    END
  END rd_out[240]
  PIN rd_out[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.655 0.070 123.725 ;
    END
  END rd_out[241]
  PIN rd_out[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.865 0.070 123.935 ;
    END
  END rd_out[242]
  PIN rd_out[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.075 0.070 124.145 ;
    END
  END rd_out[243]
  PIN rd_out[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.285 0.070 124.355 ;
    END
  END rd_out[244]
  PIN rd_out[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.495 0.070 124.565 ;
    END
  END rd_out[245]
  PIN rd_out[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.705 0.070 124.775 ;
    END
  END rd_out[246]
  PIN rd_out[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.915 0.070 124.985 ;
    END
  END rd_out[247]
  PIN rd_out[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.125 0.070 125.195 ;
    END
  END rd_out[248]
  PIN rd_out[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.335 0.070 125.405 ;
    END
  END rd_out[249]
  PIN rd_out[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.545 0.070 125.615 ;
    END
  END rd_out[250]
  PIN rd_out[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.755 0.070 125.825 ;
    END
  END rd_out[251]
  PIN rd_out[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 125.965 0.070 126.035 ;
    END
  END rd_out[252]
  PIN rd_out[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.175 0.070 126.245 ;
    END
  END rd_out[253]
  PIN rd_out[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.385 0.070 126.455 ;
    END
  END rd_out[254]
  PIN rd_out[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.595 0.070 126.665 ;
    END
  END rd_out[255]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.025 0.070 144.095 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.235 0.070 144.305 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.445 0.070 144.515 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.655 0.070 144.725 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.865 0.070 144.935 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.075 0.070 145.145 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.285 0.070 145.355 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.495 0.070 145.565 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.705 0.070 145.775 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.915 0.070 145.985 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.125 0.070 146.195 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.335 0.070 146.405 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.545 0.070 146.615 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.755 0.070 146.825 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 146.965 0.070 147.035 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.175 0.070 147.245 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.385 0.070 147.455 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.595 0.070 147.665 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.805 0.070 147.875 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.015 0.070 148.085 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.225 0.070 148.295 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.435 0.070 148.505 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.645 0.070 148.715 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.855 0.070 148.925 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.065 0.070 149.135 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.275 0.070 149.345 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.485 0.070 149.555 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.695 0.070 149.765 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 149.905 0.070 149.975 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.115 0.070 150.185 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.325 0.070 150.395 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.535 0.070 150.605 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.745 0.070 150.815 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.955 0.070 151.025 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.165 0.070 151.235 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.375 0.070 151.445 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.585 0.070 151.655 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.795 0.070 151.865 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.005 0.070 152.075 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.215 0.070 152.285 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.425 0.070 152.495 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.635 0.070 152.705 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 152.845 0.070 152.915 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.055 0.070 153.125 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.265 0.070 153.335 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.475 0.070 153.545 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.685 0.070 153.755 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.895 0.070 153.965 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.105 0.070 154.175 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.315 0.070 154.385 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.525 0.070 154.595 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.735 0.070 154.805 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.945 0.070 155.015 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.155 0.070 155.225 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.365 0.070 155.435 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.575 0.070 155.645 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.785 0.070 155.855 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 155.995 0.070 156.065 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.205 0.070 156.275 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.415 0.070 156.485 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.625 0.070 156.695 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.835 0.070 156.905 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.045 0.070 157.115 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.255 0.070 157.325 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.465 0.070 157.535 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.675 0.070 157.745 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 157.885 0.070 157.955 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.095 0.070 158.165 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.305 0.070 158.375 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.515 0.070 158.585 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.725 0.070 158.795 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.935 0.070 159.005 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.145 0.070 159.215 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.355 0.070 159.425 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.565 0.070 159.635 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.775 0.070 159.845 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.985 0.070 160.055 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.195 0.070 160.265 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.405 0.070 160.475 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.615 0.070 160.685 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 160.825 0.070 160.895 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.035 0.070 161.105 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.245 0.070 161.315 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.455 0.070 161.525 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.665 0.070 161.735 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 161.875 0.070 161.945 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.085 0.070 162.155 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.295 0.070 162.365 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.505 0.070 162.575 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.715 0.070 162.785 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 162.925 0.070 162.995 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.135 0.070 163.205 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.345 0.070 163.415 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.555 0.070 163.625 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.765 0.070 163.835 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 163.975 0.070 164.045 ;
    END
  END wd_in[95]
  PIN wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.185 0.070 164.255 ;
    END
  END wd_in[96]
  PIN wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.395 0.070 164.465 ;
    END
  END wd_in[97]
  PIN wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.605 0.070 164.675 ;
    END
  END wd_in[98]
  PIN wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 164.815 0.070 164.885 ;
    END
  END wd_in[99]
  PIN wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.025 0.070 165.095 ;
    END
  END wd_in[100]
  PIN wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.235 0.070 165.305 ;
    END
  END wd_in[101]
  PIN wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.445 0.070 165.515 ;
    END
  END wd_in[102]
  PIN wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.655 0.070 165.725 ;
    END
  END wd_in[103]
  PIN wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 165.865 0.070 165.935 ;
    END
  END wd_in[104]
  PIN wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.075 0.070 166.145 ;
    END
  END wd_in[105]
  PIN wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.285 0.070 166.355 ;
    END
  END wd_in[106]
  PIN wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.495 0.070 166.565 ;
    END
  END wd_in[107]
  PIN wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.705 0.070 166.775 ;
    END
  END wd_in[108]
  PIN wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 166.915 0.070 166.985 ;
    END
  END wd_in[109]
  PIN wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.125 0.070 167.195 ;
    END
  END wd_in[110]
  PIN wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.335 0.070 167.405 ;
    END
  END wd_in[111]
  PIN wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.545 0.070 167.615 ;
    END
  END wd_in[112]
  PIN wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.755 0.070 167.825 ;
    END
  END wd_in[113]
  PIN wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 167.965 0.070 168.035 ;
    END
  END wd_in[114]
  PIN wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.175 0.070 168.245 ;
    END
  END wd_in[115]
  PIN wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.385 0.070 168.455 ;
    END
  END wd_in[116]
  PIN wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.595 0.070 168.665 ;
    END
  END wd_in[117]
  PIN wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 168.805 0.070 168.875 ;
    END
  END wd_in[118]
  PIN wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.015 0.070 169.085 ;
    END
  END wd_in[119]
  PIN wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.225 0.070 169.295 ;
    END
  END wd_in[120]
  PIN wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.435 0.070 169.505 ;
    END
  END wd_in[121]
  PIN wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.645 0.070 169.715 ;
    END
  END wd_in[122]
  PIN wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 169.855 0.070 169.925 ;
    END
  END wd_in[123]
  PIN wd_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.065 0.070 170.135 ;
    END
  END wd_in[124]
  PIN wd_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.275 0.070 170.345 ;
    END
  END wd_in[125]
  PIN wd_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.485 0.070 170.555 ;
    END
  END wd_in[126]
  PIN wd_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.695 0.070 170.765 ;
    END
  END wd_in[127]
  PIN wd_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 170.905 0.070 170.975 ;
    END
  END wd_in[128]
  PIN wd_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.115 0.070 171.185 ;
    END
  END wd_in[129]
  PIN wd_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.325 0.070 171.395 ;
    END
  END wd_in[130]
  PIN wd_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.535 0.070 171.605 ;
    END
  END wd_in[131]
  PIN wd_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.745 0.070 171.815 ;
    END
  END wd_in[132]
  PIN wd_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 171.955 0.070 172.025 ;
    END
  END wd_in[133]
  PIN wd_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.165 0.070 172.235 ;
    END
  END wd_in[134]
  PIN wd_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.375 0.070 172.445 ;
    END
  END wd_in[135]
  PIN wd_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.585 0.070 172.655 ;
    END
  END wd_in[136]
  PIN wd_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 172.795 0.070 172.865 ;
    END
  END wd_in[137]
  PIN wd_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.005 0.070 173.075 ;
    END
  END wd_in[138]
  PIN wd_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.215 0.070 173.285 ;
    END
  END wd_in[139]
  PIN wd_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.425 0.070 173.495 ;
    END
  END wd_in[140]
  PIN wd_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.635 0.070 173.705 ;
    END
  END wd_in[141]
  PIN wd_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 173.845 0.070 173.915 ;
    END
  END wd_in[142]
  PIN wd_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.055 0.070 174.125 ;
    END
  END wd_in[143]
  PIN wd_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.265 0.070 174.335 ;
    END
  END wd_in[144]
  PIN wd_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.475 0.070 174.545 ;
    END
  END wd_in[145]
  PIN wd_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.685 0.070 174.755 ;
    END
  END wd_in[146]
  PIN wd_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 174.895 0.070 174.965 ;
    END
  END wd_in[147]
  PIN wd_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.105 0.070 175.175 ;
    END
  END wd_in[148]
  PIN wd_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.315 0.070 175.385 ;
    END
  END wd_in[149]
  PIN wd_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.525 0.070 175.595 ;
    END
  END wd_in[150]
  PIN wd_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.735 0.070 175.805 ;
    END
  END wd_in[151]
  PIN wd_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 175.945 0.070 176.015 ;
    END
  END wd_in[152]
  PIN wd_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.155 0.070 176.225 ;
    END
  END wd_in[153]
  PIN wd_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.365 0.070 176.435 ;
    END
  END wd_in[154]
  PIN wd_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.575 0.070 176.645 ;
    END
  END wd_in[155]
  PIN wd_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.785 0.070 176.855 ;
    END
  END wd_in[156]
  PIN wd_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 176.995 0.070 177.065 ;
    END
  END wd_in[157]
  PIN wd_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.205 0.070 177.275 ;
    END
  END wd_in[158]
  PIN wd_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.415 0.070 177.485 ;
    END
  END wd_in[159]
  PIN wd_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.625 0.070 177.695 ;
    END
  END wd_in[160]
  PIN wd_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 177.835 0.070 177.905 ;
    END
  END wd_in[161]
  PIN wd_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.045 0.070 178.115 ;
    END
  END wd_in[162]
  PIN wd_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.255 0.070 178.325 ;
    END
  END wd_in[163]
  PIN wd_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.465 0.070 178.535 ;
    END
  END wd_in[164]
  PIN wd_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.675 0.070 178.745 ;
    END
  END wd_in[165]
  PIN wd_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 178.885 0.070 178.955 ;
    END
  END wd_in[166]
  PIN wd_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.095 0.070 179.165 ;
    END
  END wd_in[167]
  PIN wd_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.305 0.070 179.375 ;
    END
  END wd_in[168]
  PIN wd_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.515 0.070 179.585 ;
    END
  END wd_in[169]
  PIN wd_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.725 0.070 179.795 ;
    END
  END wd_in[170]
  PIN wd_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 179.935 0.070 180.005 ;
    END
  END wd_in[171]
  PIN wd_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.145 0.070 180.215 ;
    END
  END wd_in[172]
  PIN wd_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.355 0.070 180.425 ;
    END
  END wd_in[173]
  PIN wd_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.565 0.070 180.635 ;
    END
  END wd_in[174]
  PIN wd_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.775 0.070 180.845 ;
    END
  END wd_in[175]
  PIN wd_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 180.985 0.070 181.055 ;
    END
  END wd_in[176]
  PIN wd_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.195 0.070 181.265 ;
    END
  END wd_in[177]
  PIN wd_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.405 0.070 181.475 ;
    END
  END wd_in[178]
  PIN wd_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.615 0.070 181.685 ;
    END
  END wd_in[179]
  PIN wd_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 181.825 0.070 181.895 ;
    END
  END wd_in[180]
  PIN wd_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.035 0.070 182.105 ;
    END
  END wd_in[181]
  PIN wd_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.245 0.070 182.315 ;
    END
  END wd_in[182]
  PIN wd_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.455 0.070 182.525 ;
    END
  END wd_in[183]
  PIN wd_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.665 0.070 182.735 ;
    END
  END wd_in[184]
  PIN wd_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 182.875 0.070 182.945 ;
    END
  END wd_in[185]
  PIN wd_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.085 0.070 183.155 ;
    END
  END wd_in[186]
  PIN wd_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.295 0.070 183.365 ;
    END
  END wd_in[187]
  PIN wd_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.505 0.070 183.575 ;
    END
  END wd_in[188]
  PIN wd_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.715 0.070 183.785 ;
    END
  END wd_in[189]
  PIN wd_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 183.925 0.070 183.995 ;
    END
  END wd_in[190]
  PIN wd_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.135 0.070 184.205 ;
    END
  END wd_in[191]
  PIN wd_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.345 0.070 184.415 ;
    END
  END wd_in[192]
  PIN wd_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.555 0.070 184.625 ;
    END
  END wd_in[193]
  PIN wd_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.765 0.070 184.835 ;
    END
  END wd_in[194]
  PIN wd_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 184.975 0.070 185.045 ;
    END
  END wd_in[195]
  PIN wd_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.185 0.070 185.255 ;
    END
  END wd_in[196]
  PIN wd_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.395 0.070 185.465 ;
    END
  END wd_in[197]
  PIN wd_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.605 0.070 185.675 ;
    END
  END wd_in[198]
  PIN wd_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 185.815 0.070 185.885 ;
    END
  END wd_in[199]
  PIN wd_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.025 0.070 186.095 ;
    END
  END wd_in[200]
  PIN wd_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.235 0.070 186.305 ;
    END
  END wd_in[201]
  PIN wd_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.445 0.070 186.515 ;
    END
  END wd_in[202]
  PIN wd_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.655 0.070 186.725 ;
    END
  END wd_in[203]
  PIN wd_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 186.865 0.070 186.935 ;
    END
  END wd_in[204]
  PIN wd_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.075 0.070 187.145 ;
    END
  END wd_in[205]
  PIN wd_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.285 0.070 187.355 ;
    END
  END wd_in[206]
  PIN wd_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.495 0.070 187.565 ;
    END
  END wd_in[207]
  PIN wd_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.705 0.070 187.775 ;
    END
  END wd_in[208]
  PIN wd_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 187.915 0.070 187.985 ;
    END
  END wd_in[209]
  PIN wd_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.125 0.070 188.195 ;
    END
  END wd_in[210]
  PIN wd_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.335 0.070 188.405 ;
    END
  END wd_in[211]
  PIN wd_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.545 0.070 188.615 ;
    END
  END wd_in[212]
  PIN wd_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.755 0.070 188.825 ;
    END
  END wd_in[213]
  PIN wd_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 188.965 0.070 189.035 ;
    END
  END wd_in[214]
  PIN wd_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.175 0.070 189.245 ;
    END
  END wd_in[215]
  PIN wd_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.385 0.070 189.455 ;
    END
  END wd_in[216]
  PIN wd_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.595 0.070 189.665 ;
    END
  END wd_in[217]
  PIN wd_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 189.805 0.070 189.875 ;
    END
  END wd_in[218]
  PIN wd_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.015 0.070 190.085 ;
    END
  END wd_in[219]
  PIN wd_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.225 0.070 190.295 ;
    END
  END wd_in[220]
  PIN wd_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.435 0.070 190.505 ;
    END
  END wd_in[221]
  PIN wd_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.645 0.070 190.715 ;
    END
  END wd_in[222]
  PIN wd_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 190.855 0.070 190.925 ;
    END
  END wd_in[223]
  PIN wd_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.065 0.070 191.135 ;
    END
  END wd_in[224]
  PIN wd_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.275 0.070 191.345 ;
    END
  END wd_in[225]
  PIN wd_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.485 0.070 191.555 ;
    END
  END wd_in[226]
  PIN wd_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.695 0.070 191.765 ;
    END
  END wd_in[227]
  PIN wd_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 191.905 0.070 191.975 ;
    END
  END wd_in[228]
  PIN wd_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.115 0.070 192.185 ;
    END
  END wd_in[229]
  PIN wd_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.325 0.070 192.395 ;
    END
  END wd_in[230]
  PIN wd_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.535 0.070 192.605 ;
    END
  END wd_in[231]
  PIN wd_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.745 0.070 192.815 ;
    END
  END wd_in[232]
  PIN wd_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 192.955 0.070 193.025 ;
    END
  END wd_in[233]
  PIN wd_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.165 0.070 193.235 ;
    END
  END wd_in[234]
  PIN wd_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.375 0.070 193.445 ;
    END
  END wd_in[235]
  PIN wd_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.585 0.070 193.655 ;
    END
  END wd_in[236]
  PIN wd_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 193.795 0.070 193.865 ;
    END
  END wd_in[237]
  PIN wd_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.005 0.070 194.075 ;
    END
  END wd_in[238]
  PIN wd_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.215 0.070 194.285 ;
    END
  END wd_in[239]
  PIN wd_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.425 0.070 194.495 ;
    END
  END wd_in[240]
  PIN wd_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.635 0.070 194.705 ;
    END
  END wd_in[241]
  PIN wd_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 194.845 0.070 194.915 ;
    END
  END wd_in[242]
  PIN wd_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.055 0.070 195.125 ;
    END
  END wd_in[243]
  PIN wd_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.265 0.070 195.335 ;
    END
  END wd_in[244]
  PIN wd_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.475 0.070 195.545 ;
    END
  END wd_in[245]
  PIN wd_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.685 0.070 195.755 ;
    END
  END wd_in[246]
  PIN wd_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 195.895 0.070 195.965 ;
    END
  END wd_in[247]
  PIN wd_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.105 0.070 196.175 ;
    END
  END wd_in[248]
  PIN wd_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.315 0.070 196.385 ;
    END
  END wd_in[249]
  PIN wd_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.525 0.070 196.595 ;
    END
  END wd_in[250]
  PIN wd_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.735 0.070 196.805 ;
    END
  END wd_in[251]
  PIN wd_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 196.945 0.070 197.015 ;
    END
  END wd_in[252]
  PIN wd_in[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.155 0.070 197.225 ;
    END
  END wd_in[253]
  PIN wd_in[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.365 0.070 197.435 ;
    END
  END wd_in[254]
  PIN wd_in[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 197.575 0.070 197.645 ;
    END
  END wd_in[255]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.005 0.070 215.075 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.215 0.070 215.285 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.425 0.070 215.495 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.635 0.070 215.705 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 215.845 0.070 215.915 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.055 0.070 216.125 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 216.265 0.070 216.335 ;
    END
  END addr_in[6]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 233.695 0.070 233.765 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 233.905 0.070 233.975 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 234.115 0.070 234.185 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 235.900 ;
      RECT 5.320 2.100 5.600 235.900 ;
      RECT 8.680 2.100 8.960 235.900 ;
      RECT 12.040 2.100 12.320 235.900 ;
      RECT 15.400 2.100 15.680 235.900 ;
      RECT 18.760 2.100 19.040 235.900 ;
      RECT 22.120 2.100 22.400 235.900 ;
      RECT 25.480 2.100 25.760 235.900 ;
      RECT 28.840 2.100 29.120 235.900 ;
      RECT 32.200 2.100 32.480 235.900 ;
      RECT 35.560 2.100 35.840 235.900 ;
      RECT 38.920 2.100 39.200 235.900 ;
      RECT 42.280 2.100 42.560 235.900 ;
      RECT 45.640 2.100 45.920 235.900 ;
      RECT 49.000 2.100 49.280 235.900 ;
      RECT 52.360 2.100 52.640 235.900 ;
      RECT 55.720 2.100 56.000 235.900 ;
      RECT 59.080 2.100 59.360 235.900 ;
      RECT 62.440 2.100 62.720 235.900 ;
      RECT 65.800 2.100 66.080 235.900 ;
      RECT 69.160 2.100 69.440 235.900 ;
      RECT 72.520 2.100 72.800 235.900 ;
      RECT 75.880 2.100 76.160 235.900 ;
      RECT 79.240 2.100 79.520 235.900 ;
      RECT 82.600 2.100 82.880 235.900 ;
      RECT 85.960 2.100 86.240 235.900 ;
      RECT 89.320 2.100 89.600 235.900 ;
      RECT 92.680 2.100 92.960 235.900 ;
      RECT 96.040 2.100 96.320 235.900 ;
      RECT 99.400 2.100 99.680 235.900 ;
      RECT 102.760 2.100 103.040 235.900 ;
      RECT 106.120 2.100 106.400 235.900 ;
      RECT 109.480 2.100 109.760 235.900 ;
      RECT 112.840 2.100 113.120 235.900 ;
      RECT 116.200 2.100 116.480 235.900 ;
      RECT 119.560 2.100 119.840 235.900 ;
      RECT 122.920 2.100 123.200 235.900 ;
      RECT 126.280 2.100 126.560 235.900 ;
      RECT 129.640 2.100 129.920 235.900 ;
      RECT 133.000 2.100 133.280 235.900 ;
      RECT 136.360 2.100 136.640 235.900 ;
      RECT 139.720 2.100 140.000 235.900 ;
      RECT 143.080 2.100 143.360 235.900 ;
      RECT 146.440 2.100 146.720 235.900 ;
      RECT 149.800 2.100 150.080 235.900 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 235.900 ;
      RECT 7.000 2.100 7.280 235.900 ;
      RECT 10.360 2.100 10.640 235.900 ;
      RECT 13.720 2.100 14.000 235.900 ;
      RECT 17.080 2.100 17.360 235.900 ;
      RECT 20.440 2.100 20.720 235.900 ;
      RECT 23.800 2.100 24.080 235.900 ;
      RECT 27.160 2.100 27.440 235.900 ;
      RECT 30.520 2.100 30.800 235.900 ;
      RECT 33.880 2.100 34.160 235.900 ;
      RECT 37.240 2.100 37.520 235.900 ;
      RECT 40.600 2.100 40.880 235.900 ;
      RECT 43.960 2.100 44.240 235.900 ;
      RECT 47.320 2.100 47.600 235.900 ;
      RECT 50.680 2.100 50.960 235.900 ;
      RECT 54.040 2.100 54.320 235.900 ;
      RECT 57.400 2.100 57.680 235.900 ;
      RECT 60.760 2.100 61.040 235.900 ;
      RECT 64.120 2.100 64.400 235.900 ;
      RECT 67.480 2.100 67.760 235.900 ;
      RECT 70.840 2.100 71.120 235.900 ;
      RECT 74.200 2.100 74.480 235.900 ;
      RECT 77.560 2.100 77.840 235.900 ;
      RECT 80.920 2.100 81.200 235.900 ;
      RECT 84.280 2.100 84.560 235.900 ;
      RECT 87.640 2.100 87.920 235.900 ;
      RECT 91.000 2.100 91.280 235.900 ;
      RECT 94.360 2.100 94.640 235.900 ;
      RECT 97.720 2.100 98.000 235.900 ;
      RECT 101.080 2.100 101.360 235.900 ;
      RECT 104.440 2.100 104.720 235.900 ;
      RECT 107.800 2.100 108.080 235.900 ;
      RECT 111.160 2.100 111.440 235.900 ;
      RECT 114.520 2.100 114.800 235.900 ;
      RECT 117.880 2.100 118.160 235.900 ;
      RECT 121.240 2.100 121.520 235.900 ;
      RECT 124.600 2.100 124.880 235.900 ;
      RECT 127.960 2.100 128.240 235.900 ;
      RECT 131.320 2.100 131.600 235.900 ;
      RECT 134.680 2.100 134.960 235.900 ;
      RECT 138.040 2.100 138.320 235.900 ;
      RECT 141.400 2.100 141.680 235.900 ;
      RECT 144.760 2.100 145.040 235.900 ;
      RECT 148.120 2.100 148.400 235.900 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 153.710 238.000 ;
    LAYER metal2 ;
    RECT 0 0 153.710 238.000 ;
    LAYER metal3 ;
    RECT 0.070 0 153.710 238.000 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.275 ;
    RECT 0 2.345 0.070 2.485 ;
    RECT 0 2.555 0.070 2.695 ;
    RECT 0 2.765 0.070 2.905 ;
    RECT 0 2.975 0.070 3.115 ;
    RECT 0 3.185 0.070 3.325 ;
    RECT 0 3.395 0.070 3.535 ;
    RECT 0 3.605 0.070 3.745 ;
    RECT 0 3.815 0.070 3.955 ;
    RECT 0 4.025 0.070 4.165 ;
    RECT 0 4.235 0.070 4.375 ;
    RECT 0 4.445 0.070 4.585 ;
    RECT 0 4.655 0.070 4.795 ;
    RECT 0 4.865 0.070 5.005 ;
    RECT 0 5.075 0.070 5.215 ;
    RECT 0 5.285 0.070 5.425 ;
    RECT 0 5.495 0.070 5.635 ;
    RECT 0 5.705 0.070 5.845 ;
    RECT 0 5.915 0.070 6.055 ;
    RECT 0 6.125 0.070 6.265 ;
    RECT 0 6.335 0.070 6.475 ;
    RECT 0 6.545 0.070 6.685 ;
    RECT 0 6.755 0.070 6.895 ;
    RECT 0 6.965 0.070 7.105 ;
    RECT 0 7.175 0.070 7.315 ;
    RECT 0 7.385 0.070 7.525 ;
    RECT 0 7.595 0.070 7.735 ;
    RECT 0 7.805 0.070 7.945 ;
    RECT 0 8.015 0.070 8.155 ;
    RECT 0 8.225 0.070 8.365 ;
    RECT 0 8.435 0.070 8.575 ;
    RECT 0 8.645 0.070 8.785 ;
    RECT 0 8.855 0.070 8.995 ;
    RECT 0 9.065 0.070 9.205 ;
    RECT 0 9.275 0.070 9.415 ;
    RECT 0 9.485 0.070 9.625 ;
    RECT 0 9.695 0.070 9.835 ;
    RECT 0 9.905 0.070 10.045 ;
    RECT 0 10.115 0.070 10.255 ;
    RECT 0 10.325 0.070 10.465 ;
    RECT 0 10.535 0.070 10.675 ;
    RECT 0 10.745 0.070 10.885 ;
    RECT 0 10.955 0.070 11.095 ;
    RECT 0 11.165 0.070 11.305 ;
    RECT 0 11.375 0.070 11.515 ;
    RECT 0 11.585 0.070 11.725 ;
    RECT 0 11.795 0.070 11.935 ;
    RECT 0 12.005 0.070 12.145 ;
    RECT 0 12.215 0.070 12.355 ;
    RECT 0 12.425 0.070 12.565 ;
    RECT 0 12.635 0.070 12.775 ;
    RECT 0 12.845 0.070 12.985 ;
    RECT 0 13.055 0.070 13.195 ;
    RECT 0 13.265 0.070 13.405 ;
    RECT 0 13.475 0.070 13.615 ;
    RECT 0 13.685 0.070 13.825 ;
    RECT 0 13.895 0.070 14.035 ;
    RECT 0 14.105 0.070 14.245 ;
    RECT 0 14.315 0.070 14.455 ;
    RECT 0 14.525 0.070 14.665 ;
    RECT 0 14.735 0.070 14.875 ;
    RECT 0 14.945 0.070 15.085 ;
    RECT 0 15.155 0.070 15.295 ;
    RECT 0 15.365 0.070 15.505 ;
    RECT 0 15.575 0.070 15.715 ;
    RECT 0 15.785 0.070 15.925 ;
    RECT 0 15.995 0.070 16.135 ;
    RECT 0 16.205 0.070 16.345 ;
    RECT 0 16.415 0.070 16.555 ;
    RECT 0 16.625 0.070 16.765 ;
    RECT 0 16.835 0.070 16.975 ;
    RECT 0 17.045 0.070 17.185 ;
    RECT 0 17.255 0.070 17.395 ;
    RECT 0 17.465 0.070 17.605 ;
    RECT 0 17.675 0.070 17.815 ;
    RECT 0 17.885 0.070 18.025 ;
    RECT 0 18.095 0.070 18.235 ;
    RECT 0 18.305 0.070 18.445 ;
    RECT 0 18.515 0.070 18.655 ;
    RECT 0 18.725 0.070 18.865 ;
    RECT 0 18.935 0.070 19.075 ;
    RECT 0 19.145 0.070 19.285 ;
    RECT 0 19.355 0.070 19.495 ;
    RECT 0 19.565 0.070 19.705 ;
    RECT 0 19.775 0.070 19.915 ;
    RECT 0 19.985 0.070 20.125 ;
    RECT 0 20.195 0.070 20.335 ;
    RECT 0 20.405 0.070 20.545 ;
    RECT 0 20.615 0.070 20.755 ;
    RECT 0 20.825 0.070 20.965 ;
    RECT 0 21.035 0.070 21.175 ;
    RECT 0 21.245 0.070 21.385 ;
    RECT 0 21.455 0.070 21.595 ;
    RECT 0 21.665 0.070 21.805 ;
    RECT 0 21.875 0.070 22.015 ;
    RECT 0 22.085 0.070 22.225 ;
    RECT 0 22.295 0.070 22.435 ;
    RECT 0 22.505 0.070 22.645 ;
    RECT 0 22.715 0.070 22.855 ;
    RECT 0 22.925 0.070 23.065 ;
    RECT 0 23.135 0.070 23.275 ;
    RECT 0 23.345 0.070 23.485 ;
    RECT 0 23.555 0.070 23.695 ;
    RECT 0 23.765 0.070 23.905 ;
    RECT 0 23.975 0.070 24.115 ;
    RECT 0 24.185 0.070 24.325 ;
    RECT 0 24.395 0.070 24.535 ;
    RECT 0 24.605 0.070 24.745 ;
    RECT 0 24.815 0.070 24.955 ;
    RECT 0 25.025 0.070 25.165 ;
    RECT 0 25.235 0.070 25.375 ;
    RECT 0 25.445 0.070 25.585 ;
    RECT 0 25.655 0.070 25.795 ;
    RECT 0 25.865 0.070 26.005 ;
    RECT 0 26.075 0.070 26.215 ;
    RECT 0 26.285 0.070 26.425 ;
    RECT 0 26.495 0.070 26.635 ;
    RECT 0 26.705 0.070 26.845 ;
    RECT 0 26.915 0.070 27.055 ;
    RECT 0 27.125 0.070 27.265 ;
    RECT 0 27.335 0.070 27.475 ;
    RECT 0 27.545 0.070 27.685 ;
    RECT 0 27.755 0.070 27.895 ;
    RECT 0 27.965 0.070 28.105 ;
    RECT 0 28.175 0.070 28.315 ;
    RECT 0 28.385 0.070 28.525 ;
    RECT 0 28.595 0.070 28.735 ;
    RECT 0 28.805 0.070 28.945 ;
    RECT 0 29.015 0.070 29.155 ;
    RECT 0 29.225 0.070 29.365 ;
    RECT 0 29.435 0.070 29.575 ;
    RECT 0 29.645 0.070 29.785 ;
    RECT 0 29.855 0.070 29.995 ;
    RECT 0 30.065 0.070 30.205 ;
    RECT 0 30.275 0.070 30.415 ;
    RECT 0 30.485 0.070 30.625 ;
    RECT 0 30.695 0.070 30.835 ;
    RECT 0 30.905 0.070 31.045 ;
    RECT 0 31.115 0.070 31.255 ;
    RECT 0 31.325 0.070 31.465 ;
    RECT 0 31.535 0.070 31.675 ;
    RECT 0 31.745 0.070 31.885 ;
    RECT 0 31.955 0.070 32.095 ;
    RECT 0 32.165 0.070 32.305 ;
    RECT 0 32.375 0.070 32.515 ;
    RECT 0 32.585 0.070 32.725 ;
    RECT 0 32.795 0.070 32.935 ;
    RECT 0 33.005 0.070 33.145 ;
    RECT 0 33.215 0.070 33.355 ;
    RECT 0 33.425 0.070 33.565 ;
    RECT 0 33.635 0.070 33.775 ;
    RECT 0 33.845 0.070 33.985 ;
    RECT 0 34.055 0.070 34.195 ;
    RECT 0 34.265 0.070 34.405 ;
    RECT 0 34.475 0.070 34.615 ;
    RECT 0 34.685 0.070 34.825 ;
    RECT 0 34.895 0.070 35.035 ;
    RECT 0 35.105 0.070 35.245 ;
    RECT 0 35.315 0.070 35.455 ;
    RECT 0 35.525 0.070 35.665 ;
    RECT 0 35.735 0.070 35.875 ;
    RECT 0 35.945 0.070 36.085 ;
    RECT 0 36.155 0.070 36.295 ;
    RECT 0 36.365 0.070 36.505 ;
    RECT 0 36.575 0.070 36.715 ;
    RECT 0 36.785 0.070 36.925 ;
    RECT 0 36.995 0.070 37.135 ;
    RECT 0 37.205 0.070 37.345 ;
    RECT 0 37.415 0.070 37.555 ;
    RECT 0 37.625 0.070 37.765 ;
    RECT 0 37.835 0.070 37.975 ;
    RECT 0 38.045 0.070 38.185 ;
    RECT 0 38.255 0.070 38.395 ;
    RECT 0 38.465 0.070 38.605 ;
    RECT 0 38.675 0.070 38.815 ;
    RECT 0 38.885 0.070 39.025 ;
    RECT 0 39.095 0.070 39.235 ;
    RECT 0 39.305 0.070 39.445 ;
    RECT 0 39.515 0.070 39.655 ;
    RECT 0 39.725 0.070 39.865 ;
    RECT 0 39.935 0.070 40.075 ;
    RECT 0 40.145 0.070 40.285 ;
    RECT 0 40.355 0.070 40.495 ;
    RECT 0 40.565 0.070 40.705 ;
    RECT 0 40.775 0.070 40.915 ;
    RECT 0 40.985 0.070 41.125 ;
    RECT 0 41.195 0.070 41.335 ;
    RECT 0 41.405 0.070 41.545 ;
    RECT 0 41.615 0.070 41.755 ;
    RECT 0 41.825 0.070 41.965 ;
    RECT 0 42.035 0.070 42.175 ;
    RECT 0 42.245 0.070 42.385 ;
    RECT 0 42.455 0.070 42.595 ;
    RECT 0 42.665 0.070 42.805 ;
    RECT 0 42.875 0.070 43.015 ;
    RECT 0 43.085 0.070 43.225 ;
    RECT 0 43.295 0.070 43.435 ;
    RECT 0 43.505 0.070 43.645 ;
    RECT 0 43.715 0.070 43.855 ;
    RECT 0 43.925 0.070 44.065 ;
    RECT 0 44.135 0.070 44.275 ;
    RECT 0 44.345 0.070 44.485 ;
    RECT 0 44.555 0.070 44.695 ;
    RECT 0 44.765 0.070 44.905 ;
    RECT 0 44.975 0.070 45.115 ;
    RECT 0 45.185 0.070 45.325 ;
    RECT 0 45.395 0.070 45.535 ;
    RECT 0 45.605 0.070 45.745 ;
    RECT 0 45.815 0.070 45.955 ;
    RECT 0 46.025 0.070 46.165 ;
    RECT 0 46.235 0.070 46.375 ;
    RECT 0 46.445 0.070 46.585 ;
    RECT 0 46.655 0.070 46.795 ;
    RECT 0 46.865 0.070 47.005 ;
    RECT 0 47.075 0.070 47.215 ;
    RECT 0 47.285 0.070 47.425 ;
    RECT 0 47.495 0.070 47.635 ;
    RECT 0 47.705 0.070 47.845 ;
    RECT 0 47.915 0.070 48.055 ;
    RECT 0 48.125 0.070 48.265 ;
    RECT 0 48.335 0.070 48.475 ;
    RECT 0 48.545 0.070 48.685 ;
    RECT 0 48.755 0.070 48.895 ;
    RECT 0 48.965 0.070 49.105 ;
    RECT 0 49.175 0.070 49.315 ;
    RECT 0 49.385 0.070 49.525 ;
    RECT 0 49.595 0.070 49.735 ;
    RECT 0 49.805 0.070 49.945 ;
    RECT 0 50.015 0.070 50.155 ;
    RECT 0 50.225 0.070 50.365 ;
    RECT 0 50.435 0.070 50.575 ;
    RECT 0 50.645 0.070 50.785 ;
    RECT 0 50.855 0.070 50.995 ;
    RECT 0 51.065 0.070 51.205 ;
    RECT 0 51.275 0.070 51.415 ;
    RECT 0 51.485 0.070 51.625 ;
    RECT 0 51.695 0.070 51.835 ;
    RECT 0 51.905 0.070 52.045 ;
    RECT 0 52.115 0.070 52.255 ;
    RECT 0 52.325 0.070 52.465 ;
    RECT 0 52.535 0.070 52.675 ;
    RECT 0 52.745 0.070 52.885 ;
    RECT 0 52.955 0.070 53.095 ;
    RECT 0 53.165 0.070 53.305 ;
    RECT 0 53.375 0.070 53.515 ;
    RECT 0 53.585 0.070 53.725 ;
    RECT 0 53.795 0.070 53.935 ;
    RECT 0 54.005 0.070 54.145 ;
    RECT 0 54.215 0.070 54.355 ;
    RECT 0 54.425 0.070 54.565 ;
    RECT 0 54.635 0.070 54.775 ;
    RECT 0 54.845 0.070 54.985 ;
    RECT 0 55.055 0.070 55.195 ;
    RECT 0 55.265 0.070 55.405 ;
    RECT 0 55.475 0.070 55.615 ;
    RECT 0 55.685 0.070 73.045 ;
    RECT 0 73.115 0.070 73.255 ;
    RECT 0 73.325 0.070 73.465 ;
    RECT 0 73.535 0.070 73.675 ;
    RECT 0 73.745 0.070 73.885 ;
    RECT 0 73.955 0.070 74.095 ;
    RECT 0 74.165 0.070 74.305 ;
    RECT 0 74.375 0.070 74.515 ;
    RECT 0 74.585 0.070 74.725 ;
    RECT 0 74.795 0.070 74.935 ;
    RECT 0 75.005 0.070 75.145 ;
    RECT 0 75.215 0.070 75.355 ;
    RECT 0 75.425 0.070 75.565 ;
    RECT 0 75.635 0.070 75.775 ;
    RECT 0 75.845 0.070 75.985 ;
    RECT 0 76.055 0.070 76.195 ;
    RECT 0 76.265 0.070 76.405 ;
    RECT 0 76.475 0.070 76.615 ;
    RECT 0 76.685 0.070 76.825 ;
    RECT 0 76.895 0.070 77.035 ;
    RECT 0 77.105 0.070 77.245 ;
    RECT 0 77.315 0.070 77.455 ;
    RECT 0 77.525 0.070 77.665 ;
    RECT 0 77.735 0.070 77.875 ;
    RECT 0 77.945 0.070 78.085 ;
    RECT 0 78.155 0.070 78.295 ;
    RECT 0 78.365 0.070 78.505 ;
    RECT 0 78.575 0.070 78.715 ;
    RECT 0 78.785 0.070 78.925 ;
    RECT 0 78.995 0.070 79.135 ;
    RECT 0 79.205 0.070 79.345 ;
    RECT 0 79.415 0.070 79.555 ;
    RECT 0 79.625 0.070 79.765 ;
    RECT 0 79.835 0.070 79.975 ;
    RECT 0 80.045 0.070 80.185 ;
    RECT 0 80.255 0.070 80.395 ;
    RECT 0 80.465 0.070 80.605 ;
    RECT 0 80.675 0.070 80.815 ;
    RECT 0 80.885 0.070 81.025 ;
    RECT 0 81.095 0.070 81.235 ;
    RECT 0 81.305 0.070 81.445 ;
    RECT 0 81.515 0.070 81.655 ;
    RECT 0 81.725 0.070 81.865 ;
    RECT 0 81.935 0.070 82.075 ;
    RECT 0 82.145 0.070 82.285 ;
    RECT 0 82.355 0.070 82.495 ;
    RECT 0 82.565 0.070 82.705 ;
    RECT 0 82.775 0.070 82.915 ;
    RECT 0 82.985 0.070 83.125 ;
    RECT 0 83.195 0.070 83.335 ;
    RECT 0 83.405 0.070 83.545 ;
    RECT 0 83.615 0.070 83.755 ;
    RECT 0 83.825 0.070 83.965 ;
    RECT 0 84.035 0.070 84.175 ;
    RECT 0 84.245 0.070 84.385 ;
    RECT 0 84.455 0.070 84.595 ;
    RECT 0 84.665 0.070 84.805 ;
    RECT 0 84.875 0.070 85.015 ;
    RECT 0 85.085 0.070 85.225 ;
    RECT 0 85.295 0.070 85.435 ;
    RECT 0 85.505 0.070 85.645 ;
    RECT 0 85.715 0.070 85.855 ;
    RECT 0 85.925 0.070 86.065 ;
    RECT 0 86.135 0.070 86.275 ;
    RECT 0 86.345 0.070 86.485 ;
    RECT 0 86.555 0.070 86.695 ;
    RECT 0 86.765 0.070 86.905 ;
    RECT 0 86.975 0.070 87.115 ;
    RECT 0 87.185 0.070 87.325 ;
    RECT 0 87.395 0.070 87.535 ;
    RECT 0 87.605 0.070 87.745 ;
    RECT 0 87.815 0.070 87.955 ;
    RECT 0 88.025 0.070 88.165 ;
    RECT 0 88.235 0.070 88.375 ;
    RECT 0 88.445 0.070 88.585 ;
    RECT 0 88.655 0.070 88.795 ;
    RECT 0 88.865 0.070 89.005 ;
    RECT 0 89.075 0.070 89.215 ;
    RECT 0 89.285 0.070 89.425 ;
    RECT 0 89.495 0.070 89.635 ;
    RECT 0 89.705 0.070 89.845 ;
    RECT 0 89.915 0.070 90.055 ;
    RECT 0 90.125 0.070 90.265 ;
    RECT 0 90.335 0.070 90.475 ;
    RECT 0 90.545 0.070 90.685 ;
    RECT 0 90.755 0.070 90.895 ;
    RECT 0 90.965 0.070 91.105 ;
    RECT 0 91.175 0.070 91.315 ;
    RECT 0 91.385 0.070 91.525 ;
    RECT 0 91.595 0.070 91.735 ;
    RECT 0 91.805 0.070 91.945 ;
    RECT 0 92.015 0.070 92.155 ;
    RECT 0 92.225 0.070 92.365 ;
    RECT 0 92.435 0.070 92.575 ;
    RECT 0 92.645 0.070 92.785 ;
    RECT 0 92.855 0.070 92.995 ;
    RECT 0 93.065 0.070 93.205 ;
    RECT 0 93.275 0.070 93.415 ;
    RECT 0 93.485 0.070 93.625 ;
    RECT 0 93.695 0.070 93.835 ;
    RECT 0 93.905 0.070 94.045 ;
    RECT 0 94.115 0.070 94.255 ;
    RECT 0 94.325 0.070 94.465 ;
    RECT 0 94.535 0.070 94.675 ;
    RECT 0 94.745 0.070 94.885 ;
    RECT 0 94.955 0.070 95.095 ;
    RECT 0 95.165 0.070 95.305 ;
    RECT 0 95.375 0.070 95.515 ;
    RECT 0 95.585 0.070 95.725 ;
    RECT 0 95.795 0.070 95.935 ;
    RECT 0 96.005 0.070 96.145 ;
    RECT 0 96.215 0.070 96.355 ;
    RECT 0 96.425 0.070 96.565 ;
    RECT 0 96.635 0.070 96.775 ;
    RECT 0 96.845 0.070 96.985 ;
    RECT 0 97.055 0.070 97.195 ;
    RECT 0 97.265 0.070 97.405 ;
    RECT 0 97.475 0.070 97.615 ;
    RECT 0 97.685 0.070 97.825 ;
    RECT 0 97.895 0.070 98.035 ;
    RECT 0 98.105 0.070 98.245 ;
    RECT 0 98.315 0.070 98.455 ;
    RECT 0 98.525 0.070 98.665 ;
    RECT 0 98.735 0.070 98.875 ;
    RECT 0 98.945 0.070 99.085 ;
    RECT 0 99.155 0.070 99.295 ;
    RECT 0 99.365 0.070 99.505 ;
    RECT 0 99.575 0.070 99.715 ;
    RECT 0 99.785 0.070 99.925 ;
    RECT 0 99.995 0.070 100.135 ;
    RECT 0 100.205 0.070 100.345 ;
    RECT 0 100.415 0.070 100.555 ;
    RECT 0 100.625 0.070 100.765 ;
    RECT 0 100.835 0.070 100.975 ;
    RECT 0 101.045 0.070 101.185 ;
    RECT 0 101.255 0.070 101.395 ;
    RECT 0 101.465 0.070 101.605 ;
    RECT 0 101.675 0.070 101.815 ;
    RECT 0 101.885 0.070 102.025 ;
    RECT 0 102.095 0.070 102.235 ;
    RECT 0 102.305 0.070 102.445 ;
    RECT 0 102.515 0.070 102.655 ;
    RECT 0 102.725 0.070 102.865 ;
    RECT 0 102.935 0.070 103.075 ;
    RECT 0 103.145 0.070 103.285 ;
    RECT 0 103.355 0.070 103.495 ;
    RECT 0 103.565 0.070 103.705 ;
    RECT 0 103.775 0.070 103.915 ;
    RECT 0 103.985 0.070 104.125 ;
    RECT 0 104.195 0.070 104.335 ;
    RECT 0 104.405 0.070 104.545 ;
    RECT 0 104.615 0.070 104.755 ;
    RECT 0 104.825 0.070 104.965 ;
    RECT 0 105.035 0.070 105.175 ;
    RECT 0 105.245 0.070 105.385 ;
    RECT 0 105.455 0.070 105.595 ;
    RECT 0 105.665 0.070 105.805 ;
    RECT 0 105.875 0.070 106.015 ;
    RECT 0 106.085 0.070 106.225 ;
    RECT 0 106.295 0.070 106.435 ;
    RECT 0 106.505 0.070 106.645 ;
    RECT 0 106.715 0.070 106.855 ;
    RECT 0 106.925 0.070 107.065 ;
    RECT 0 107.135 0.070 107.275 ;
    RECT 0 107.345 0.070 107.485 ;
    RECT 0 107.555 0.070 107.695 ;
    RECT 0 107.765 0.070 107.905 ;
    RECT 0 107.975 0.070 108.115 ;
    RECT 0 108.185 0.070 108.325 ;
    RECT 0 108.395 0.070 108.535 ;
    RECT 0 108.605 0.070 108.745 ;
    RECT 0 108.815 0.070 108.955 ;
    RECT 0 109.025 0.070 109.165 ;
    RECT 0 109.235 0.070 109.375 ;
    RECT 0 109.445 0.070 109.585 ;
    RECT 0 109.655 0.070 109.795 ;
    RECT 0 109.865 0.070 110.005 ;
    RECT 0 110.075 0.070 110.215 ;
    RECT 0 110.285 0.070 110.425 ;
    RECT 0 110.495 0.070 110.635 ;
    RECT 0 110.705 0.070 110.845 ;
    RECT 0 110.915 0.070 111.055 ;
    RECT 0 111.125 0.070 111.265 ;
    RECT 0 111.335 0.070 111.475 ;
    RECT 0 111.545 0.070 111.685 ;
    RECT 0 111.755 0.070 111.895 ;
    RECT 0 111.965 0.070 112.105 ;
    RECT 0 112.175 0.070 112.315 ;
    RECT 0 112.385 0.070 112.525 ;
    RECT 0 112.595 0.070 112.735 ;
    RECT 0 112.805 0.070 112.945 ;
    RECT 0 113.015 0.070 113.155 ;
    RECT 0 113.225 0.070 113.365 ;
    RECT 0 113.435 0.070 113.575 ;
    RECT 0 113.645 0.070 113.785 ;
    RECT 0 113.855 0.070 113.995 ;
    RECT 0 114.065 0.070 114.205 ;
    RECT 0 114.275 0.070 114.415 ;
    RECT 0 114.485 0.070 114.625 ;
    RECT 0 114.695 0.070 114.835 ;
    RECT 0 114.905 0.070 115.045 ;
    RECT 0 115.115 0.070 115.255 ;
    RECT 0 115.325 0.070 115.465 ;
    RECT 0 115.535 0.070 115.675 ;
    RECT 0 115.745 0.070 115.885 ;
    RECT 0 115.955 0.070 116.095 ;
    RECT 0 116.165 0.070 116.305 ;
    RECT 0 116.375 0.070 116.515 ;
    RECT 0 116.585 0.070 116.725 ;
    RECT 0 116.795 0.070 116.935 ;
    RECT 0 117.005 0.070 117.145 ;
    RECT 0 117.215 0.070 117.355 ;
    RECT 0 117.425 0.070 117.565 ;
    RECT 0 117.635 0.070 117.775 ;
    RECT 0 117.845 0.070 117.985 ;
    RECT 0 118.055 0.070 118.195 ;
    RECT 0 118.265 0.070 118.405 ;
    RECT 0 118.475 0.070 118.615 ;
    RECT 0 118.685 0.070 118.825 ;
    RECT 0 118.895 0.070 119.035 ;
    RECT 0 119.105 0.070 119.245 ;
    RECT 0 119.315 0.070 119.455 ;
    RECT 0 119.525 0.070 119.665 ;
    RECT 0 119.735 0.070 119.875 ;
    RECT 0 119.945 0.070 120.085 ;
    RECT 0 120.155 0.070 120.295 ;
    RECT 0 120.365 0.070 120.505 ;
    RECT 0 120.575 0.070 120.715 ;
    RECT 0 120.785 0.070 120.925 ;
    RECT 0 120.995 0.070 121.135 ;
    RECT 0 121.205 0.070 121.345 ;
    RECT 0 121.415 0.070 121.555 ;
    RECT 0 121.625 0.070 121.765 ;
    RECT 0 121.835 0.070 121.975 ;
    RECT 0 122.045 0.070 122.185 ;
    RECT 0 122.255 0.070 122.395 ;
    RECT 0 122.465 0.070 122.605 ;
    RECT 0 122.675 0.070 122.815 ;
    RECT 0 122.885 0.070 123.025 ;
    RECT 0 123.095 0.070 123.235 ;
    RECT 0 123.305 0.070 123.445 ;
    RECT 0 123.515 0.070 123.655 ;
    RECT 0 123.725 0.070 123.865 ;
    RECT 0 123.935 0.070 124.075 ;
    RECT 0 124.145 0.070 124.285 ;
    RECT 0 124.355 0.070 124.495 ;
    RECT 0 124.565 0.070 124.705 ;
    RECT 0 124.775 0.070 124.915 ;
    RECT 0 124.985 0.070 125.125 ;
    RECT 0 125.195 0.070 125.335 ;
    RECT 0 125.405 0.070 125.545 ;
    RECT 0 125.615 0.070 125.755 ;
    RECT 0 125.825 0.070 125.965 ;
    RECT 0 126.035 0.070 126.175 ;
    RECT 0 126.245 0.070 126.385 ;
    RECT 0 126.455 0.070 126.595 ;
    RECT 0 126.665 0.070 144.025 ;
    RECT 0 144.095 0.070 144.235 ;
    RECT 0 144.305 0.070 144.445 ;
    RECT 0 144.515 0.070 144.655 ;
    RECT 0 144.725 0.070 144.865 ;
    RECT 0 144.935 0.070 145.075 ;
    RECT 0 145.145 0.070 145.285 ;
    RECT 0 145.355 0.070 145.495 ;
    RECT 0 145.565 0.070 145.705 ;
    RECT 0 145.775 0.070 145.915 ;
    RECT 0 145.985 0.070 146.125 ;
    RECT 0 146.195 0.070 146.335 ;
    RECT 0 146.405 0.070 146.545 ;
    RECT 0 146.615 0.070 146.755 ;
    RECT 0 146.825 0.070 146.965 ;
    RECT 0 147.035 0.070 147.175 ;
    RECT 0 147.245 0.070 147.385 ;
    RECT 0 147.455 0.070 147.595 ;
    RECT 0 147.665 0.070 147.805 ;
    RECT 0 147.875 0.070 148.015 ;
    RECT 0 148.085 0.070 148.225 ;
    RECT 0 148.295 0.070 148.435 ;
    RECT 0 148.505 0.070 148.645 ;
    RECT 0 148.715 0.070 148.855 ;
    RECT 0 148.925 0.070 149.065 ;
    RECT 0 149.135 0.070 149.275 ;
    RECT 0 149.345 0.070 149.485 ;
    RECT 0 149.555 0.070 149.695 ;
    RECT 0 149.765 0.070 149.905 ;
    RECT 0 149.975 0.070 150.115 ;
    RECT 0 150.185 0.070 150.325 ;
    RECT 0 150.395 0.070 150.535 ;
    RECT 0 150.605 0.070 150.745 ;
    RECT 0 150.815 0.070 150.955 ;
    RECT 0 151.025 0.070 151.165 ;
    RECT 0 151.235 0.070 151.375 ;
    RECT 0 151.445 0.070 151.585 ;
    RECT 0 151.655 0.070 151.795 ;
    RECT 0 151.865 0.070 152.005 ;
    RECT 0 152.075 0.070 152.215 ;
    RECT 0 152.285 0.070 152.425 ;
    RECT 0 152.495 0.070 152.635 ;
    RECT 0 152.705 0.070 152.845 ;
    RECT 0 152.915 0.070 153.055 ;
    RECT 0 153.125 0.070 153.265 ;
    RECT 0 153.335 0.070 153.475 ;
    RECT 0 153.545 0.070 153.685 ;
    RECT 0 153.755 0.070 153.895 ;
    RECT 0 153.965 0.070 154.105 ;
    RECT 0 154.175 0.070 154.315 ;
    RECT 0 154.385 0.070 154.525 ;
    RECT 0 154.595 0.070 154.735 ;
    RECT 0 154.805 0.070 154.945 ;
    RECT 0 155.015 0.070 155.155 ;
    RECT 0 155.225 0.070 155.365 ;
    RECT 0 155.435 0.070 155.575 ;
    RECT 0 155.645 0.070 155.785 ;
    RECT 0 155.855 0.070 155.995 ;
    RECT 0 156.065 0.070 156.205 ;
    RECT 0 156.275 0.070 156.415 ;
    RECT 0 156.485 0.070 156.625 ;
    RECT 0 156.695 0.070 156.835 ;
    RECT 0 156.905 0.070 157.045 ;
    RECT 0 157.115 0.070 157.255 ;
    RECT 0 157.325 0.070 157.465 ;
    RECT 0 157.535 0.070 157.675 ;
    RECT 0 157.745 0.070 157.885 ;
    RECT 0 157.955 0.070 158.095 ;
    RECT 0 158.165 0.070 158.305 ;
    RECT 0 158.375 0.070 158.515 ;
    RECT 0 158.585 0.070 158.725 ;
    RECT 0 158.795 0.070 158.935 ;
    RECT 0 159.005 0.070 159.145 ;
    RECT 0 159.215 0.070 159.355 ;
    RECT 0 159.425 0.070 159.565 ;
    RECT 0 159.635 0.070 159.775 ;
    RECT 0 159.845 0.070 159.985 ;
    RECT 0 160.055 0.070 160.195 ;
    RECT 0 160.265 0.070 160.405 ;
    RECT 0 160.475 0.070 160.615 ;
    RECT 0 160.685 0.070 160.825 ;
    RECT 0 160.895 0.070 161.035 ;
    RECT 0 161.105 0.070 161.245 ;
    RECT 0 161.315 0.070 161.455 ;
    RECT 0 161.525 0.070 161.665 ;
    RECT 0 161.735 0.070 161.875 ;
    RECT 0 161.945 0.070 162.085 ;
    RECT 0 162.155 0.070 162.295 ;
    RECT 0 162.365 0.070 162.505 ;
    RECT 0 162.575 0.070 162.715 ;
    RECT 0 162.785 0.070 162.925 ;
    RECT 0 162.995 0.070 163.135 ;
    RECT 0 163.205 0.070 163.345 ;
    RECT 0 163.415 0.070 163.555 ;
    RECT 0 163.625 0.070 163.765 ;
    RECT 0 163.835 0.070 163.975 ;
    RECT 0 164.045 0.070 164.185 ;
    RECT 0 164.255 0.070 164.395 ;
    RECT 0 164.465 0.070 164.605 ;
    RECT 0 164.675 0.070 164.815 ;
    RECT 0 164.885 0.070 165.025 ;
    RECT 0 165.095 0.070 165.235 ;
    RECT 0 165.305 0.070 165.445 ;
    RECT 0 165.515 0.070 165.655 ;
    RECT 0 165.725 0.070 165.865 ;
    RECT 0 165.935 0.070 166.075 ;
    RECT 0 166.145 0.070 166.285 ;
    RECT 0 166.355 0.070 166.495 ;
    RECT 0 166.565 0.070 166.705 ;
    RECT 0 166.775 0.070 166.915 ;
    RECT 0 166.985 0.070 167.125 ;
    RECT 0 167.195 0.070 167.335 ;
    RECT 0 167.405 0.070 167.545 ;
    RECT 0 167.615 0.070 167.755 ;
    RECT 0 167.825 0.070 167.965 ;
    RECT 0 168.035 0.070 168.175 ;
    RECT 0 168.245 0.070 168.385 ;
    RECT 0 168.455 0.070 168.595 ;
    RECT 0 168.665 0.070 168.805 ;
    RECT 0 168.875 0.070 169.015 ;
    RECT 0 169.085 0.070 169.225 ;
    RECT 0 169.295 0.070 169.435 ;
    RECT 0 169.505 0.070 169.645 ;
    RECT 0 169.715 0.070 169.855 ;
    RECT 0 169.925 0.070 170.065 ;
    RECT 0 170.135 0.070 170.275 ;
    RECT 0 170.345 0.070 170.485 ;
    RECT 0 170.555 0.070 170.695 ;
    RECT 0 170.765 0.070 170.905 ;
    RECT 0 170.975 0.070 171.115 ;
    RECT 0 171.185 0.070 171.325 ;
    RECT 0 171.395 0.070 171.535 ;
    RECT 0 171.605 0.070 171.745 ;
    RECT 0 171.815 0.070 171.955 ;
    RECT 0 172.025 0.070 172.165 ;
    RECT 0 172.235 0.070 172.375 ;
    RECT 0 172.445 0.070 172.585 ;
    RECT 0 172.655 0.070 172.795 ;
    RECT 0 172.865 0.070 173.005 ;
    RECT 0 173.075 0.070 173.215 ;
    RECT 0 173.285 0.070 173.425 ;
    RECT 0 173.495 0.070 173.635 ;
    RECT 0 173.705 0.070 173.845 ;
    RECT 0 173.915 0.070 174.055 ;
    RECT 0 174.125 0.070 174.265 ;
    RECT 0 174.335 0.070 174.475 ;
    RECT 0 174.545 0.070 174.685 ;
    RECT 0 174.755 0.070 174.895 ;
    RECT 0 174.965 0.070 175.105 ;
    RECT 0 175.175 0.070 175.315 ;
    RECT 0 175.385 0.070 175.525 ;
    RECT 0 175.595 0.070 175.735 ;
    RECT 0 175.805 0.070 175.945 ;
    RECT 0 176.015 0.070 176.155 ;
    RECT 0 176.225 0.070 176.365 ;
    RECT 0 176.435 0.070 176.575 ;
    RECT 0 176.645 0.070 176.785 ;
    RECT 0 176.855 0.070 176.995 ;
    RECT 0 177.065 0.070 177.205 ;
    RECT 0 177.275 0.070 177.415 ;
    RECT 0 177.485 0.070 177.625 ;
    RECT 0 177.695 0.070 177.835 ;
    RECT 0 177.905 0.070 178.045 ;
    RECT 0 178.115 0.070 178.255 ;
    RECT 0 178.325 0.070 178.465 ;
    RECT 0 178.535 0.070 178.675 ;
    RECT 0 178.745 0.070 178.885 ;
    RECT 0 178.955 0.070 179.095 ;
    RECT 0 179.165 0.070 179.305 ;
    RECT 0 179.375 0.070 179.515 ;
    RECT 0 179.585 0.070 179.725 ;
    RECT 0 179.795 0.070 179.935 ;
    RECT 0 180.005 0.070 180.145 ;
    RECT 0 180.215 0.070 180.355 ;
    RECT 0 180.425 0.070 180.565 ;
    RECT 0 180.635 0.070 180.775 ;
    RECT 0 180.845 0.070 180.985 ;
    RECT 0 181.055 0.070 181.195 ;
    RECT 0 181.265 0.070 181.405 ;
    RECT 0 181.475 0.070 181.615 ;
    RECT 0 181.685 0.070 181.825 ;
    RECT 0 181.895 0.070 182.035 ;
    RECT 0 182.105 0.070 182.245 ;
    RECT 0 182.315 0.070 182.455 ;
    RECT 0 182.525 0.070 182.665 ;
    RECT 0 182.735 0.070 182.875 ;
    RECT 0 182.945 0.070 183.085 ;
    RECT 0 183.155 0.070 183.295 ;
    RECT 0 183.365 0.070 183.505 ;
    RECT 0 183.575 0.070 183.715 ;
    RECT 0 183.785 0.070 183.925 ;
    RECT 0 183.995 0.070 184.135 ;
    RECT 0 184.205 0.070 184.345 ;
    RECT 0 184.415 0.070 184.555 ;
    RECT 0 184.625 0.070 184.765 ;
    RECT 0 184.835 0.070 184.975 ;
    RECT 0 185.045 0.070 185.185 ;
    RECT 0 185.255 0.070 185.395 ;
    RECT 0 185.465 0.070 185.605 ;
    RECT 0 185.675 0.070 185.815 ;
    RECT 0 185.885 0.070 186.025 ;
    RECT 0 186.095 0.070 186.235 ;
    RECT 0 186.305 0.070 186.445 ;
    RECT 0 186.515 0.070 186.655 ;
    RECT 0 186.725 0.070 186.865 ;
    RECT 0 186.935 0.070 187.075 ;
    RECT 0 187.145 0.070 187.285 ;
    RECT 0 187.355 0.070 187.495 ;
    RECT 0 187.565 0.070 187.705 ;
    RECT 0 187.775 0.070 187.915 ;
    RECT 0 187.985 0.070 188.125 ;
    RECT 0 188.195 0.070 188.335 ;
    RECT 0 188.405 0.070 188.545 ;
    RECT 0 188.615 0.070 188.755 ;
    RECT 0 188.825 0.070 188.965 ;
    RECT 0 189.035 0.070 189.175 ;
    RECT 0 189.245 0.070 189.385 ;
    RECT 0 189.455 0.070 189.595 ;
    RECT 0 189.665 0.070 189.805 ;
    RECT 0 189.875 0.070 190.015 ;
    RECT 0 190.085 0.070 190.225 ;
    RECT 0 190.295 0.070 190.435 ;
    RECT 0 190.505 0.070 190.645 ;
    RECT 0 190.715 0.070 190.855 ;
    RECT 0 190.925 0.070 191.065 ;
    RECT 0 191.135 0.070 191.275 ;
    RECT 0 191.345 0.070 191.485 ;
    RECT 0 191.555 0.070 191.695 ;
    RECT 0 191.765 0.070 191.905 ;
    RECT 0 191.975 0.070 192.115 ;
    RECT 0 192.185 0.070 192.325 ;
    RECT 0 192.395 0.070 192.535 ;
    RECT 0 192.605 0.070 192.745 ;
    RECT 0 192.815 0.070 192.955 ;
    RECT 0 193.025 0.070 193.165 ;
    RECT 0 193.235 0.070 193.375 ;
    RECT 0 193.445 0.070 193.585 ;
    RECT 0 193.655 0.070 193.795 ;
    RECT 0 193.865 0.070 194.005 ;
    RECT 0 194.075 0.070 194.215 ;
    RECT 0 194.285 0.070 194.425 ;
    RECT 0 194.495 0.070 194.635 ;
    RECT 0 194.705 0.070 194.845 ;
    RECT 0 194.915 0.070 195.055 ;
    RECT 0 195.125 0.070 195.265 ;
    RECT 0 195.335 0.070 195.475 ;
    RECT 0 195.545 0.070 195.685 ;
    RECT 0 195.755 0.070 195.895 ;
    RECT 0 195.965 0.070 196.105 ;
    RECT 0 196.175 0.070 196.315 ;
    RECT 0 196.385 0.070 196.525 ;
    RECT 0 196.595 0.070 196.735 ;
    RECT 0 196.805 0.070 196.945 ;
    RECT 0 197.015 0.070 197.155 ;
    RECT 0 197.225 0.070 197.365 ;
    RECT 0 197.435 0.070 197.575 ;
    RECT 0 197.645 0.070 215.005 ;
    RECT 0 215.075 0.070 215.215 ;
    RECT 0 215.285 0.070 215.425 ;
    RECT 0 215.495 0.070 215.635 ;
    RECT 0 215.705 0.070 215.845 ;
    RECT 0 215.915 0.070 216.055 ;
    RECT 0 216.125 0.070 216.265 ;
    RECT 0 216.335 0.070 233.695 ;
    RECT 0 233.765 0.070 233.905 ;
    RECT 0 233.975 0.070 234.115 ;
    RECT 0 234.185 0.070 238.000 ;
    LAYER metal4 ;
    RECT 0 0 153.710 2.100 ;
    RECT 0 235.900 153.710 238.000 ;
    RECT 0.000 2.100 1.960 235.900 ;
    RECT 2.240 2.100 3.640 235.900 ;
    RECT 3.920 2.100 5.320 235.900 ;
    RECT 5.600 2.100 7.000 235.900 ;
    RECT 7.280 2.100 8.680 235.900 ;
    RECT 8.960 2.100 10.360 235.900 ;
    RECT 10.640 2.100 12.040 235.900 ;
    RECT 12.320 2.100 13.720 235.900 ;
    RECT 14.000 2.100 15.400 235.900 ;
    RECT 15.680 2.100 17.080 235.900 ;
    RECT 17.360 2.100 18.760 235.900 ;
    RECT 19.040 2.100 20.440 235.900 ;
    RECT 20.720 2.100 22.120 235.900 ;
    RECT 22.400 2.100 23.800 235.900 ;
    RECT 24.080 2.100 25.480 235.900 ;
    RECT 25.760 2.100 27.160 235.900 ;
    RECT 27.440 2.100 28.840 235.900 ;
    RECT 29.120 2.100 30.520 235.900 ;
    RECT 30.800 2.100 32.200 235.900 ;
    RECT 32.480 2.100 33.880 235.900 ;
    RECT 34.160 2.100 35.560 235.900 ;
    RECT 35.840 2.100 37.240 235.900 ;
    RECT 37.520 2.100 38.920 235.900 ;
    RECT 39.200 2.100 40.600 235.900 ;
    RECT 40.880 2.100 42.280 235.900 ;
    RECT 42.560 2.100 43.960 235.900 ;
    RECT 44.240 2.100 45.640 235.900 ;
    RECT 45.920 2.100 47.320 235.900 ;
    RECT 47.600 2.100 49.000 235.900 ;
    RECT 49.280 2.100 50.680 235.900 ;
    RECT 50.960 2.100 52.360 235.900 ;
    RECT 52.640 2.100 54.040 235.900 ;
    RECT 54.320 2.100 55.720 235.900 ;
    RECT 56.000 2.100 57.400 235.900 ;
    RECT 57.680 2.100 59.080 235.900 ;
    RECT 59.360 2.100 60.760 235.900 ;
    RECT 61.040 2.100 62.440 235.900 ;
    RECT 62.720 2.100 64.120 235.900 ;
    RECT 64.400 2.100 65.800 235.900 ;
    RECT 66.080 2.100 67.480 235.900 ;
    RECT 67.760 2.100 69.160 235.900 ;
    RECT 69.440 2.100 70.840 235.900 ;
    RECT 71.120 2.100 72.520 235.900 ;
    RECT 72.800 2.100 74.200 235.900 ;
    RECT 74.480 2.100 75.880 235.900 ;
    RECT 76.160 2.100 77.560 235.900 ;
    RECT 77.840 2.100 79.240 235.900 ;
    RECT 79.520 2.100 80.920 235.900 ;
    RECT 81.200 2.100 82.600 235.900 ;
    RECT 82.880 2.100 84.280 235.900 ;
    RECT 84.560 2.100 85.960 235.900 ;
    RECT 86.240 2.100 87.640 235.900 ;
    RECT 87.920 2.100 89.320 235.900 ;
    RECT 89.600 2.100 91.000 235.900 ;
    RECT 91.280 2.100 92.680 235.900 ;
    RECT 92.960 2.100 94.360 235.900 ;
    RECT 94.640 2.100 96.040 235.900 ;
    RECT 96.320 2.100 97.720 235.900 ;
    RECT 98.000 2.100 99.400 235.900 ;
    RECT 99.680 2.100 101.080 235.900 ;
    RECT 101.360 2.100 102.760 235.900 ;
    RECT 103.040 2.100 104.440 235.900 ;
    RECT 104.720 2.100 106.120 235.900 ;
    RECT 106.400 2.100 107.800 235.900 ;
    RECT 108.080 2.100 109.480 235.900 ;
    RECT 109.760 2.100 111.160 235.900 ;
    RECT 111.440 2.100 112.840 235.900 ;
    RECT 113.120 2.100 114.520 235.900 ;
    RECT 114.800 2.100 116.200 235.900 ;
    RECT 116.480 2.100 117.880 235.900 ;
    RECT 118.160 2.100 119.560 235.900 ;
    RECT 119.840 2.100 121.240 235.900 ;
    RECT 121.520 2.100 122.920 235.900 ;
    RECT 123.200 2.100 124.600 235.900 ;
    RECT 124.880 2.100 126.280 235.900 ;
    RECT 126.560 2.100 127.960 235.900 ;
    RECT 128.240 2.100 129.640 235.900 ;
    RECT 129.920 2.100 131.320 235.900 ;
    RECT 131.600 2.100 133.000 235.900 ;
    RECT 133.280 2.100 134.680 235.900 ;
    RECT 134.960 2.100 136.360 235.900 ;
    RECT 136.640 2.100 138.040 235.900 ;
    RECT 138.320 2.100 139.720 235.900 ;
    RECT 140.000 2.100 141.400 235.900 ;
    RECT 141.680 2.100 143.080 235.900 ;
    RECT 143.360 2.100 144.760 235.900 ;
    RECT 145.040 2.100 146.440 235.900 ;
    RECT 146.720 2.100 148.120 235.900 ;
    RECT 148.400 2.100 149.800 235.900 ;
    RECT 150.080 2.100 153.710 235.900 ;
    LAYER OVERLAP ;
    RECT 0 0 153.710 238.000 ;
  END
END fakeram45_128x256

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_128x116
  FOREIGN fakeram45_128x116 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 121.030 BY 117.600 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.275 0.070 2.345 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.695 0.070 2.765 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.115 0.070 3.185 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.535 0.070 3.605 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.955 0.070 4.025 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.375 0.070 4.445 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.795 0.070 4.865 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.215 0.070 5.285 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.635 0.070 5.705 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.055 0.070 6.125 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.475 0.070 6.545 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.895 0.070 6.965 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.315 0.070 7.385 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.735 0.070 7.805 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.155 0.070 8.225 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.575 0.070 8.645 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.785 0.070 8.855 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.995 0.070 9.065 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.415 0.070 9.485 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.835 0.070 9.905 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.255 0.070 10.325 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.675 0.070 10.745 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.095 0.070 11.165 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.515 0.070 11.585 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.935 0.070 12.005 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.355 0.070 12.425 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.775 0.070 12.845 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.985 0.070 13.055 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.195 0.070 13.265 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.615 0.070 13.685 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.035 0.070 14.105 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.455 0.070 14.525 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.875 0.070 14.945 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.295 0.070 15.365 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.505 0.070 15.575 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.715 0.070 15.785 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.135 0.070 16.205 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.345 0.070 16.415 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.555 0.070 16.625 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.975 0.070 17.045 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.185 0.070 17.255 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.395 0.070 17.465 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.605 0.070 17.675 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.815 0.070 17.885 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.025 0.070 18.095 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.235 0.070 18.305 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.655 0.070 18.725 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.075 0.070 19.145 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.495 0.070 19.565 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.915 0.070 19.985 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.335 0.070 20.405 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.545 0.070 20.615 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.755 0.070 20.825 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.175 0.070 21.245 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.595 0.070 21.665 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.015 0.070 22.085 ;
    END
  END w_mask_in[95]
  PIN w_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.225 0.070 22.295 ;
    END
  END w_mask_in[96]
  PIN w_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.435 0.070 22.505 ;
    END
  END w_mask_in[97]
  PIN w_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END w_mask_in[98]
  PIN w_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.855 0.070 22.925 ;
    END
  END w_mask_in[99]
  PIN w_mask_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END w_mask_in[100]
  PIN w_mask_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.275 0.070 23.345 ;
    END
  END w_mask_in[101]
  PIN w_mask_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END w_mask_in[102]
  PIN w_mask_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.695 0.070 23.765 ;
    END
  END w_mask_in[103]
  PIN w_mask_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.905 0.070 23.975 ;
    END
  END w_mask_in[104]
  PIN w_mask_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.115 0.070 24.185 ;
    END
  END w_mask_in[105]
  PIN w_mask_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END w_mask_in[106]
  PIN w_mask_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.535 0.070 24.605 ;
    END
  END w_mask_in[107]
  PIN w_mask_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END w_mask_in[108]
  PIN w_mask_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.955 0.070 25.025 ;
    END
  END w_mask_in[109]
  PIN w_mask_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END w_mask_in[110]
  PIN w_mask_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.375 0.070 25.445 ;
    END
  END w_mask_in[111]
  PIN w_mask_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END w_mask_in[112]
  PIN w_mask_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.795 0.070 25.865 ;
    END
  END w_mask_in[113]
  PIN w_mask_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END w_mask_in[114]
  PIN w_mask_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.215 0.070 26.285 ;
    END
  END w_mask_in[115]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.875 0.070 35.945 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.295 0.070 36.365 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.505 0.070 36.575 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.715 0.070 36.785 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.135 0.070 37.205 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.555 0.070 37.625 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.975 0.070 38.045 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.185 0.070 38.255 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.395 0.070 38.465 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.815 0.070 38.885 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.235 0.070 39.305 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.655 0.070 39.725 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.075 0.070 40.145 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.495 0.070 40.565 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.915 0.070 40.985 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.335 0.070 41.405 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.755 0.070 41.825 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.175 0.070 42.245 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.595 0.070 42.665 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.015 0.070 43.085 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.435 0.070 43.505 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.855 0.070 43.925 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.275 0.070 44.345 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.695 0.070 44.765 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.115 0.070 45.185 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.325 0.070 45.395 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.535 0.070 45.605 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.745 0.070 45.815 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.955 0.070 46.025 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.375 0.070 46.445 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.585 0.070 46.655 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.795 0.070 46.865 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.215 0.070 47.285 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.635 0.070 47.705 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.055 0.070 48.125 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.265 0.070 48.335 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.475 0.070 48.545 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.895 0.070 48.965 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.315 0.070 49.385 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.735 0.070 49.805 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.945 0.070 50.015 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.155 0.070 50.225 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.575 0.070 50.645 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.785 0.070 50.855 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.995 0.070 51.065 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.205 0.070 51.275 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.415 0.070 51.485 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.625 0.070 51.695 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.835 0.070 51.905 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.045 0.070 52.115 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.255 0.070 52.325 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.675 0.070 52.745 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.095 0.070 53.165 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.305 0.070 53.375 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.515 0.070 53.585 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.935 0.070 54.005 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.145 0.070 54.215 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.355 0.070 54.425 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.775 0.070 54.845 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.985 0.070 55.055 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.195 0.070 55.265 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.615 0.070 55.685 ;
    END
  END rd_out[95]
  PIN rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.825 0.070 55.895 ;
    END
  END rd_out[96]
  PIN rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.035 0.070 56.105 ;
    END
  END rd_out[97]
  PIN rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END rd_out[98]
  PIN rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.455 0.070 56.525 ;
    END
  END rd_out[99]
  PIN rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.665 0.070 56.735 ;
    END
  END rd_out[100]
  PIN rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.875 0.070 56.945 ;
    END
  END rd_out[101]
  PIN rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.085 0.070 57.155 ;
    END
  END rd_out[102]
  PIN rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.295 0.070 57.365 ;
    END
  END rd_out[103]
  PIN rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.505 0.070 57.575 ;
    END
  END rd_out[104]
  PIN rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.715 0.070 57.785 ;
    END
  END rd_out[105]
  PIN rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END rd_out[106]
  PIN rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.135 0.070 58.205 ;
    END
  END rd_out[107]
  PIN rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.345 0.070 58.415 ;
    END
  END rd_out[108]
  PIN rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.555 0.070 58.625 ;
    END
  END rd_out[109]
  PIN rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.765 0.070 58.835 ;
    END
  END rd_out[110]
  PIN rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.975 0.070 59.045 ;
    END
  END rd_out[111]
  PIN rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.185 0.070 59.255 ;
    END
  END rd_out[112]
  PIN rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.395 0.070 59.465 ;
    END
  END rd_out[113]
  PIN rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.605 0.070 59.675 ;
    END
  END rd_out[114]
  PIN rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.815 0.070 59.885 ;
    END
  END rd_out[115]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.265 0.070 69.335 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.475 0.070 69.545 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.685 0.070 69.755 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.895 0.070 69.965 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.105 0.070 70.175 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.315 0.070 70.385 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.735 0.070 70.805 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.945 0.070 71.015 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.155 0.070 71.225 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.575 0.070 71.645 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.785 0.070 71.855 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.995 0.070 72.065 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.205 0.070 72.275 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.415 0.070 72.485 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.625 0.070 72.695 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.835 0.070 72.905 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.255 0.070 73.325 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.465 0.070 73.535 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.675 0.070 73.745 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.095 0.070 74.165 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.305 0.070 74.375 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.515 0.070 74.585 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.725 0.070 74.795 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.935 0.070 75.005 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.145 0.070 75.215 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.355 0.070 75.425 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.775 0.070 75.845 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.195 0.070 76.265 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.405 0.070 76.475 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.615 0.070 76.685 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.825 0.070 76.895 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.035 0.070 77.105 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.245 0.070 77.315 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.455 0.070 77.525 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.665 0.070 77.735 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.875 0.070 77.945 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.085 0.070 78.155 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.295 0.070 78.365 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.505 0.070 78.575 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.715 0.070 78.785 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.925 0.070 78.995 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.135 0.070 79.205 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.345 0.070 79.415 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.555 0.070 79.625 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.975 0.070 80.045 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.185 0.070 80.255 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.395 0.070 80.465 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.605 0.070 80.675 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.815 0.070 80.885 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.025 0.070 81.095 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.235 0.070 81.305 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.445 0.070 81.515 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.655 0.070 81.725 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.075 0.070 82.145 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.285 0.070 82.355 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.495 0.070 82.565 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.705 0.070 82.775 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.915 0.070 82.985 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.125 0.070 83.195 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.335 0.070 83.405 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.545 0.070 83.615 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.755 0.070 83.825 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.965 0.070 84.035 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.175 0.070 84.245 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.385 0.070 84.455 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.595 0.070 84.665 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.015 0.070 85.085 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.225 0.070 85.295 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.435 0.070 85.505 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.855 0.070 85.925 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.065 0.070 86.135 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.275 0.070 86.345 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.485 0.070 86.555 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.695 0.070 86.765 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.905 0.070 86.975 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.115 0.070 87.185 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.325 0.070 87.395 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.535 0.070 87.605 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.745 0.070 87.815 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.955 0.070 88.025 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.165 0.070 88.235 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.375 0.070 88.445 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.585 0.070 88.655 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.795 0.070 88.865 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.005 0.070 89.075 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.215 0.070 89.285 ;
    END
  END wd_in[95]
  PIN wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.425 0.070 89.495 ;
    END
  END wd_in[96]
  PIN wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.635 0.070 89.705 ;
    END
  END wd_in[97]
  PIN wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.845 0.070 89.915 ;
    END
  END wd_in[98]
  PIN wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.055 0.070 90.125 ;
    END
  END wd_in[99]
  PIN wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.265 0.070 90.335 ;
    END
  END wd_in[100]
  PIN wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.475 0.070 90.545 ;
    END
  END wd_in[101]
  PIN wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.685 0.070 90.755 ;
    END
  END wd_in[102]
  PIN wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.895 0.070 90.965 ;
    END
  END wd_in[103]
  PIN wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.105 0.070 91.175 ;
    END
  END wd_in[104]
  PIN wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.315 0.070 91.385 ;
    END
  END wd_in[105]
  PIN wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.525 0.070 91.595 ;
    END
  END wd_in[106]
  PIN wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.735 0.070 91.805 ;
    END
  END wd_in[107]
  PIN wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.945 0.070 92.015 ;
    END
  END wd_in[108]
  PIN wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.155 0.070 92.225 ;
    END
  END wd_in[109]
  PIN wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.365 0.070 92.435 ;
    END
  END wd_in[110]
  PIN wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.575 0.070 92.645 ;
    END
  END wd_in[111]
  PIN wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.785 0.070 92.855 ;
    END
  END wd_in[112]
  PIN wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.995 0.070 93.065 ;
    END
  END wd_in[113]
  PIN wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.205 0.070 93.275 ;
    END
  END wd_in[114]
  PIN wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.415 0.070 93.485 ;
    END
  END wd_in[115]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.865 0.070 102.935 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.075 0.070 103.145 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.285 0.070 103.355 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.495 0.070 103.565 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.705 0.070 103.775 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 103.915 0.070 103.985 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.125 0.070 104.195 ;
    END
  END addr_in[6]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.575 0.070 113.645 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.785 0.070 113.855 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.995 0.070 114.065 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 115.500 ;
      RECT 5.320 2.100 5.600 115.500 ;
      RECT 8.680 2.100 8.960 115.500 ;
      RECT 12.040 2.100 12.320 115.500 ;
      RECT 15.400 2.100 15.680 115.500 ;
      RECT 18.760 2.100 19.040 115.500 ;
      RECT 22.120 2.100 22.400 115.500 ;
      RECT 25.480 2.100 25.760 115.500 ;
      RECT 28.840 2.100 29.120 115.500 ;
      RECT 32.200 2.100 32.480 115.500 ;
      RECT 35.560 2.100 35.840 115.500 ;
      RECT 38.920 2.100 39.200 115.500 ;
      RECT 42.280 2.100 42.560 115.500 ;
      RECT 45.640 2.100 45.920 115.500 ;
      RECT 49.000 2.100 49.280 115.500 ;
      RECT 52.360 2.100 52.640 115.500 ;
      RECT 55.720 2.100 56.000 115.500 ;
      RECT 59.080 2.100 59.360 115.500 ;
      RECT 62.440 2.100 62.720 115.500 ;
      RECT 65.800 2.100 66.080 115.500 ;
      RECT 69.160 2.100 69.440 115.500 ;
      RECT 72.520 2.100 72.800 115.500 ;
      RECT 75.880 2.100 76.160 115.500 ;
      RECT 79.240 2.100 79.520 115.500 ;
      RECT 82.600 2.100 82.880 115.500 ;
      RECT 85.960 2.100 86.240 115.500 ;
      RECT 89.320 2.100 89.600 115.500 ;
      RECT 92.680 2.100 92.960 115.500 ;
      RECT 96.040 2.100 96.320 115.500 ;
      RECT 99.400 2.100 99.680 115.500 ;
      RECT 102.760 2.100 103.040 115.500 ;
      RECT 106.120 2.100 106.400 115.500 ;
      RECT 109.480 2.100 109.760 115.500 ;
      RECT 112.840 2.100 113.120 115.500 ;
      RECT 116.200 2.100 116.480 115.500 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 115.500 ;
      RECT 7.000 2.100 7.280 115.500 ;
      RECT 10.360 2.100 10.640 115.500 ;
      RECT 13.720 2.100 14.000 115.500 ;
      RECT 17.080 2.100 17.360 115.500 ;
      RECT 20.440 2.100 20.720 115.500 ;
      RECT 23.800 2.100 24.080 115.500 ;
      RECT 27.160 2.100 27.440 115.500 ;
      RECT 30.520 2.100 30.800 115.500 ;
      RECT 33.880 2.100 34.160 115.500 ;
      RECT 37.240 2.100 37.520 115.500 ;
      RECT 40.600 2.100 40.880 115.500 ;
      RECT 43.960 2.100 44.240 115.500 ;
      RECT 47.320 2.100 47.600 115.500 ;
      RECT 50.680 2.100 50.960 115.500 ;
      RECT 54.040 2.100 54.320 115.500 ;
      RECT 57.400 2.100 57.680 115.500 ;
      RECT 60.760 2.100 61.040 115.500 ;
      RECT 64.120 2.100 64.400 115.500 ;
      RECT 67.480 2.100 67.760 115.500 ;
      RECT 70.840 2.100 71.120 115.500 ;
      RECT 74.200 2.100 74.480 115.500 ;
      RECT 77.560 2.100 77.840 115.500 ;
      RECT 80.920 2.100 81.200 115.500 ;
      RECT 84.280 2.100 84.560 115.500 ;
      RECT 87.640 2.100 87.920 115.500 ;
      RECT 91.000 2.100 91.280 115.500 ;
      RECT 94.360 2.100 94.640 115.500 ;
      RECT 97.720 2.100 98.000 115.500 ;
      RECT 101.080 2.100 101.360 115.500 ;
      RECT 104.440 2.100 104.720 115.500 ;
      RECT 107.800 2.100 108.080 115.500 ;
      RECT 111.160 2.100 111.440 115.500 ;
      RECT 114.520 2.100 114.800 115.500 ;
      RECT 117.880 2.100 118.160 115.500 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 121.030 117.600 ;
    LAYER metal2 ;
    RECT 0 0 121.030 117.600 ;
    LAYER metal3 ;
    RECT 0.070 0 121.030 117.600 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.275 ;
    RECT 0 2.345 0.070 2.485 ;
    RECT 0 2.555 0.070 2.695 ;
    RECT 0 2.765 0.070 2.905 ;
    RECT 0 2.975 0.070 3.115 ;
    RECT 0 3.185 0.070 3.325 ;
    RECT 0 3.395 0.070 3.535 ;
    RECT 0 3.605 0.070 3.745 ;
    RECT 0 3.815 0.070 3.955 ;
    RECT 0 4.025 0.070 4.165 ;
    RECT 0 4.235 0.070 4.375 ;
    RECT 0 4.445 0.070 4.585 ;
    RECT 0 4.655 0.070 4.795 ;
    RECT 0 4.865 0.070 5.005 ;
    RECT 0 5.075 0.070 5.215 ;
    RECT 0 5.285 0.070 5.425 ;
    RECT 0 5.495 0.070 5.635 ;
    RECT 0 5.705 0.070 5.845 ;
    RECT 0 5.915 0.070 6.055 ;
    RECT 0 6.125 0.070 6.265 ;
    RECT 0 6.335 0.070 6.475 ;
    RECT 0 6.545 0.070 6.685 ;
    RECT 0 6.755 0.070 6.895 ;
    RECT 0 6.965 0.070 7.105 ;
    RECT 0 7.175 0.070 7.315 ;
    RECT 0 7.385 0.070 7.525 ;
    RECT 0 7.595 0.070 7.735 ;
    RECT 0 7.805 0.070 7.945 ;
    RECT 0 8.015 0.070 8.155 ;
    RECT 0 8.225 0.070 8.365 ;
    RECT 0 8.435 0.070 8.575 ;
    RECT 0 8.645 0.070 8.785 ;
    RECT 0 8.855 0.070 8.995 ;
    RECT 0 9.065 0.070 9.205 ;
    RECT 0 9.275 0.070 9.415 ;
    RECT 0 9.485 0.070 9.625 ;
    RECT 0 9.695 0.070 9.835 ;
    RECT 0 9.905 0.070 10.045 ;
    RECT 0 10.115 0.070 10.255 ;
    RECT 0 10.325 0.070 10.465 ;
    RECT 0 10.535 0.070 10.675 ;
    RECT 0 10.745 0.070 10.885 ;
    RECT 0 10.955 0.070 11.095 ;
    RECT 0 11.165 0.070 11.305 ;
    RECT 0 11.375 0.070 11.515 ;
    RECT 0 11.585 0.070 11.725 ;
    RECT 0 11.795 0.070 11.935 ;
    RECT 0 12.005 0.070 12.145 ;
    RECT 0 12.215 0.070 12.355 ;
    RECT 0 12.425 0.070 12.565 ;
    RECT 0 12.635 0.070 12.775 ;
    RECT 0 12.845 0.070 12.985 ;
    RECT 0 13.055 0.070 13.195 ;
    RECT 0 13.265 0.070 13.405 ;
    RECT 0 13.475 0.070 13.615 ;
    RECT 0 13.685 0.070 13.825 ;
    RECT 0 13.895 0.070 14.035 ;
    RECT 0 14.105 0.070 14.245 ;
    RECT 0 14.315 0.070 14.455 ;
    RECT 0 14.525 0.070 14.665 ;
    RECT 0 14.735 0.070 14.875 ;
    RECT 0 14.945 0.070 15.085 ;
    RECT 0 15.155 0.070 15.295 ;
    RECT 0 15.365 0.070 15.505 ;
    RECT 0 15.575 0.070 15.715 ;
    RECT 0 15.785 0.070 15.925 ;
    RECT 0 15.995 0.070 16.135 ;
    RECT 0 16.205 0.070 16.345 ;
    RECT 0 16.415 0.070 16.555 ;
    RECT 0 16.625 0.070 16.765 ;
    RECT 0 16.835 0.070 16.975 ;
    RECT 0 17.045 0.070 17.185 ;
    RECT 0 17.255 0.070 17.395 ;
    RECT 0 17.465 0.070 17.605 ;
    RECT 0 17.675 0.070 17.815 ;
    RECT 0 17.885 0.070 18.025 ;
    RECT 0 18.095 0.070 18.235 ;
    RECT 0 18.305 0.070 18.445 ;
    RECT 0 18.515 0.070 18.655 ;
    RECT 0 18.725 0.070 18.865 ;
    RECT 0 18.935 0.070 19.075 ;
    RECT 0 19.145 0.070 19.285 ;
    RECT 0 19.355 0.070 19.495 ;
    RECT 0 19.565 0.070 19.705 ;
    RECT 0 19.775 0.070 19.915 ;
    RECT 0 19.985 0.070 20.125 ;
    RECT 0 20.195 0.070 20.335 ;
    RECT 0 20.405 0.070 20.545 ;
    RECT 0 20.615 0.070 20.755 ;
    RECT 0 20.825 0.070 20.965 ;
    RECT 0 21.035 0.070 21.175 ;
    RECT 0 21.245 0.070 21.385 ;
    RECT 0 21.455 0.070 21.595 ;
    RECT 0 21.665 0.070 21.805 ;
    RECT 0 21.875 0.070 22.015 ;
    RECT 0 22.085 0.070 22.225 ;
    RECT 0 22.295 0.070 22.435 ;
    RECT 0 22.505 0.070 22.645 ;
    RECT 0 22.715 0.070 22.855 ;
    RECT 0 22.925 0.070 23.065 ;
    RECT 0 23.135 0.070 23.275 ;
    RECT 0 23.345 0.070 23.485 ;
    RECT 0 23.555 0.070 23.695 ;
    RECT 0 23.765 0.070 23.905 ;
    RECT 0 23.975 0.070 24.115 ;
    RECT 0 24.185 0.070 24.325 ;
    RECT 0 24.395 0.070 24.535 ;
    RECT 0 24.605 0.070 24.745 ;
    RECT 0 24.815 0.070 24.955 ;
    RECT 0 25.025 0.070 25.165 ;
    RECT 0 25.235 0.070 25.375 ;
    RECT 0 25.445 0.070 25.585 ;
    RECT 0 25.655 0.070 25.795 ;
    RECT 0 25.865 0.070 26.005 ;
    RECT 0 26.075 0.070 26.215 ;
    RECT 0 26.285 0.070 35.665 ;
    RECT 0 35.735 0.070 35.875 ;
    RECT 0 35.945 0.070 36.085 ;
    RECT 0 36.155 0.070 36.295 ;
    RECT 0 36.365 0.070 36.505 ;
    RECT 0 36.575 0.070 36.715 ;
    RECT 0 36.785 0.070 36.925 ;
    RECT 0 36.995 0.070 37.135 ;
    RECT 0 37.205 0.070 37.345 ;
    RECT 0 37.415 0.070 37.555 ;
    RECT 0 37.625 0.070 37.765 ;
    RECT 0 37.835 0.070 37.975 ;
    RECT 0 38.045 0.070 38.185 ;
    RECT 0 38.255 0.070 38.395 ;
    RECT 0 38.465 0.070 38.605 ;
    RECT 0 38.675 0.070 38.815 ;
    RECT 0 38.885 0.070 39.025 ;
    RECT 0 39.095 0.070 39.235 ;
    RECT 0 39.305 0.070 39.445 ;
    RECT 0 39.515 0.070 39.655 ;
    RECT 0 39.725 0.070 39.865 ;
    RECT 0 39.935 0.070 40.075 ;
    RECT 0 40.145 0.070 40.285 ;
    RECT 0 40.355 0.070 40.495 ;
    RECT 0 40.565 0.070 40.705 ;
    RECT 0 40.775 0.070 40.915 ;
    RECT 0 40.985 0.070 41.125 ;
    RECT 0 41.195 0.070 41.335 ;
    RECT 0 41.405 0.070 41.545 ;
    RECT 0 41.615 0.070 41.755 ;
    RECT 0 41.825 0.070 41.965 ;
    RECT 0 42.035 0.070 42.175 ;
    RECT 0 42.245 0.070 42.385 ;
    RECT 0 42.455 0.070 42.595 ;
    RECT 0 42.665 0.070 42.805 ;
    RECT 0 42.875 0.070 43.015 ;
    RECT 0 43.085 0.070 43.225 ;
    RECT 0 43.295 0.070 43.435 ;
    RECT 0 43.505 0.070 43.645 ;
    RECT 0 43.715 0.070 43.855 ;
    RECT 0 43.925 0.070 44.065 ;
    RECT 0 44.135 0.070 44.275 ;
    RECT 0 44.345 0.070 44.485 ;
    RECT 0 44.555 0.070 44.695 ;
    RECT 0 44.765 0.070 44.905 ;
    RECT 0 44.975 0.070 45.115 ;
    RECT 0 45.185 0.070 45.325 ;
    RECT 0 45.395 0.070 45.535 ;
    RECT 0 45.605 0.070 45.745 ;
    RECT 0 45.815 0.070 45.955 ;
    RECT 0 46.025 0.070 46.165 ;
    RECT 0 46.235 0.070 46.375 ;
    RECT 0 46.445 0.070 46.585 ;
    RECT 0 46.655 0.070 46.795 ;
    RECT 0 46.865 0.070 47.005 ;
    RECT 0 47.075 0.070 47.215 ;
    RECT 0 47.285 0.070 47.425 ;
    RECT 0 47.495 0.070 47.635 ;
    RECT 0 47.705 0.070 47.845 ;
    RECT 0 47.915 0.070 48.055 ;
    RECT 0 48.125 0.070 48.265 ;
    RECT 0 48.335 0.070 48.475 ;
    RECT 0 48.545 0.070 48.685 ;
    RECT 0 48.755 0.070 48.895 ;
    RECT 0 48.965 0.070 49.105 ;
    RECT 0 49.175 0.070 49.315 ;
    RECT 0 49.385 0.070 49.525 ;
    RECT 0 49.595 0.070 49.735 ;
    RECT 0 49.805 0.070 49.945 ;
    RECT 0 50.015 0.070 50.155 ;
    RECT 0 50.225 0.070 50.365 ;
    RECT 0 50.435 0.070 50.575 ;
    RECT 0 50.645 0.070 50.785 ;
    RECT 0 50.855 0.070 50.995 ;
    RECT 0 51.065 0.070 51.205 ;
    RECT 0 51.275 0.070 51.415 ;
    RECT 0 51.485 0.070 51.625 ;
    RECT 0 51.695 0.070 51.835 ;
    RECT 0 51.905 0.070 52.045 ;
    RECT 0 52.115 0.070 52.255 ;
    RECT 0 52.325 0.070 52.465 ;
    RECT 0 52.535 0.070 52.675 ;
    RECT 0 52.745 0.070 52.885 ;
    RECT 0 52.955 0.070 53.095 ;
    RECT 0 53.165 0.070 53.305 ;
    RECT 0 53.375 0.070 53.515 ;
    RECT 0 53.585 0.070 53.725 ;
    RECT 0 53.795 0.070 53.935 ;
    RECT 0 54.005 0.070 54.145 ;
    RECT 0 54.215 0.070 54.355 ;
    RECT 0 54.425 0.070 54.565 ;
    RECT 0 54.635 0.070 54.775 ;
    RECT 0 54.845 0.070 54.985 ;
    RECT 0 55.055 0.070 55.195 ;
    RECT 0 55.265 0.070 55.405 ;
    RECT 0 55.475 0.070 55.615 ;
    RECT 0 55.685 0.070 55.825 ;
    RECT 0 55.895 0.070 56.035 ;
    RECT 0 56.105 0.070 56.245 ;
    RECT 0 56.315 0.070 56.455 ;
    RECT 0 56.525 0.070 56.665 ;
    RECT 0 56.735 0.070 56.875 ;
    RECT 0 56.945 0.070 57.085 ;
    RECT 0 57.155 0.070 57.295 ;
    RECT 0 57.365 0.070 57.505 ;
    RECT 0 57.575 0.070 57.715 ;
    RECT 0 57.785 0.070 57.925 ;
    RECT 0 57.995 0.070 58.135 ;
    RECT 0 58.205 0.070 58.345 ;
    RECT 0 58.415 0.070 58.555 ;
    RECT 0 58.625 0.070 58.765 ;
    RECT 0 58.835 0.070 58.975 ;
    RECT 0 59.045 0.070 59.185 ;
    RECT 0 59.255 0.070 59.395 ;
    RECT 0 59.465 0.070 59.605 ;
    RECT 0 59.675 0.070 59.815 ;
    RECT 0 59.885 0.070 69.265 ;
    RECT 0 69.335 0.070 69.475 ;
    RECT 0 69.545 0.070 69.685 ;
    RECT 0 69.755 0.070 69.895 ;
    RECT 0 69.965 0.070 70.105 ;
    RECT 0 70.175 0.070 70.315 ;
    RECT 0 70.385 0.070 70.525 ;
    RECT 0 70.595 0.070 70.735 ;
    RECT 0 70.805 0.070 70.945 ;
    RECT 0 71.015 0.070 71.155 ;
    RECT 0 71.225 0.070 71.365 ;
    RECT 0 71.435 0.070 71.575 ;
    RECT 0 71.645 0.070 71.785 ;
    RECT 0 71.855 0.070 71.995 ;
    RECT 0 72.065 0.070 72.205 ;
    RECT 0 72.275 0.070 72.415 ;
    RECT 0 72.485 0.070 72.625 ;
    RECT 0 72.695 0.070 72.835 ;
    RECT 0 72.905 0.070 73.045 ;
    RECT 0 73.115 0.070 73.255 ;
    RECT 0 73.325 0.070 73.465 ;
    RECT 0 73.535 0.070 73.675 ;
    RECT 0 73.745 0.070 73.885 ;
    RECT 0 73.955 0.070 74.095 ;
    RECT 0 74.165 0.070 74.305 ;
    RECT 0 74.375 0.070 74.515 ;
    RECT 0 74.585 0.070 74.725 ;
    RECT 0 74.795 0.070 74.935 ;
    RECT 0 75.005 0.070 75.145 ;
    RECT 0 75.215 0.070 75.355 ;
    RECT 0 75.425 0.070 75.565 ;
    RECT 0 75.635 0.070 75.775 ;
    RECT 0 75.845 0.070 75.985 ;
    RECT 0 76.055 0.070 76.195 ;
    RECT 0 76.265 0.070 76.405 ;
    RECT 0 76.475 0.070 76.615 ;
    RECT 0 76.685 0.070 76.825 ;
    RECT 0 76.895 0.070 77.035 ;
    RECT 0 77.105 0.070 77.245 ;
    RECT 0 77.315 0.070 77.455 ;
    RECT 0 77.525 0.070 77.665 ;
    RECT 0 77.735 0.070 77.875 ;
    RECT 0 77.945 0.070 78.085 ;
    RECT 0 78.155 0.070 78.295 ;
    RECT 0 78.365 0.070 78.505 ;
    RECT 0 78.575 0.070 78.715 ;
    RECT 0 78.785 0.070 78.925 ;
    RECT 0 78.995 0.070 79.135 ;
    RECT 0 79.205 0.070 79.345 ;
    RECT 0 79.415 0.070 79.555 ;
    RECT 0 79.625 0.070 79.765 ;
    RECT 0 79.835 0.070 79.975 ;
    RECT 0 80.045 0.070 80.185 ;
    RECT 0 80.255 0.070 80.395 ;
    RECT 0 80.465 0.070 80.605 ;
    RECT 0 80.675 0.070 80.815 ;
    RECT 0 80.885 0.070 81.025 ;
    RECT 0 81.095 0.070 81.235 ;
    RECT 0 81.305 0.070 81.445 ;
    RECT 0 81.515 0.070 81.655 ;
    RECT 0 81.725 0.070 81.865 ;
    RECT 0 81.935 0.070 82.075 ;
    RECT 0 82.145 0.070 82.285 ;
    RECT 0 82.355 0.070 82.495 ;
    RECT 0 82.565 0.070 82.705 ;
    RECT 0 82.775 0.070 82.915 ;
    RECT 0 82.985 0.070 83.125 ;
    RECT 0 83.195 0.070 83.335 ;
    RECT 0 83.405 0.070 83.545 ;
    RECT 0 83.615 0.070 83.755 ;
    RECT 0 83.825 0.070 83.965 ;
    RECT 0 84.035 0.070 84.175 ;
    RECT 0 84.245 0.070 84.385 ;
    RECT 0 84.455 0.070 84.595 ;
    RECT 0 84.665 0.070 84.805 ;
    RECT 0 84.875 0.070 85.015 ;
    RECT 0 85.085 0.070 85.225 ;
    RECT 0 85.295 0.070 85.435 ;
    RECT 0 85.505 0.070 85.645 ;
    RECT 0 85.715 0.070 85.855 ;
    RECT 0 85.925 0.070 86.065 ;
    RECT 0 86.135 0.070 86.275 ;
    RECT 0 86.345 0.070 86.485 ;
    RECT 0 86.555 0.070 86.695 ;
    RECT 0 86.765 0.070 86.905 ;
    RECT 0 86.975 0.070 87.115 ;
    RECT 0 87.185 0.070 87.325 ;
    RECT 0 87.395 0.070 87.535 ;
    RECT 0 87.605 0.070 87.745 ;
    RECT 0 87.815 0.070 87.955 ;
    RECT 0 88.025 0.070 88.165 ;
    RECT 0 88.235 0.070 88.375 ;
    RECT 0 88.445 0.070 88.585 ;
    RECT 0 88.655 0.070 88.795 ;
    RECT 0 88.865 0.070 89.005 ;
    RECT 0 89.075 0.070 89.215 ;
    RECT 0 89.285 0.070 89.425 ;
    RECT 0 89.495 0.070 89.635 ;
    RECT 0 89.705 0.070 89.845 ;
    RECT 0 89.915 0.070 90.055 ;
    RECT 0 90.125 0.070 90.265 ;
    RECT 0 90.335 0.070 90.475 ;
    RECT 0 90.545 0.070 90.685 ;
    RECT 0 90.755 0.070 90.895 ;
    RECT 0 90.965 0.070 91.105 ;
    RECT 0 91.175 0.070 91.315 ;
    RECT 0 91.385 0.070 91.525 ;
    RECT 0 91.595 0.070 91.735 ;
    RECT 0 91.805 0.070 91.945 ;
    RECT 0 92.015 0.070 92.155 ;
    RECT 0 92.225 0.070 92.365 ;
    RECT 0 92.435 0.070 92.575 ;
    RECT 0 92.645 0.070 92.785 ;
    RECT 0 92.855 0.070 92.995 ;
    RECT 0 93.065 0.070 93.205 ;
    RECT 0 93.275 0.070 93.415 ;
    RECT 0 93.485 0.070 102.865 ;
    RECT 0 102.935 0.070 103.075 ;
    RECT 0 103.145 0.070 103.285 ;
    RECT 0 103.355 0.070 103.495 ;
    RECT 0 103.565 0.070 103.705 ;
    RECT 0 103.775 0.070 103.915 ;
    RECT 0 103.985 0.070 104.125 ;
    RECT 0 104.195 0.070 113.575 ;
    RECT 0 113.645 0.070 113.785 ;
    RECT 0 113.855 0.070 113.995 ;
    RECT 0 114.065 0.070 117.600 ;
    LAYER metal4 ;
    RECT 0 0 121.030 2.100 ;
    RECT 0 115.500 121.030 117.600 ;
    RECT 0.000 2.100 1.960 115.500 ;
    RECT 2.240 2.100 3.640 115.500 ;
    RECT 3.920 2.100 5.320 115.500 ;
    RECT 5.600 2.100 7.000 115.500 ;
    RECT 7.280 2.100 8.680 115.500 ;
    RECT 8.960 2.100 10.360 115.500 ;
    RECT 10.640 2.100 12.040 115.500 ;
    RECT 12.320 2.100 13.720 115.500 ;
    RECT 14.000 2.100 15.400 115.500 ;
    RECT 15.680 2.100 17.080 115.500 ;
    RECT 17.360 2.100 18.760 115.500 ;
    RECT 19.040 2.100 20.440 115.500 ;
    RECT 20.720 2.100 22.120 115.500 ;
    RECT 22.400 2.100 23.800 115.500 ;
    RECT 24.080 2.100 25.480 115.500 ;
    RECT 25.760 2.100 27.160 115.500 ;
    RECT 27.440 2.100 28.840 115.500 ;
    RECT 29.120 2.100 30.520 115.500 ;
    RECT 30.800 2.100 32.200 115.500 ;
    RECT 32.480 2.100 33.880 115.500 ;
    RECT 34.160 2.100 35.560 115.500 ;
    RECT 35.840 2.100 37.240 115.500 ;
    RECT 37.520 2.100 38.920 115.500 ;
    RECT 39.200 2.100 40.600 115.500 ;
    RECT 40.880 2.100 42.280 115.500 ;
    RECT 42.560 2.100 43.960 115.500 ;
    RECT 44.240 2.100 45.640 115.500 ;
    RECT 45.920 2.100 47.320 115.500 ;
    RECT 47.600 2.100 49.000 115.500 ;
    RECT 49.280 2.100 50.680 115.500 ;
    RECT 50.960 2.100 52.360 115.500 ;
    RECT 52.640 2.100 54.040 115.500 ;
    RECT 54.320 2.100 55.720 115.500 ;
    RECT 56.000 2.100 57.400 115.500 ;
    RECT 57.680 2.100 59.080 115.500 ;
    RECT 59.360 2.100 60.760 115.500 ;
    RECT 61.040 2.100 62.440 115.500 ;
    RECT 62.720 2.100 64.120 115.500 ;
    RECT 64.400 2.100 65.800 115.500 ;
    RECT 66.080 2.100 67.480 115.500 ;
    RECT 67.760 2.100 69.160 115.500 ;
    RECT 69.440 2.100 70.840 115.500 ;
    RECT 71.120 2.100 72.520 115.500 ;
    RECT 72.800 2.100 74.200 115.500 ;
    RECT 74.480 2.100 75.880 115.500 ;
    RECT 76.160 2.100 77.560 115.500 ;
    RECT 77.840 2.100 79.240 115.500 ;
    RECT 79.520 2.100 80.920 115.500 ;
    RECT 81.200 2.100 82.600 115.500 ;
    RECT 82.880 2.100 84.280 115.500 ;
    RECT 84.560 2.100 85.960 115.500 ;
    RECT 86.240 2.100 87.640 115.500 ;
    RECT 87.920 2.100 89.320 115.500 ;
    RECT 89.600 2.100 91.000 115.500 ;
    RECT 91.280 2.100 92.680 115.500 ;
    RECT 92.960 2.100 94.360 115.500 ;
    RECT 94.640 2.100 96.040 115.500 ;
    RECT 96.320 2.100 97.720 115.500 ;
    RECT 98.000 2.100 99.400 115.500 ;
    RECT 99.680 2.100 101.080 115.500 ;
    RECT 101.360 2.100 102.760 115.500 ;
    RECT 103.040 2.100 104.440 115.500 ;
    RECT 104.720 2.100 106.120 115.500 ;
    RECT 106.400 2.100 107.800 115.500 ;
    RECT 108.080 2.100 109.480 115.500 ;
    RECT 109.760 2.100 111.160 115.500 ;
    RECT 111.440 2.100 112.840 115.500 ;
    RECT 113.120 2.100 114.520 115.500 ;
    RECT 114.800 2.100 116.200 115.500 ;
    RECT 116.480 2.100 117.880 115.500 ;
    RECT 118.160 2.100 121.030 115.500 ;
    LAYER OVERLAP ;
    RECT 0 0 121.030 117.600 ;
  END
END fakeram45_128x116

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_128x32
  FOREIGN fakeram45_128x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 59.660 BY 82.600 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.695 0.070 2.765 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.955 0.070 4.025 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.215 0.070 5.285 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.475 0.070 6.545 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.735 0.070 7.805 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.995 0.070 9.065 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.255 0.070 10.325 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.515 0.070 11.585 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.775 0.070 12.845 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.035 0.070 14.105 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.295 0.070 15.365 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.555 0.070 16.625 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.185 0.070 17.255 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.815 0.070 17.885 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.075 0.070 19.145 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.335 0.070 20.405 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.595 0.070 21.665 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.955 0.070 25.025 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.215 0.070 26.285 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.475 0.070 27.545 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.105 0.070 28.175 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.735 0.070 28.805 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.995 0.070 30.065 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.625 0.070 30.695 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.255 0.070 31.325 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.885 0.070 31.955 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.515 0.070 32.585 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.145 0.070 33.215 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.775 0.070 33.845 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.035 0.070 35.105 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.295 0.070 36.365 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.555 0.070 37.625 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.185 0.070 38.255 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.815 0.070 38.885 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.075 0.070 40.145 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.335 0.070 41.405 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.595 0.070 42.665 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.855 0.070 43.925 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.585 0.070 46.655 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.215 0.070 47.285 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.475 0.070 48.545 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.735 0.070 49.805 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.995 0.070 51.065 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.625 0.070 51.695 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.255 0.070 52.325 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.515 0.070 53.585 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.145 0.070 54.215 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.775 0.070 54.845 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.035 0.070 56.105 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.665 0.070 56.735 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.295 0.070 57.365 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.555 0.070 58.625 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.185 0.070 59.255 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.815 0.070 59.885 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.445 0.070 60.515 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.075 0.070 61.145 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.705 0.070 61.775 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.335 0.070 62.405 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.965 0.070 63.035 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.595 0.070 63.665 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.225 0.070 64.295 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.855 0.070 64.925 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.485 0.070 65.555 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.115 0.070 66.185 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.845 0.070 68.915 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.475 0.070 69.545 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.105 0.070 70.175 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.735 0.070 70.805 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.995 0.070 72.065 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.625 0.070 72.695 ;
    END
  END addr_in[6]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.355 0.070 75.425 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.615 0.070 76.685 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 80.500 ;
      RECT 5.320 2.100 5.600 80.500 ;
      RECT 8.680 2.100 8.960 80.500 ;
      RECT 12.040 2.100 12.320 80.500 ;
      RECT 15.400 2.100 15.680 80.500 ;
      RECT 18.760 2.100 19.040 80.500 ;
      RECT 22.120 2.100 22.400 80.500 ;
      RECT 25.480 2.100 25.760 80.500 ;
      RECT 28.840 2.100 29.120 80.500 ;
      RECT 32.200 2.100 32.480 80.500 ;
      RECT 35.560 2.100 35.840 80.500 ;
      RECT 38.920 2.100 39.200 80.500 ;
      RECT 42.280 2.100 42.560 80.500 ;
      RECT 45.640 2.100 45.920 80.500 ;
      RECT 49.000 2.100 49.280 80.500 ;
      RECT 52.360 2.100 52.640 80.500 ;
      RECT 55.720 2.100 56.000 80.500 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 80.500 ;
      RECT 7.000 2.100 7.280 80.500 ;
      RECT 10.360 2.100 10.640 80.500 ;
      RECT 13.720 2.100 14.000 80.500 ;
      RECT 17.080 2.100 17.360 80.500 ;
      RECT 20.440 2.100 20.720 80.500 ;
      RECT 23.800 2.100 24.080 80.500 ;
      RECT 27.160 2.100 27.440 80.500 ;
      RECT 30.520 2.100 30.800 80.500 ;
      RECT 33.880 2.100 34.160 80.500 ;
      RECT 37.240 2.100 37.520 80.500 ;
      RECT 40.600 2.100 40.880 80.500 ;
      RECT 43.960 2.100 44.240 80.500 ;
      RECT 47.320 2.100 47.600 80.500 ;
      RECT 50.680 2.100 50.960 80.500 ;
      RECT 54.040 2.100 54.320 80.500 ;
      RECT 57.400 2.100 57.680 80.500 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 59.660 82.600 ;
    LAYER metal2 ;
    RECT 0 0 59.660 82.600 ;
    LAYER metal3 ;
    RECT 0.070 0 59.660 82.600 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.695 ;
    RECT 0 2.765 0.070 3.325 ;
    RECT 0 3.395 0.070 3.955 ;
    RECT 0 4.025 0.070 4.585 ;
    RECT 0 4.655 0.070 5.215 ;
    RECT 0 5.285 0.070 5.845 ;
    RECT 0 5.915 0.070 6.475 ;
    RECT 0 6.545 0.070 7.105 ;
    RECT 0 7.175 0.070 7.735 ;
    RECT 0 7.805 0.070 8.365 ;
    RECT 0 8.435 0.070 8.995 ;
    RECT 0 9.065 0.070 9.625 ;
    RECT 0 9.695 0.070 10.255 ;
    RECT 0 10.325 0.070 10.885 ;
    RECT 0 10.955 0.070 11.515 ;
    RECT 0 11.585 0.070 12.145 ;
    RECT 0 12.215 0.070 12.775 ;
    RECT 0 12.845 0.070 13.405 ;
    RECT 0 13.475 0.070 14.035 ;
    RECT 0 14.105 0.070 14.665 ;
    RECT 0 14.735 0.070 15.295 ;
    RECT 0 15.365 0.070 15.925 ;
    RECT 0 15.995 0.070 16.555 ;
    RECT 0 16.625 0.070 17.185 ;
    RECT 0 17.255 0.070 17.815 ;
    RECT 0 17.885 0.070 18.445 ;
    RECT 0 18.515 0.070 19.075 ;
    RECT 0 19.145 0.070 19.705 ;
    RECT 0 19.775 0.070 20.335 ;
    RECT 0 20.405 0.070 20.965 ;
    RECT 0 21.035 0.070 21.595 ;
    RECT 0 21.665 0.070 24.325 ;
    RECT 0 24.395 0.070 24.955 ;
    RECT 0 25.025 0.070 25.585 ;
    RECT 0 25.655 0.070 26.215 ;
    RECT 0 26.285 0.070 26.845 ;
    RECT 0 26.915 0.070 27.475 ;
    RECT 0 27.545 0.070 28.105 ;
    RECT 0 28.175 0.070 28.735 ;
    RECT 0 28.805 0.070 29.365 ;
    RECT 0 29.435 0.070 29.995 ;
    RECT 0 30.065 0.070 30.625 ;
    RECT 0 30.695 0.070 31.255 ;
    RECT 0 31.325 0.070 31.885 ;
    RECT 0 31.955 0.070 32.515 ;
    RECT 0 32.585 0.070 33.145 ;
    RECT 0 33.215 0.070 33.775 ;
    RECT 0 33.845 0.070 34.405 ;
    RECT 0 34.475 0.070 35.035 ;
    RECT 0 35.105 0.070 35.665 ;
    RECT 0 35.735 0.070 36.295 ;
    RECT 0 36.365 0.070 36.925 ;
    RECT 0 36.995 0.070 37.555 ;
    RECT 0 37.625 0.070 38.185 ;
    RECT 0 38.255 0.070 38.815 ;
    RECT 0 38.885 0.070 39.445 ;
    RECT 0 39.515 0.070 40.075 ;
    RECT 0 40.145 0.070 40.705 ;
    RECT 0 40.775 0.070 41.335 ;
    RECT 0 41.405 0.070 41.965 ;
    RECT 0 42.035 0.070 42.595 ;
    RECT 0 42.665 0.070 43.225 ;
    RECT 0 43.295 0.070 43.855 ;
    RECT 0 43.925 0.070 46.585 ;
    RECT 0 46.655 0.070 47.215 ;
    RECT 0 47.285 0.070 47.845 ;
    RECT 0 47.915 0.070 48.475 ;
    RECT 0 48.545 0.070 49.105 ;
    RECT 0 49.175 0.070 49.735 ;
    RECT 0 49.805 0.070 50.365 ;
    RECT 0 50.435 0.070 50.995 ;
    RECT 0 51.065 0.070 51.625 ;
    RECT 0 51.695 0.070 52.255 ;
    RECT 0 52.325 0.070 52.885 ;
    RECT 0 52.955 0.070 53.515 ;
    RECT 0 53.585 0.070 54.145 ;
    RECT 0 54.215 0.070 54.775 ;
    RECT 0 54.845 0.070 55.405 ;
    RECT 0 55.475 0.070 56.035 ;
    RECT 0 56.105 0.070 56.665 ;
    RECT 0 56.735 0.070 57.295 ;
    RECT 0 57.365 0.070 57.925 ;
    RECT 0 57.995 0.070 58.555 ;
    RECT 0 58.625 0.070 59.185 ;
    RECT 0 59.255 0.070 59.815 ;
    RECT 0 59.885 0.070 60.445 ;
    RECT 0 60.515 0.070 61.075 ;
    RECT 0 61.145 0.070 61.705 ;
    RECT 0 61.775 0.070 62.335 ;
    RECT 0 62.405 0.070 62.965 ;
    RECT 0 63.035 0.070 63.595 ;
    RECT 0 63.665 0.070 64.225 ;
    RECT 0 64.295 0.070 64.855 ;
    RECT 0 64.925 0.070 65.485 ;
    RECT 0 65.555 0.070 66.115 ;
    RECT 0 66.185 0.070 68.845 ;
    RECT 0 68.915 0.070 69.475 ;
    RECT 0 69.545 0.070 70.105 ;
    RECT 0 70.175 0.070 70.735 ;
    RECT 0 70.805 0.070 71.365 ;
    RECT 0 71.435 0.070 71.995 ;
    RECT 0 72.065 0.070 72.625 ;
    RECT 0 72.695 0.070 75.355 ;
    RECT 0 75.425 0.070 75.985 ;
    RECT 0 76.055 0.070 76.615 ;
    RECT 0 76.685 0.070 82.600 ;
    LAYER metal4 ;
    RECT 0 0 59.660 2.100 ;
    RECT 0 80.500 59.660 82.600 ;
    RECT 0.000 2.100 1.960 80.500 ;
    RECT 2.240 2.100 3.640 80.500 ;
    RECT 3.920 2.100 5.320 80.500 ;
    RECT 5.600 2.100 7.000 80.500 ;
    RECT 7.280 2.100 8.680 80.500 ;
    RECT 8.960 2.100 10.360 80.500 ;
    RECT 10.640 2.100 12.040 80.500 ;
    RECT 12.320 2.100 13.720 80.500 ;
    RECT 14.000 2.100 15.400 80.500 ;
    RECT 15.680 2.100 17.080 80.500 ;
    RECT 17.360 2.100 18.760 80.500 ;
    RECT 19.040 2.100 20.440 80.500 ;
    RECT 20.720 2.100 22.120 80.500 ;
    RECT 22.400 2.100 23.800 80.500 ;
    RECT 24.080 2.100 25.480 80.500 ;
    RECT 25.760 2.100 27.160 80.500 ;
    RECT 27.440 2.100 28.840 80.500 ;
    RECT 29.120 2.100 30.520 80.500 ;
    RECT 30.800 2.100 32.200 80.500 ;
    RECT 32.480 2.100 33.880 80.500 ;
    RECT 34.160 2.100 35.560 80.500 ;
    RECT 35.840 2.100 37.240 80.500 ;
    RECT 37.520 2.100 38.920 80.500 ;
    RECT 39.200 2.100 40.600 80.500 ;
    RECT 40.880 2.100 42.280 80.500 ;
    RECT 42.560 2.100 43.960 80.500 ;
    RECT 44.240 2.100 45.640 80.500 ;
    RECT 45.920 2.100 47.320 80.500 ;
    RECT 47.600 2.100 49.000 80.500 ;
    RECT 49.280 2.100 50.680 80.500 ;
    RECT 50.960 2.100 52.360 80.500 ;
    RECT 52.640 2.100 54.040 80.500 ;
    RECT 54.320 2.100 55.720 80.500 ;
    RECT 56.000 2.100 57.400 80.500 ;
    RECT 57.680 2.100 59.660 80.500 ;
    LAYER OVERLAP ;
    RECT 0 0 59.660 82.600 ;
  END
END fakeram45_128x32

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_64x124
  FOREIGN fakeram45_64x124 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 80.560 BY 121.800 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.275 0.070 2.345 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.695 0.070 2.765 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.115 0.070 3.185 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.535 0.070 3.605 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.955 0.070 4.025 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.375 0.070 4.445 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.795 0.070 4.865 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.215 0.070 5.285 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.635 0.070 5.705 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.055 0.070 6.125 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.475 0.070 6.545 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.895 0.070 6.965 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.315 0.070 7.385 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.735 0.070 7.805 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.155 0.070 8.225 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.575 0.070 8.645 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.785 0.070 8.855 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.995 0.070 9.065 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.415 0.070 9.485 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.835 0.070 9.905 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.255 0.070 10.325 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.675 0.070 10.745 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.095 0.070 11.165 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.515 0.070 11.585 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.935 0.070 12.005 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.355 0.070 12.425 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.775 0.070 12.845 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.985 0.070 13.055 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.195 0.070 13.265 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.615 0.070 13.685 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.035 0.070 14.105 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.455 0.070 14.525 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.875 0.070 14.945 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.295 0.070 15.365 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.505 0.070 15.575 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.715 0.070 15.785 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.135 0.070 16.205 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.345 0.070 16.415 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.555 0.070 16.625 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.975 0.070 17.045 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.185 0.070 17.255 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.395 0.070 17.465 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.605 0.070 17.675 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.815 0.070 17.885 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.025 0.070 18.095 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.235 0.070 18.305 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.655 0.070 18.725 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.075 0.070 19.145 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.495 0.070 19.565 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.915 0.070 19.985 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.335 0.070 20.405 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.545 0.070 20.615 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.755 0.070 20.825 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.175 0.070 21.245 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.595 0.070 21.665 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.015 0.070 22.085 ;
    END
  END w_mask_in[95]
  PIN w_mask_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.225 0.070 22.295 ;
    END
  END w_mask_in[96]
  PIN w_mask_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.435 0.070 22.505 ;
    END
  END w_mask_in[97]
  PIN w_mask_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END w_mask_in[98]
  PIN w_mask_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.855 0.070 22.925 ;
    END
  END w_mask_in[99]
  PIN w_mask_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END w_mask_in[100]
  PIN w_mask_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.275 0.070 23.345 ;
    END
  END w_mask_in[101]
  PIN w_mask_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END w_mask_in[102]
  PIN w_mask_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.695 0.070 23.765 ;
    END
  END w_mask_in[103]
  PIN w_mask_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.905 0.070 23.975 ;
    END
  END w_mask_in[104]
  PIN w_mask_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.115 0.070 24.185 ;
    END
  END w_mask_in[105]
  PIN w_mask_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END w_mask_in[106]
  PIN w_mask_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.535 0.070 24.605 ;
    END
  END w_mask_in[107]
  PIN w_mask_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END w_mask_in[108]
  PIN w_mask_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.955 0.070 25.025 ;
    END
  END w_mask_in[109]
  PIN w_mask_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END w_mask_in[110]
  PIN w_mask_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.375 0.070 25.445 ;
    END
  END w_mask_in[111]
  PIN w_mask_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END w_mask_in[112]
  PIN w_mask_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.795 0.070 25.865 ;
    END
  END w_mask_in[113]
  PIN w_mask_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END w_mask_in[114]
  PIN w_mask_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.215 0.070 26.285 ;
    END
  END w_mask_in[115]
  PIN w_mask_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.425 0.070 26.495 ;
    END
  END w_mask_in[116]
  PIN w_mask_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.635 0.070 26.705 ;
    END
  END w_mask_in[117]
  PIN w_mask_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END w_mask_in[118]
  PIN w_mask_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.055 0.070 27.125 ;
    END
  END w_mask_in[119]
  PIN w_mask_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END w_mask_in[120]
  PIN w_mask_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.475 0.070 27.545 ;
    END
  END w_mask_in[121]
  PIN w_mask_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.685 0.070 27.755 ;
    END
  END w_mask_in[122]
  PIN w_mask_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.895 0.070 27.965 ;
    END
  END w_mask_in[123]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.135 0.070 37.205 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.555 0.070 37.625 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.975 0.070 38.045 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.185 0.070 38.255 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.395 0.070 38.465 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.815 0.070 38.885 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.235 0.070 39.305 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.655 0.070 39.725 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.075 0.070 40.145 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.495 0.070 40.565 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.915 0.070 40.985 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.335 0.070 41.405 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.755 0.070 41.825 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.175 0.070 42.245 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.595 0.070 42.665 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.015 0.070 43.085 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.435 0.070 43.505 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.855 0.070 43.925 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.275 0.070 44.345 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.695 0.070 44.765 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.115 0.070 45.185 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.325 0.070 45.395 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.535 0.070 45.605 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.745 0.070 45.815 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.955 0.070 46.025 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.375 0.070 46.445 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.585 0.070 46.655 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.795 0.070 46.865 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.215 0.070 47.285 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.635 0.070 47.705 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.055 0.070 48.125 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.265 0.070 48.335 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.475 0.070 48.545 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.895 0.070 48.965 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.315 0.070 49.385 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.735 0.070 49.805 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.945 0.070 50.015 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.155 0.070 50.225 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.575 0.070 50.645 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.785 0.070 50.855 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.995 0.070 51.065 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.205 0.070 51.275 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.415 0.070 51.485 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.625 0.070 51.695 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.835 0.070 51.905 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.045 0.070 52.115 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.255 0.070 52.325 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.675 0.070 52.745 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.095 0.070 53.165 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.305 0.070 53.375 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.515 0.070 53.585 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.935 0.070 54.005 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.145 0.070 54.215 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.355 0.070 54.425 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.775 0.070 54.845 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.985 0.070 55.055 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.195 0.070 55.265 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.615 0.070 55.685 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.825 0.070 55.895 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.035 0.070 56.105 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.455 0.070 56.525 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.665 0.070 56.735 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.875 0.070 56.945 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.085 0.070 57.155 ;
    END
  END rd_out[95]
  PIN rd_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.295 0.070 57.365 ;
    END
  END rd_out[96]
  PIN rd_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.505 0.070 57.575 ;
    END
  END rd_out[97]
  PIN rd_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.715 0.070 57.785 ;
    END
  END rd_out[98]
  PIN rd_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END rd_out[99]
  PIN rd_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.135 0.070 58.205 ;
    END
  END rd_out[100]
  PIN rd_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.345 0.070 58.415 ;
    END
  END rd_out[101]
  PIN rd_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.555 0.070 58.625 ;
    END
  END rd_out[102]
  PIN rd_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.765 0.070 58.835 ;
    END
  END rd_out[103]
  PIN rd_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.975 0.070 59.045 ;
    END
  END rd_out[104]
  PIN rd_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.185 0.070 59.255 ;
    END
  END rd_out[105]
  PIN rd_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.395 0.070 59.465 ;
    END
  END rd_out[106]
  PIN rd_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.605 0.070 59.675 ;
    END
  END rd_out[107]
  PIN rd_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.815 0.070 59.885 ;
    END
  END rd_out[108]
  PIN rd_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.025 0.070 60.095 ;
    END
  END rd_out[109]
  PIN rd_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.235 0.070 60.305 ;
    END
  END rd_out[110]
  PIN rd_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.445 0.070 60.515 ;
    END
  END rd_out[111]
  PIN rd_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.655 0.070 60.725 ;
    END
  END rd_out[112]
  PIN rd_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.865 0.070 60.935 ;
    END
  END rd_out[113]
  PIN rd_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.075 0.070 61.145 ;
    END
  END rd_out[114]
  PIN rd_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.285 0.070 61.355 ;
    END
  END rd_out[115]
  PIN rd_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.495 0.070 61.565 ;
    END
  END rd_out[116]
  PIN rd_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.705 0.070 61.775 ;
    END
  END rd_out[117]
  PIN rd_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.915 0.070 61.985 ;
    END
  END rd_out[118]
  PIN rd_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.125 0.070 62.195 ;
    END
  END rd_out[119]
  PIN rd_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.335 0.070 62.405 ;
    END
  END rd_out[120]
  PIN rd_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.545 0.070 62.615 ;
    END
  END rd_out[121]
  PIN rd_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.755 0.070 62.825 ;
    END
  END rd_out[122]
  PIN rd_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.965 0.070 63.035 ;
    END
  END rd_out[123]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.205 0.070 72.275 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.415 0.070 72.485 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.625 0.070 72.695 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.835 0.070 72.905 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.255 0.070 73.325 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.465 0.070 73.535 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.675 0.070 73.745 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.095 0.070 74.165 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.305 0.070 74.375 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.515 0.070 74.585 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.725 0.070 74.795 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.935 0.070 75.005 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.145 0.070 75.215 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.355 0.070 75.425 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.775 0.070 75.845 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.195 0.070 76.265 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.405 0.070 76.475 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.615 0.070 76.685 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.825 0.070 76.895 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.035 0.070 77.105 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.245 0.070 77.315 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.455 0.070 77.525 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.665 0.070 77.735 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.875 0.070 77.945 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.085 0.070 78.155 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.295 0.070 78.365 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.505 0.070 78.575 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.715 0.070 78.785 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.925 0.070 78.995 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.135 0.070 79.205 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.345 0.070 79.415 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.555 0.070 79.625 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.975 0.070 80.045 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.185 0.070 80.255 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.395 0.070 80.465 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.605 0.070 80.675 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.815 0.070 80.885 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.025 0.070 81.095 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.235 0.070 81.305 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.445 0.070 81.515 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.655 0.070 81.725 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.075 0.070 82.145 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.285 0.070 82.355 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.495 0.070 82.565 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.705 0.070 82.775 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.915 0.070 82.985 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.125 0.070 83.195 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.335 0.070 83.405 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.545 0.070 83.615 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.755 0.070 83.825 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.965 0.070 84.035 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.175 0.070 84.245 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.385 0.070 84.455 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.595 0.070 84.665 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.015 0.070 85.085 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.225 0.070 85.295 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.435 0.070 85.505 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.855 0.070 85.925 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.065 0.070 86.135 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.275 0.070 86.345 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.485 0.070 86.555 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.695 0.070 86.765 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.905 0.070 86.975 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.115 0.070 87.185 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.325 0.070 87.395 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.535 0.070 87.605 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.745 0.070 87.815 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.955 0.070 88.025 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.165 0.070 88.235 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.375 0.070 88.445 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.585 0.070 88.655 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.795 0.070 88.865 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.005 0.070 89.075 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.215 0.070 89.285 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.425 0.070 89.495 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.635 0.070 89.705 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.845 0.070 89.915 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.055 0.070 90.125 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.265 0.070 90.335 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.475 0.070 90.545 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.685 0.070 90.755 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.895 0.070 90.965 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.105 0.070 91.175 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.315 0.070 91.385 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.525 0.070 91.595 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.735 0.070 91.805 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.945 0.070 92.015 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.155 0.070 92.225 ;
    END
  END wd_in[95]
  PIN wd_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.365 0.070 92.435 ;
    END
  END wd_in[96]
  PIN wd_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.575 0.070 92.645 ;
    END
  END wd_in[97]
  PIN wd_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.785 0.070 92.855 ;
    END
  END wd_in[98]
  PIN wd_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.995 0.070 93.065 ;
    END
  END wd_in[99]
  PIN wd_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.205 0.070 93.275 ;
    END
  END wd_in[100]
  PIN wd_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.415 0.070 93.485 ;
    END
  END wd_in[101]
  PIN wd_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.625 0.070 93.695 ;
    END
  END wd_in[102]
  PIN wd_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.835 0.070 93.905 ;
    END
  END wd_in[103]
  PIN wd_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.045 0.070 94.115 ;
    END
  END wd_in[104]
  PIN wd_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.255 0.070 94.325 ;
    END
  END wd_in[105]
  PIN wd_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.465 0.070 94.535 ;
    END
  END wd_in[106]
  PIN wd_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.675 0.070 94.745 ;
    END
  END wd_in[107]
  PIN wd_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.885 0.070 94.955 ;
    END
  END wd_in[108]
  PIN wd_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.095 0.070 95.165 ;
    END
  END wd_in[109]
  PIN wd_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.305 0.070 95.375 ;
    END
  END wd_in[110]
  PIN wd_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.515 0.070 95.585 ;
    END
  END wd_in[111]
  PIN wd_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.725 0.070 95.795 ;
    END
  END wd_in[112]
  PIN wd_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.935 0.070 96.005 ;
    END
  END wd_in[113]
  PIN wd_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.145 0.070 96.215 ;
    END
  END wd_in[114]
  PIN wd_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.355 0.070 96.425 ;
    END
  END wd_in[115]
  PIN wd_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.565 0.070 96.635 ;
    END
  END wd_in[116]
  PIN wd_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.775 0.070 96.845 ;
    END
  END wd_in[117]
  PIN wd_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.985 0.070 97.055 ;
    END
  END wd_in[118]
  PIN wd_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.195 0.070 97.265 ;
    END
  END wd_in[119]
  PIN wd_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.405 0.070 97.475 ;
    END
  END wd_in[120]
  PIN wd_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.615 0.070 97.685 ;
    END
  END wd_in[121]
  PIN wd_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.825 0.070 97.895 ;
    END
  END wd_in[122]
  PIN wd_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.035 0.070 98.105 ;
    END
  END wd_in[123]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.275 0.070 107.345 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.485 0.070 107.555 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.695 0.070 107.765 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.905 0.070 107.975 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.115 0.070 108.185 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.325 0.070 108.395 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.565 0.070 117.635 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.775 0.070 117.845 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.985 0.070 118.055 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 119.700 ;
      RECT 5.320 2.100 5.600 119.700 ;
      RECT 8.680 2.100 8.960 119.700 ;
      RECT 12.040 2.100 12.320 119.700 ;
      RECT 15.400 2.100 15.680 119.700 ;
      RECT 18.760 2.100 19.040 119.700 ;
      RECT 22.120 2.100 22.400 119.700 ;
      RECT 25.480 2.100 25.760 119.700 ;
      RECT 28.840 2.100 29.120 119.700 ;
      RECT 32.200 2.100 32.480 119.700 ;
      RECT 35.560 2.100 35.840 119.700 ;
      RECT 38.920 2.100 39.200 119.700 ;
      RECT 42.280 2.100 42.560 119.700 ;
      RECT 45.640 2.100 45.920 119.700 ;
      RECT 49.000 2.100 49.280 119.700 ;
      RECT 52.360 2.100 52.640 119.700 ;
      RECT 55.720 2.100 56.000 119.700 ;
      RECT 59.080 2.100 59.360 119.700 ;
      RECT 62.440 2.100 62.720 119.700 ;
      RECT 65.800 2.100 66.080 119.700 ;
      RECT 69.160 2.100 69.440 119.700 ;
      RECT 72.520 2.100 72.800 119.700 ;
      RECT 75.880 2.100 76.160 119.700 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 119.700 ;
      RECT 7.000 2.100 7.280 119.700 ;
      RECT 10.360 2.100 10.640 119.700 ;
      RECT 13.720 2.100 14.000 119.700 ;
      RECT 17.080 2.100 17.360 119.700 ;
      RECT 20.440 2.100 20.720 119.700 ;
      RECT 23.800 2.100 24.080 119.700 ;
      RECT 27.160 2.100 27.440 119.700 ;
      RECT 30.520 2.100 30.800 119.700 ;
      RECT 33.880 2.100 34.160 119.700 ;
      RECT 37.240 2.100 37.520 119.700 ;
      RECT 40.600 2.100 40.880 119.700 ;
      RECT 43.960 2.100 44.240 119.700 ;
      RECT 47.320 2.100 47.600 119.700 ;
      RECT 50.680 2.100 50.960 119.700 ;
      RECT 54.040 2.100 54.320 119.700 ;
      RECT 57.400 2.100 57.680 119.700 ;
      RECT 60.760 2.100 61.040 119.700 ;
      RECT 64.120 2.100 64.400 119.700 ;
      RECT 67.480 2.100 67.760 119.700 ;
      RECT 70.840 2.100 71.120 119.700 ;
      RECT 74.200 2.100 74.480 119.700 ;
      RECT 77.560 2.100 77.840 119.700 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 80.560 121.800 ;
    LAYER metal2 ;
    RECT 0 0 80.560 121.800 ;
    LAYER metal3 ;
    RECT 0.070 0 80.560 121.800 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.275 ;
    RECT 0 2.345 0.070 2.485 ;
    RECT 0 2.555 0.070 2.695 ;
    RECT 0 2.765 0.070 2.905 ;
    RECT 0 2.975 0.070 3.115 ;
    RECT 0 3.185 0.070 3.325 ;
    RECT 0 3.395 0.070 3.535 ;
    RECT 0 3.605 0.070 3.745 ;
    RECT 0 3.815 0.070 3.955 ;
    RECT 0 4.025 0.070 4.165 ;
    RECT 0 4.235 0.070 4.375 ;
    RECT 0 4.445 0.070 4.585 ;
    RECT 0 4.655 0.070 4.795 ;
    RECT 0 4.865 0.070 5.005 ;
    RECT 0 5.075 0.070 5.215 ;
    RECT 0 5.285 0.070 5.425 ;
    RECT 0 5.495 0.070 5.635 ;
    RECT 0 5.705 0.070 5.845 ;
    RECT 0 5.915 0.070 6.055 ;
    RECT 0 6.125 0.070 6.265 ;
    RECT 0 6.335 0.070 6.475 ;
    RECT 0 6.545 0.070 6.685 ;
    RECT 0 6.755 0.070 6.895 ;
    RECT 0 6.965 0.070 7.105 ;
    RECT 0 7.175 0.070 7.315 ;
    RECT 0 7.385 0.070 7.525 ;
    RECT 0 7.595 0.070 7.735 ;
    RECT 0 7.805 0.070 7.945 ;
    RECT 0 8.015 0.070 8.155 ;
    RECT 0 8.225 0.070 8.365 ;
    RECT 0 8.435 0.070 8.575 ;
    RECT 0 8.645 0.070 8.785 ;
    RECT 0 8.855 0.070 8.995 ;
    RECT 0 9.065 0.070 9.205 ;
    RECT 0 9.275 0.070 9.415 ;
    RECT 0 9.485 0.070 9.625 ;
    RECT 0 9.695 0.070 9.835 ;
    RECT 0 9.905 0.070 10.045 ;
    RECT 0 10.115 0.070 10.255 ;
    RECT 0 10.325 0.070 10.465 ;
    RECT 0 10.535 0.070 10.675 ;
    RECT 0 10.745 0.070 10.885 ;
    RECT 0 10.955 0.070 11.095 ;
    RECT 0 11.165 0.070 11.305 ;
    RECT 0 11.375 0.070 11.515 ;
    RECT 0 11.585 0.070 11.725 ;
    RECT 0 11.795 0.070 11.935 ;
    RECT 0 12.005 0.070 12.145 ;
    RECT 0 12.215 0.070 12.355 ;
    RECT 0 12.425 0.070 12.565 ;
    RECT 0 12.635 0.070 12.775 ;
    RECT 0 12.845 0.070 12.985 ;
    RECT 0 13.055 0.070 13.195 ;
    RECT 0 13.265 0.070 13.405 ;
    RECT 0 13.475 0.070 13.615 ;
    RECT 0 13.685 0.070 13.825 ;
    RECT 0 13.895 0.070 14.035 ;
    RECT 0 14.105 0.070 14.245 ;
    RECT 0 14.315 0.070 14.455 ;
    RECT 0 14.525 0.070 14.665 ;
    RECT 0 14.735 0.070 14.875 ;
    RECT 0 14.945 0.070 15.085 ;
    RECT 0 15.155 0.070 15.295 ;
    RECT 0 15.365 0.070 15.505 ;
    RECT 0 15.575 0.070 15.715 ;
    RECT 0 15.785 0.070 15.925 ;
    RECT 0 15.995 0.070 16.135 ;
    RECT 0 16.205 0.070 16.345 ;
    RECT 0 16.415 0.070 16.555 ;
    RECT 0 16.625 0.070 16.765 ;
    RECT 0 16.835 0.070 16.975 ;
    RECT 0 17.045 0.070 17.185 ;
    RECT 0 17.255 0.070 17.395 ;
    RECT 0 17.465 0.070 17.605 ;
    RECT 0 17.675 0.070 17.815 ;
    RECT 0 17.885 0.070 18.025 ;
    RECT 0 18.095 0.070 18.235 ;
    RECT 0 18.305 0.070 18.445 ;
    RECT 0 18.515 0.070 18.655 ;
    RECT 0 18.725 0.070 18.865 ;
    RECT 0 18.935 0.070 19.075 ;
    RECT 0 19.145 0.070 19.285 ;
    RECT 0 19.355 0.070 19.495 ;
    RECT 0 19.565 0.070 19.705 ;
    RECT 0 19.775 0.070 19.915 ;
    RECT 0 19.985 0.070 20.125 ;
    RECT 0 20.195 0.070 20.335 ;
    RECT 0 20.405 0.070 20.545 ;
    RECT 0 20.615 0.070 20.755 ;
    RECT 0 20.825 0.070 20.965 ;
    RECT 0 21.035 0.070 21.175 ;
    RECT 0 21.245 0.070 21.385 ;
    RECT 0 21.455 0.070 21.595 ;
    RECT 0 21.665 0.070 21.805 ;
    RECT 0 21.875 0.070 22.015 ;
    RECT 0 22.085 0.070 22.225 ;
    RECT 0 22.295 0.070 22.435 ;
    RECT 0 22.505 0.070 22.645 ;
    RECT 0 22.715 0.070 22.855 ;
    RECT 0 22.925 0.070 23.065 ;
    RECT 0 23.135 0.070 23.275 ;
    RECT 0 23.345 0.070 23.485 ;
    RECT 0 23.555 0.070 23.695 ;
    RECT 0 23.765 0.070 23.905 ;
    RECT 0 23.975 0.070 24.115 ;
    RECT 0 24.185 0.070 24.325 ;
    RECT 0 24.395 0.070 24.535 ;
    RECT 0 24.605 0.070 24.745 ;
    RECT 0 24.815 0.070 24.955 ;
    RECT 0 25.025 0.070 25.165 ;
    RECT 0 25.235 0.070 25.375 ;
    RECT 0 25.445 0.070 25.585 ;
    RECT 0 25.655 0.070 25.795 ;
    RECT 0 25.865 0.070 26.005 ;
    RECT 0 26.075 0.070 26.215 ;
    RECT 0 26.285 0.070 26.425 ;
    RECT 0 26.495 0.070 26.635 ;
    RECT 0 26.705 0.070 26.845 ;
    RECT 0 26.915 0.070 27.055 ;
    RECT 0 27.125 0.070 27.265 ;
    RECT 0 27.335 0.070 27.475 ;
    RECT 0 27.545 0.070 27.685 ;
    RECT 0 27.755 0.070 27.895 ;
    RECT 0 27.965 0.070 37.135 ;
    RECT 0 37.205 0.070 37.345 ;
    RECT 0 37.415 0.070 37.555 ;
    RECT 0 37.625 0.070 37.765 ;
    RECT 0 37.835 0.070 37.975 ;
    RECT 0 38.045 0.070 38.185 ;
    RECT 0 38.255 0.070 38.395 ;
    RECT 0 38.465 0.070 38.605 ;
    RECT 0 38.675 0.070 38.815 ;
    RECT 0 38.885 0.070 39.025 ;
    RECT 0 39.095 0.070 39.235 ;
    RECT 0 39.305 0.070 39.445 ;
    RECT 0 39.515 0.070 39.655 ;
    RECT 0 39.725 0.070 39.865 ;
    RECT 0 39.935 0.070 40.075 ;
    RECT 0 40.145 0.070 40.285 ;
    RECT 0 40.355 0.070 40.495 ;
    RECT 0 40.565 0.070 40.705 ;
    RECT 0 40.775 0.070 40.915 ;
    RECT 0 40.985 0.070 41.125 ;
    RECT 0 41.195 0.070 41.335 ;
    RECT 0 41.405 0.070 41.545 ;
    RECT 0 41.615 0.070 41.755 ;
    RECT 0 41.825 0.070 41.965 ;
    RECT 0 42.035 0.070 42.175 ;
    RECT 0 42.245 0.070 42.385 ;
    RECT 0 42.455 0.070 42.595 ;
    RECT 0 42.665 0.070 42.805 ;
    RECT 0 42.875 0.070 43.015 ;
    RECT 0 43.085 0.070 43.225 ;
    RECT 0 43.295 0.070 43.435 ;
    RECT 0 43.505 0.070 43.645 ;
    RECT 0 43.715 0.070 43.855 ;
    RECT 0 43.925 0.070 44.065 ;
    RECT 0 44.135 0.070 44.275 ;
    RECT 0 44.345 0.070 44.485 ;
    RECT 0 44.555 0.070 44.695 ;
    RECT 0 44.765 0.070 44.905 ;
    RECT 0 44.975 0.070 45.115 ;
    RECT 0 45.185 0.070 45.325 ;
    RECT 0 45.395 0.070 45.535 ;
    RECT 0 45.605 0.070 45.745 ;
    RECT 0 45.815 0.070 45.955 ;
    RECT 0 46.025 0.070 46.165 ;
    RECT 0 46.235 0.070 46.375 ;
    RECT 0 46.445 0.070 46.585 ;
    RECT 0 46.655 0.070 46.795 ;
    RECT 0 46.865 0.070 47.005 ;
    RECT 0 47.075 0.070 47.215 ;
    RECT 0 47.285 0.070 47.425 ;
    RECT 0 47.495 0.070 47.635 ;
    RECT 0 47.705 0.070 47.845 ;
    RECT 0 47.915 0.070 48.055 ;
    RECT 0 48.125 0.070 48.265 ;
    RECT 0 48.335 0.070 48.475 ;
    RECT 0 48.545 0.070 48.685 ;
    RECT 0 48.755 0.070 48.895 ;
    RECT 0 48.965 0.070 49.105 ;
    RECT 0 49.175 0.070 49.315 ;
    RECT 0 49.385 0.070 49.525 ;
    RECT 0 49.595 0.070 49.735 ;
    RECT 0 49.805 0.070 49.945 ;
    RECT 0 50.015 0.070 50.155 ;
    RECT 0 50.225 0.070 50.365 ;
    RECT 0 50.435 0.070 50.575 ;
    RECT 0 50.645 0.070 50.785 ;
    RECT 0 50.855 0.070 50.995 ;
    RECT 0 51.065 0.070 51.205 ;
    RECT 0 51.275 0.070 51.415 ;
    RECT 0 51.485 0.070 51.625 ;
    RECT 0 51.695 0.070 51.835 ;
    RECT 0 51.905 0.070 52.045 ;
    RECT 0 52.115 0.070 52.255 ;
    RECT 0 52.325 0.070 52.465 ;
    RECT 0 52.535 0.070 52.675 ;
    RECT 0 52.745 0.070 52.885 ;
    RECT 0 52.955 0.070 53.095 ;
    RECT 0 53.165 0.070 53.305 ;
    RECT 0 53.375 0.070 53.515 ;
    RECT 0 53.585 0.070 53.725 ;
    RECT 0 53.795 0.070 53.935 ;
    RECT 0 54.005 0.070 54.145 ;
    RECT 0 54.215 0.070 54.355 ;
    RECT 0 54.425 0.070 54.565 ;
    RECT 0 54.635 0.070 54.775 ;
    RECT 0 54.845 0.070 54.985 ;
    RECT 0 55.055 0.070 55.195 ;
    RECT 0 55.265 0.070 55.405 ;
    RECT 0 55.475 0.070 55.615 ;
    RECT 0 55.685 0.070 55.825 ;
    RECT 0 55.895 0.070 56.035 ;
    RECT 0 56.105 0.070 56.245 ;
    RECT 0 56.315 0.070 56.455 ;
    RECT 0 56.525 0.070 56.665 ;
    RECT 0 56.735 0.070 56.875 ;
    RECT 0 56.945 0.070 57.085 ;
    RECT 0 57.155 0.070 57.295 ;
    RECT 0 57.365 0.070 57.505 ;
    RECT 0 57.575 0.070 57.715 ;
    RECT 0 57.785 0.070 57.925 ;
    RECT 0 57.995 0.070 58.135 ;
    RECT 0 58.205 0.070 58.345 ;
    RECT 0 58.415 0.070 58.555 ;
    RECT 0 58.625 0.070 58.765 ;
    RECT 0 58.835 0.070 58.975 ;
    RECT 0 59.045 0.070 59.185 ;
    RECT 0 59.255 0.070 59.395 ;
    RECT 0 59.465 0.070 59.605 ;
    RECT 0 59.675 0.070 59.815 ;
    RECT 0 59.885 0.070 60.025 ;
    RECT 0 60.095 0.070 60.235 ;
    RECT 0 60.305 0.070 60.445 ;
    RECT 0 60.515 0.070 60.655 ;
    RECT 0 60.725 0.070 60.865 ;
    RECT 0 60.935 0.070 61.075 ;
    RECT 0 61.145 0.070 61.285 ;
    RECT 0 61.355 0.070 61.495 ;
    RECT 0 61.565 0.070 61.705 ;
    RECT 0 61.775 0.070 61.915 ;
    RECT 0 61.985 0.070 62.125 ;
    RECT 0 62.195 0.070 62.335 ;
    RECT 0 62.405 0.070 62.545 ;
    RECT 0 62.615 0.070 62.755 ;
    RECT 0 62.825 0.070 62.965 ;
    RECT 0 63.035 0.070 72.205 ;
    RECT 0 72.275 0.070 72.415 ;
    RECT 0 72.485 0.070 72.625 ;
    RECT 0 72.695 0.070 72.835 ;
    RECT 0 72.905 0.070 73.045 ;
    RECT 0 73.115 0.070 73.255 ;
    RECT 0 73.325 0.070 73.465 ;
    RECT 0 73.535 0.070 73.675 ;
    RECT 0 73.745 0.070 73.885 ;
    RECT 0 73.955 0.070 74.095 ;
    RECT 0 74.165 0.070 74.305 ;
    RECT 0 74.375 0.070 74.515 ;
    RECT 0 74.585 0.070 74.725 ;
    RECT 0 74.795 0.070 74.935 ;
    RECT 0 75.005 0.070 75.145 ;
    RECT 0 75.215 0.070 75.355 ;
    RECT 0 75.425 0.070 75.565 ;
    RECT 0 75.635 0.070 75.775 ;
    RECT 0 75.845 0.070 75.985 ;
    RECT 0 76.055 0.070 76.195 ;
    RECT 0 76.265 0.070 76.405 ;
    RECT 0 76.475 0.070 76.615 ;
    RECT 0 76.685 0.070 76.825 ;
    RECT 0 76.895 0.070 77.035 ;
    RECT 0 77.105 0.070 77.245 ;
    RECT 0 77.315 0.070 77.455 ;
    RECT 0 77.525 0.070 77.665 ;
    RECT 0 77.735 0.070 77.875 ;
    RECT 0 77.945 0.070 78.085 ;
    RECT 0 78.155 0.070 78.295 ;
    RECT 0 78.365 0.070 78.505 ;
    RECT 0 78.575 0.070 78.715 ;
    RECT 0 78.785 0.070 78.925 ;
    RECT 0 78.995 0.070 79.135 ;
    RECT 0 79.205 0.070 79.345 ;
    RECT 0 79.415 0.070 79.555 ;
    RECT 0 79.625 0.070 79.765 ;
    RECT 0 79.835 0.070 79.975 ;
    RECT 0 80.045 0.070 80.185 ;
    RECT 0 80.255 0.070 80.395 ;
    RECT 0 80.465 0.070 80.605 ;
    RECT 0 80.675 0.070 80.815 ;
    RECT 0 80.885 0.070 81.025 ;
    RECT 0 81.095 0.070 81.235 ;
    RECT 0 81.305 0.070 81.445 ;
    RECT 0 81.515 0.070 81.655 ;
    RECT 0 81.725 0.070 81.865 ;
    RECT 0 81.935 0.070 82.075 ;
    RECT 0 82.145 0.070 82.285 ;
    RECT 0 82.355 0.070 82.495 ;
    RECT 0 82.565 0.070 82.705 ;
    RECT 0 82.775 0.070 82.915 ;
    RECT 0 82.985 0.070 83.125 ;
    RECT 0 83.195 0.070 83.335 ;
    RECT 0 83.405 0.070 83.545 ;
    RECT 0 83.615 0.070 83.755 ;
    RECT 0 83.825 0.070 83.965 ;
    RECT 0 84.035 0.070 84.175 ;
    RECT 0 84.245 0.070 84.385 ;
    RECT 0 84.455 0.070 84.595 ;
    RECT 0 84.665 0.070 84.805 ;
    RECT 0 84.875 0.070 85.015 ;
    RECT 0 85.085 0.070 85.225 ;
    RECT 0 85.295 0.070 85.435 ;
    RECT 0 85.505 0.070 85.645 ;
    RECT 0 85.715 0.070 85.855 ;
    RECT 0 85.925 0.070 86.065 ;
    RECT 0 86.135 0.070 86.275 ;
    RECT 0 86.345 0.070 86.485 ;
    RECT 0 86.555 0.070 86.695 ;
    RECT 0 86.765 0.070 86.905 ;
    RECT 0 86.975 0.070 87.115 ;
    RECT 0 87.185 0.070 87.325 ;
    RECT 0 87.395 0.070 87.535 ;
    RECT 0 87.605 0.070 87.745 ;
    RECT 0 87.815 0.070 87.955 ;
    RECT 0 88.025 0.070 88.165 ;
    RECT 0 88.235 0.070 88.375 ;
    RECT 0 88.445 0.070 88.585 ;
    RECT 0 88.655 0.070 88.795 ;
    RECT 0 88.865 0.070 89.005 ;
    RECT 0 89.075 0.070 89.215 ;
    RECT 0 89.285 0.070 89.425 ;
    RECT 0 89.495 0.070 89.635 ;
    RECT 0 89.705 0.070 89.845 ;
    RECT 0 89.915 0.070 90.055 ;
    RECT 0 90.125 0.070 90.265 ;
    RECT 0 90.335 0.070 90.475 ;
    RECT 0 90.545 0.070 90.685 ;
    RECT 0 90.755 0.070 90.895 ;
    RECT 0 90.965 0.070 91.105 ;
    RECT 0 91.175 0.070 91.315 ;
    RECT 0 91.385 0.070 91.525 ;
    RECT 0 91.595 0.070 91.735 ;
    RECT 0 91.805 0.070 91.945 ;
    RECT 0 92.015 0.070 92.155 ;
    RECT 0 92.225 0.070 92.365 ;
    RECT 0 92.435 0.070 92.575 ;
    RECT 0 92.645 0.070 92.785 ;
    RECT 0 92.855 0.070 92.995 ;
    RECT 0 93.065 0.070 93.205 ;
    RECT 0 93.275 0.070 93.415 ;
    RECT 0 93.485 0.070 93.625 ;
    RECT 0 93.695 0.070 93.835 ;
    RECT 0 93.905 0.070 94.045 ;
    RECT 0 94.115 0.070 94.255 ;
    RECT 0 94.325 0.070 94.465 ;
    RECT 0 94.535 0.070 94.675 ;
    RECT 0 94.745 0.070 94.885 ;
    RECT 0 94.955 0.070 95.095 ;
    RECT 0 95.165 0.070 95.305 ;
    RECT 0 95.375 0.070 95.515 ;
    RECT 0 95.585 0.070 95.725 ;
    RECT 0 95.795 0.070 95.935 ;
    RECT 0 96.005 0.070 96.145 ;
    RECT 0 96.215 0.070 96.355 ;
    RECT 0 96.425 0.070 96.565 ;
    RECT 0 96.635 0.070 96.775 ;
    RECT 0 96.845 0.070 96.985 ;
    RECT 0 97.055 0.070 97.195 ;
    RECT 0 97.265 0.070 97.405 ;
    RECT 0 97.475 0.070 97.615 ;
    RECT 0 97.685 0.070 97.825 ;
    RECT 0 97.895 0.070 98.035 ;
    RECT 0 98.105 0.070 107.275 ;
    RECT 0 107.345 0.070 107.485 ;
    RECT 0 107.555 0.070 107.695 ;
    RECT 0 107.765 0.070 107.905 ;
    RECT 0 107.975 0.070 108.115 ;
    RECT 0 108.185 0.070 108.325 ;
    RECT 0 108.395 0.070 117.565 ;
    RECT 0 117.635 0.070 117.775 ;
    RECT 0 117.845 0.070 117.985 ;
    RECT 0 118.055 0.070 121.800 ;
    LAYER metal4 ;
    RECT 0 0 80.560 2.100 ;
    RECT 0 119.700 80.560 121.800 ;
    RECT 0.000 2.100 1.960 119.700 ;
    RECT 2.240 2.100 3.640 119.700 ;
    RECT 3.920 2.100 5.320 119.700 ;
    RECT 5.600 2.100 7.000 119.700 ;
    RECT 7.280 2.100 8.680 119.700 ;
    RECT 8.960 2.100 10.360 119.700 ;
    RECT 10.640 2.100 12.040 119.700 ;
    RECT 12.320 2.100 13.720 119.700 ;
    RECT 14.000 2.100 15.400 119.700 ;
    RECT 15.680 2.100 17.080 119.700 ;
    RECT 17.360 2.100 18.760 119.700 ;
    RECT 19.040 2.100 20.440 119.700 ;
    RECT 20.720 2.100 22.120 119.700 ;
    RECT 22.400 2.100 23.800 119.700 ;
    RECT 24.080 2.100 25.480 119.700 ;
    RECT 25.760 2.100 27.160 119.700 ;
    RECT 27.440 2.100 28.840 119.700 ;
    RECT 29.120 2.100 30.520 119.700 ;
    RECT 30.800 2.100 32.200 119.700 ;
    RECT 32.480 2.100 33.880 119.700 ;
    RECT 34.160 2.100 35.560 119.700 ;
    RECT 35.840 2.100 37.240 119.700 ;
    RECT 37.520 2.100 38.920 119.700 ;
    RECT 39.200 2.100 40.600 119.700 ;
    RECT 40.880 2.100 42.280 119.700 ;
    RECT 42.560 2.100 43.960 119.700 ;
    RECT 44.240 2.100 45.640 119.700 ;
    RECT 45.920 2.100 47.320 119.700 ;
    RECT 47.600 2.100 49.000 119.700 ;
    RECT 49.280 2.100 50.680 119.700 ;
    RECT 50.960 2.100 52.360 119.700 ;
    RECT 52.640 2.100 54.040 119.700 ;
    RECT 54.320 2.100 55.720 119.700 ;
    RECT 56.000 2.100 57.400 119.700 ;
    RECT 57.680 2.100 59.080 119.700 ;
    RECT 59.360 2.100 60.760 119.700 ;
    RECT 61.040 2.100 62.440 119.700 ;
    RECT 62.720 2.100 64.120 119.700 ;
    RECT 64.400 2.100 65.800 119.700 ;
    RECT 66.080 2.100 67.480 119.700 ;
    RECT 67.760 2.100 69.160 119.700 ;
    RECT 69.440 2.100 70.840 119.700 ;
    RECT 71.120 2.100 72.520 119.700 ;
    RECT 72.800 2.100 74.200 119.700 ;
    RECT 74.480 2.100 75.880 119.700 ;
    RECT 76.160 2.100 77.560 119.700 ;
    RECT 77.840 2.100 80.560 119.700 ;
    LAYER OVERLAP ;
    RECT 0 0 80.560 121.800 ;
  END
END fakeram45_64x124

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_64x96
  FOREIGN fakeram45_64x96 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 54.530 BY 77.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.275 0.070 2.345 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.695 0.070 2.765 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.115 0.070 3.185 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.535 0.070 3.605 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.955 0.070 4.025 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.375 0.070 4.445 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.795 0.070 4.865 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.215 0.070 5.285 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.635 0.070 5.705 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.055 0.070 6.125 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.475 0.070 6.545 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.895 0.070 6.965 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.315 0.070 7.385 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.735 0.070 7.805 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.155 0.070 8.225 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.575 0.070 8.645 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.785 0.070 8.855 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.995 0.070 9.065 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.415 0.070 9.485 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.835 0.070 9.905 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.255 0.070 10.325 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.675 0.070 10.745 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.095 0.070 11.165 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.515 0.070 11.585 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.935 0.070 12.005 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.355 0.070 12.425 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.775 0.070 12.845 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.985 0.070 13.055 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.195 0.070 13.265 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.615 0.070 13.685 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.035 0.070 14.105 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.455 0.070 14.525 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.875 0.070 14.945 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.295 0.070 15.365 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.505 0.070 15.575 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.715 0.070 15.785 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.135 0.070 16.205 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.345 0.070 16.415 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.555 0.070 16.625 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.975 0.070 17.045 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.185 0.070 17.255 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.395 0.070 17.465 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.605 0.070 17.675 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.815 0.070 17.885 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.025 0.070 18.095 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.235 0.070 18.305 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.655 0.070 18.725 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.075 0.070 19.145 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.495 0.070 19.565 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.915 0.070 19.985 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.335 0.070 20.405 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.545 0.070 20.615 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.755 0.070 20.825 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.175 0.070 21.245 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.595 0.070 21.665 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END w_mask_in[94]
  PIN w_mask_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.015 0.070 22.085 ;
    END
  END w_mask_in[95]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.535 0.070 24.605 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.955 0.070 25.025 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.375 0.070 25.445 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.795 0.070 25.865 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.215 0.070 26.285 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.425 0.070 26.495 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.635 0.070 26.705 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.055 0.070 27.125 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.475 0.070 27.545 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.685 0.070 27.755 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.895 0.070 27.965 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.105 0.070 28.175 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.315 0.070 28.385 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.735 0.070 28.805 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.945 0.070 29.015 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.155 0.070 29.225 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.575 0.070 29.645 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.785 0.070 29.855 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.995 0.070 30.065 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.205 0.070 30.275 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.415 0.070 30.485 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.625 0.070 30.695 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.835 0.070 30.905 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.045 0.070 31.115 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.255 0.070 31.325 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.465 0.070 31.535 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.675 0.070 31.745 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.885 0.070 31.955 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.095 0.070 32.165 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.305 0.070 32.375 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.515 0.070 32.585 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.935 0.070 33.005 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.145 0.070 33.215 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.355 0.070 33.425 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.775 0.070 33.845 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.985 0.070 34.055 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.195 0.070 34.265 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.615 0.070 34.685 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.825 0.070 34.895 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.035 0.070 35.105 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.455 0.070 35.525 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.875 0.070 35.945 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.295 0.070 36.365 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.505 0.070 36.575 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.715 0.070 36.785 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.135 0.070 37.205 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.555 0.070 37.625 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.975 0.070 38.045 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.185 0.070 38.255 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.395 0.070 38.465 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.815 0.070 38.885 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.235 0.070 39.305 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.655 0.070 39.725 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.075 0.070 40.145 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.495 0.070 40.565 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.915 0.070 40.985 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.335 0.070 41.405 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.755 0.070 41.825 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.175 0.070 42.245 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.595 0.070 42.665 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.015 0.070 43.085 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.435 0.070 43.505 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.855 0.070 43.925 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.275 0.070 44.345 ;
    END
  END rd_out[94]
  PIN rd_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END rd_out[95]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.215 0.070 47.285 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.635 0.070 47.705 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.055 0.070 48.125 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.265 0.070 48.335 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.475 0.070 48.545 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.895 0.070 48.965 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.315 0.070 49.385 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.735 0.070 49.805 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.945 0.070 50.015 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.155 0.070 50.225 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.575 0.070 50.645 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.785 0.070 50.855 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.995 0.070 51.065 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.205 0.070 51.275 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.415 0.070 51.485 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.625 0.070 51.695 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.835 0.070 51.905 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.045 0.070 52.115 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.255 0.070 52.325 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.675 0.070 52.745 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.095 0.070 53.165 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.305 0.070 53.375 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.515 0.070 53.585 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.935 0.070 54.005 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.145 0.070 54.215 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.355 0.070 54.425 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.775 0.070 54.845 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.985 0.070 55.055 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.195 0.070 55.265 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.615 0.070 55.685 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.825 0.070 55.895 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.035 0.070 56.105 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.455 0.070 56.525 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.665 0.070 56.735 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.875 0.070 56.945 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.085 0.070 57.155 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.295 0.070 57.365 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.505 0.070 57.575 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.715 0.070 57.785 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.135 0.070 58.205 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.345 0.070 58.415 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.555 0.070 58.625 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.765 0.070 58.835 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.975 0.070 59.045 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.185 0.070 59.255 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.395 0.070 59.465 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.605 0.070 59.675 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.815 0.070 59.885 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.025 0.070 60.095 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.235 0.070 60.305 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.445 0.070 60.515 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.655 0.070 60.725 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.865 0.070 60.935 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.075 0.070 61.145 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.285 0.070 61.355 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.495 0.070 61.565 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.705 0.070 61.775 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.915 0.070 61.985 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.125 0.070 62.195 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.335 0.070 62.405 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.545 0.070 62.615 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.755 0.070 62.825 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.965 0.070 63.035 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.175 0.070 63.245 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.385 0.070 63.455 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.595 0.070 63.665 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.805 0.070 63.875 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.015 0.070 64.085 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.225 0.070 64.295 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.435 0.070 64.505 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.645 0.070 64.715 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.855 0.070 64.925 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.065 0.070 65.135 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.275 0.070 65.345 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.485 0.070 65.555 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.695 0.070 65.765 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.905 0.070 65.975 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.115 0.070 66.185 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.325 0.070 66.395 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.535 0.070 66.605 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.745 0.070 66.815 ;
    END
  END wd_in[94]
  PIN wd_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.955 0.070 67.025 ;
    END
  END wd_in[95]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.475 0.070 69.545 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.685 0.070 69.755 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.895 0.070 69.965 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.105 0.070 70.175 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.315 0.070 70.385 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.255 0.070 73.325 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.465 0.070 73.535 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 74.900 ;
      RECT 5.320 2.100 5.600 74.900 ;
      RECT 8.680 2.100 8.960 74.900 ;
      RECT 12.040 2.100 12.320 74.900 ;
      RECT 15.400 2.100 15.680 74.900 ;
      RECT 18.760 2.100 19.040 74.900 ;
      RECT 22.120 2.100 22.400 74.900 ;
      RECT 25.480 2.100 25.760 74.900 ;
      RECT 28.840 2.100 29.120 74.900 ;
      RECT 32.200 2.100 32.480 74.900 ;
      RECT 35.560 2.100 35.840 74.900 ;
      RECT 38.920 2.100 39.200 74.900 ;
      RECT 42.280 2.100 42.560 74.900 ;
      RECT 45.640 2.100 45.920 74.900 ;
      RECT 49.000 2.100 49.280 74.900 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 74.900 ;
      RECT 7.000 2.100 7.280 74.900 ;
      RECT 10.360 2.100 10.640 74.900 ;
      RECT 13.720 2.100 14.000 74.900 ;
      RECT 17.080 2.100 17.360 74.900 ;
      RECT 20.440 2.100 20.720 74.900 ;
      RECT 23.800 2.100 24.080 74.900 ;
      RECT 27.160 2.100 27.440 74.900 ;
      RECT 30.520 2.100 30.800 74.900 ;
      RECT 33.880 2.100 34.160 74.900 ;
      RECT 37.240 2.100 37.520 74.900 ;
      RECT 40.600 2.100 40.880 74.900 ;
      RECT 43.960 2.100 44.240 74.900 ;
      RECT 47.320 2.100 47.600 74.900 ;
      RECT 50.680 2.100 50.960 74.900 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 54.530 77.000 ;
    LAYER metal2 ;
    RECT 0 0 54.530 77.000 ;
    LAYER metal3 ;
    RECT 0.070 0 54.530 77.000 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.275 ;
    RECT 0 2.345 0.070 2.485 ;
    RECT 0 2.555 0.070 2.695 ;
    RECT 0 2.765 0.070 2.905 ;
    RECT 0 2.975 0.070 3.115 ;
    RECT 0 3.185 0.070 3.325 ;
    RECT 0 3.395 0.070 3.535 ;
    RECT 0 3.605 0.070 3.745 ;
    RECT 0 3.815 0.070 3.955 ;
    RECT 0 4.025 0.070 4.165 ;
    RECT 0 4.235 0.070 4.375 ;
    RECT 0 4.445 0.070 4.585 ;
    RECT 0 4.655 0.070 4.795 ;
    RECT 0 4.865 0.070 5.005 ;
    RECT 0 5.075 0.070 5.215 ;
    RECT 0 5.285 0.070 5.425 ;
    RECT 0 5.495 0.070 5.635 ;
    RECT 0 5.705 0.070 5.845 ;
    RECT 0 5.915 0.070 6.055 ;
    RECT 0 6.125 0.070 6.265 ;
    RECT 0 6.335 0.070 6.475 ;
    RECT 0 6.545 0.070 6.685 ;
    RECT 0 6.755 0.070 6.895 ;
    RECT 0 6.965 0.070 7.105 ;
    RECT 0 7.175 0.070 7.315 ;
    RECT 0 7.385 0.070 7.525 ;
    RECT 0 7.595 0.070 7.735 ;
    RECT 0 7.805 0.070 7.945 ;
    RECT 0 8.015 0.070 8.155 ;
    RECT 0 8.225 0.070 8.365 ;
    RECT 0 8.435 0.070 8.575 ;
    RECT 0 8.645 0.070 8.785 ;
    RECT 0 8.855 0.070 8.995 ;
    RECT 0 9.065 0.070 9.205 ;
    RECT 0 9.275 0.070 9.415 ;
    RECT 0 9.485 0.070 9.625 ;
    RECT 0 9.695 0.070 9.835 ;
    RECT 0 9.905 0.070 10.045 ;
    RECT 0 10.115 0.070 10.255 ;
    RECT 0 10.325 0.070 10.465 ;
    RECT 0 10.535 0.070 10.675 ;
    RECT 0 10.745 0.070 10.885 ;
    RECT 0 10.955 0.070 11.095 ;
    RECT 0 11.165 0.070 11.305 ;
    RECT 0 11.375 0.070 11.515 ;
    RECT 0 11.585 0.070 11.725 ;
    RECT 0 11.795 0.070 11.935 ;
    RECT 0 12.005 0.070 12.145 ;
    RECT 0 12.215 0.070 12.355 ;
    RECT 0 12.425 0.070 12.565 ;
    RECT 0 12.635 0.070 12.775 ;
    RECT 0 12.845 0.070 12.985 ;
    RECT 0 13.055 0.070 13.195 ;
    RECT 0 13.265 0.070 13.405 ;
    RECT 0 13.475 0.070 13.615 ;
    RECT 0 13.685 0.070 13.825 ;
    RECT 0 13.895 0.070 14.035 ;
    RECT 0 14.105 0.070 14.245 ;
    RECT 0 14.315 0.070 14.455 ;
    RECT 0 14.525 0.070 14.665 ;
    RECT 0 14.735 0.070 14.875 ;
    RECT 0 14.945 0.070 15.085 ;
    RECT 0 15.155 0.070 15.295 ;
    RECT 0 15.365 0.070 15.505 ;
    RECT 0 15.575 0.070 15.715 ;
    RECT 0 15.785 0.070 15.925 ;
    RECT 0 15.995 0.070 16.135 ;
    RECT 0 16.205 0.070 16.345 ;
    RECT 0 16.415 0.070 16.555 ;
    RECT 0 16.625 0.070 16.765 ;
    RECT 0 16.835 0.070 16.975 ;
    RECT 0 17.045 0.070 17.185 ;
    RECT 0 17.255 0.070 17.395 ;
    RECT 0 17.465 0.070 17.605 ;
    RECT 0 17.675 0.070 17.815 ;
    RECT 0 17.885 0.070 18.025 ;
    RECT 0 18.095 0.070 18.235 ;
    RECT 0 18.305 0.070 18.445 ;
    RECT 0 18.515 0.070 18.655 ;
    RECT 0 18.725 0.070 18.865 ;
    RECT 0 18.935 0.070 19.075 ;
    RECT 0 19.145 0.070 19.285 ;
    RECT 0 19.355 0.070 19.495 ;
    RECT 0 19.565 0.070 19.705 ;
    RECT 0 19.775 0.070 19.915 ;
    RECT 0 19.985 0.070 20.125 ;
    RECT 0 20.195 0.070 20.335 ;
    RECT 0 20.405 0.070 20.545 ;
    RECT 0 20.615 0.070 20.755 ;
    RECT 0 20.825 0.070 20.965 ;
    RECT 0 21.035 0.070 21.175 ;
    RECT 0 21.245 0.070 21.385 ;
    RECT 0 21.455 0.070 21.595 ;
    RECT 0 21.665 0.070 21.805 ;
    RECT 0 21.875 0.070 22.015 ;
    RECT 0 22.085 0.070 24.535 ;
    RECT 0 24.605 0.070 24.745 ;
    RECT 0 24.815 0.070 24.955 ;
    RECT 0 25.025 0.070 25.165 ;
    RECT 0 25.235 0.070 25.375 ;
    RECT 0 25.445 0.070 25.585 ;
    RECT 0 25.655 0.070 25.795 ;
    RECT 0 25.865 0.070 26.005 ;
    RECT 0 26.075 0.070 26.215 ;
    RECT 0 26.285 0.070 26.425 ;
    RECT 0 26.495 0.070 26.635 ;
    RECT 0 26.705 0.070 26.845 ;
    RECT 0 26.915 0.070 27.055 ;
    RECT 0 27.125 0.070 27.265 ;
    RECT 0 27.335 0.070 27.475 ;
    RECT 0 27.545 0.070 27.685 ;
    RECT 0 27.755 0.070 27.895 ;
    RECT 0 27.965 0.070 28.105 ;
    RECT 0 28.175 0.070 28.315 ;
    RECT 0 28.385 0.070 28.525 ;
    RECT 0 28.595 0.070 28.735 ;
    RECT 0 28.805 0.070 28.945 ;
    RECT 0 29.015 0.070 29.155 ;
    RECT 0 29.225 0.070 29.365 ;
    RECT 0 29.435 0.070 29.575 ;
    RECT 0 29.645 0.070 29.785 ;
    RECT 0 29.855 0.070 29.995 ;
    RECT 0 30.065 0.070 30.205 ;
    RECT 0 30.275 0.070 30.415 ;
    RECT 0 30.485 0.070 30.625 ;
    RECT 0 30.695 0.070 30.835 ;
    RECT 0 30.905 0.070 31.045 ;
    RECT 0 31.115 0.070 31.255 ;
    RECT 0 31.325 0.070 31.465 ;
    RECT 0 31.535 0.070 31.675 ;
    RECT 0 31.745 0.070 31.885 ;
    RECT 0 31.955 0.070 32.095 ;
    RECT 0 32.165 0.070 32.305 ;
    RECT 0 32.375 0.070 32.515 ;
    RECT 0 32.585 0.070 32.725 ;
    RECT 0 32.795 0.070 32.935 ;
    RECT 0 33.005 0.070 33.145 ;
    RECT 0 33.215 0.070 33.355 ;
    RECT 0 33.425 0.070 33.565 ;
    RECT 0 33.635 0.070 33.775 ;
    RECT 0 33.845 0.070 33.985 ;
    RECT 0 34.055 0.070 34.195 ;
    RECT 0 34.265 0.070 34.405 ;
    RECT 0 34.475 0.070 34.615 ;
    RECT 0 34.685 0.070 34.825 ;
    RECT 0 34.895 0.070 35.035 ;
    RECT 0 35.105 0.070 35.245 ;
    RECT 0 35.315 0.070 35.455 ;
    RECT 0 35.525 0.070 35.665 ;
    RECT 0 35.735 0.070 35.875 ;
    RECT 0 35.945 0.070 36.085 ;
    RECT 0 36.155 0.070 36.295 ;
    RECT 0 36.365 0.070 36.505 ;
    RECT 0 36.575 0.070 36.715 ;
    RECT 0 36.785 0.070 36.925 ;
    RECT 0 36.995 0.070 37.135 ;
    RECT 0 37.205 0.070 37.345 ;
    RECT 0 37.415 0.070 37.555 ;
    RECT 0 37.625 0.070 37.765 ;
    RECT 0 37.835 0.070 37.975 ;
    RECT 0 38.045 0.070 38.185 ;
    RECT 0 38.255 0.070 38.395 ;
    RECT 0 38.465 0.070 38.605 ;
    RECT 0 38.675 0.070 38.815 ;
    RECT 0 38.885 0.070 39.025 ;
    RECT 0 39.095 0.070 39.235 ;
    RECT 0 39.305 0.070 39.445 ;
    RECT 0 39.515 0.070 39.655 ;
    RECT 0 39.725 0.070 39.865 ;
    RECT 0 39.935 0.070 40.075 ;
    RECT 0 40.145 0.070 40.285 ;
    RECT 0 40.355 0.070 40.495 ;
    RECT 0 40.565 0.070 40.705 ;
    RECT 0 40.775 0.070 40.915 ;
    RECT 0 40.985 0.070 41.125 ;
    RECT 0 41.195 0.070 41.335 ;
    RECT 0 41.405 0.070 41.545 ;
    RECT 0 41.615 0.070 41.755 ;
    RECT 0 41.825 0.070 41.965 ;
    RECT 0 42.035 0.070 42.175 ;
    RECT 0 42.245 0.070 42.385 ;
    RECT 0 42.455 0.070 42.595 ;
    RECT 0 42.665 0.070 42.805 ;
    RECT 0 42.875 0.070 43.015 ;
    RECT 0 43.085 0.070 43.225 ;
    RECT 0 43.295 0.070 43.435 ;
    RECT 0 43.505 0.070 43.645 ;
    RECT 0 43.715 0.070 43.855 ;
    RECT 0 43.925 0.070 44.065 ;
    RECT 0 44.135 0.070 44.275 ;
    RECT 0 44.345 0.070 44.485 ;
    RECT 0 44.555 0.070 47.005 ;
    RECT 0 47.075 0.070 47.215 ;
    RECT 0 47.285 0.070 47.425 ;
    RECT 0 47.495 0.070 47.635 ;
    RECT 0 47.705 0.070 47.845 ;
    RECT 0 47.915 0.070 48.055 ;
    RECT 0 48.125 0.070 48.265 ;
    RECT 0 48.335 0.070 48.475 ;
    RECT 0 48.545 0.070 48.685 ;
    RECT 0 48.755 0.070 48.895 ;
    RECT 0 48.965 0.070 49.105 ;
    RECT 0 49.175 0.070 49.315 ;
    RECT 0 49.385 0.070 49.525 ;
    RECT 0 49.595 0.070 49.735 ;
    RECT 0 49.805 0.070 49.945 ;
    RECT 0 50.015 0.070 50.155 ;
    RECT 0 50.225 0.070 50.365 ;
    RECT 0 50.435 0.070 50.575 ;
    RECT 0 50.645 0.070 50.785 ;
    RECT 0 50.855 0.070 50.995 ;
    RECT 0 51.065 0.070 51.205 ;
    RECT 0 51.275 0.070 51.415 ;
    RECT 0 51.485 0.070 51.625 ;
    RECT 0 51.695 0.070 51.835 ;
    RECT 0 51.905 0.070 52.045 ;
    RECT 0 52.115 0.070 52.255 ;
    RECT 0 52.325 0.070 52.465 ;
    RECT 0 52.535 0.070 52.675 ;
    RECT 0 52.745 0.070 52.885 ;
    RECT 0 52.955 0.070 53.095 ;
    RECT 0 53.165 0.070 53.305 ;
    RECT 0 53.375 0.070 53.515 ;
    RECT 0 53.585 0.070 53.725 ;
    RECT 0 53.795 0.070 53.935 ;
    RECT 0 54.005 0.070 54.145 ;
    RECT 0 54.215 0.070 54.355 ;
    RECT 0 54.425 0.070 54.565 ;
    RECT 0 54.635 0.070 54.775 ;
    RECT 0 54.845 0.070 54.985 ;
    RECT 0 55.055 0.070 55.195 ;
    RECT 0 55.265 0.070 55.405 ;
    RECT 0 55.475 0.070 55.615 ;
    RECT 0 55.685 0.070 55.825 ;
    RECT 0 55.895 0.070 56.035 ;
    RECT 0 56.105 0.070 56.245 ;
    RECT 0 56.315 0.070 56.455 ;
    RECT 0 56.525 0.070 56.665 ;
    RECT 0 56.735 0.070 56.875 ;
    RECT 0 56.945 0.070 57.085 ;
    RECT 0 57.155 0.070 57.295 ;
    RECT 0 57.365 0.070 57.505 ;
    RECT 0 57.575 0.070 57.715 ;
    RECT 0 57.785 0.070 57.925 ;
    RECT 0 57.995 0.070 58.135 ;
    RECT 0 58.205 0.070 58.345 ;
    RECT 0 58.415 0.070 58.555 ;
    RECT 0 58.625 0.070 58.765 ;
    RECT 0 58.835 0.070 58.975 ;
    RECT 0 59.045 0.070 59.185 ;
    RECT 0 59.255 0.070 59.395 ;
    RECT 0 59.465 0.070 59.605 ;
    RECT 0 59.675 0.070 59.815 ;
    RECT 0 59.885 0.070 60.025 ;
    RECT 0 60.095 0.070 60.235 ;
    RECT 0 60.305 0.070 60.445 ;
    RECT 0 60.515 0.070 60.655 ;
    RECT 0 60.725 0.070 60.865 ;
    RECT 0 60.935 0.070 61.075 ;
    RECT 0 61.145 0.070 61.285 ;
    RECT 0 61.355 0.070 61.495 ;
    RECT 0 61.565 0.070 61.705 ;
    RECT 0 61.775 0.070 61.915 ;
    RECT 0 61.985 0.070 62.125 ;
    RECT 0 62.195 0.070 62.335 ;
    RECT 0 62.405 0.070 62.545 ;
    RECT 0 62.615 0.070 62.755 ;
    RECT 0 62.825 0.070 62.965 ;
    RECT 0 63.035 0.070 63.175 ;
    RECT 0 63.245 0.070 63.385 ;
    RECT 0 63.455 0.070 63.595 ;
    RECT 0 63.665 0.070 63.805 ;
    RECT 0 63.875 0.070 64.015 ;
    RECT 0 64.085 0.070 64.225 ;
    RECT 0 64.295 0.070 64.435 ;
    RECT 0 64.505 0.070 64.645 ;
    RECT 0 64.715 0.070 64.855 ;
    RECT 0 64.925 0.070 65.065 ;
    RECT 0 65.135 0.070 65.275 ;
    RECT 0 65.345 0.070 65.485 ;
    RECT 0 65.555 0.070 65.695 ;
    RECT 0 65.765 0.070 65.905 ;
    RECT 0 65.975 0.070 66.115 ;
    RECT 0 66.185 0.070 66.325 ;
    RECT 0 66.395 0.070 66.535 ;
    RECT 0 66.605 0.070 66.745 ;
    RECT 0 66.815 0.070 66.955 ;
    RECT 0 67.025 0.070 69.475 ;
    RECT 0 69.545 0.070 69.685 ;
    RECT 0 69.755 0.070 69.895 ;
    RECT 0 69.965 0.070 70.105 ;
    RECT 0 70.175 0.070 70.315 ;
    RECT 0 70.385 0.070 70.525 ;
    RECT 0 70.595 0.070 73.045 ;
    RECT 0 73.115 0.070 73.255 ;
    RECT 0 73.325 0.070 73.465 ;
    RECT 0 73.535 0.070 77.000 ;
    LAYER metal4 ;
    RECT 0 0 54.530 2.100 ;
    RECT 0 74.900 54.530 77.000 ;
    RECT 0.000 2.100 1.960 74.900 ;
    RECT 2.240 2.100 3.640 74.900 ;
    RECT 3.920 2.100 5.320 74.900 ;
    RECT 5.600 2.100 7.000 74.900 ;
    RECT 7.280 2.100 8.680 74.900 ;
    RECT 8.960 2.100 10.360 74.900 ;
    RECT 10.640 2.100 12.040 74.900 ;
    RECT 12.320 2.100 13.720 74.900 ;
    RECT 14.000 2.100 15.400 74.900 ;
    RECT 15.680 2.100 17.080 74.900 ;
    RECT 17.360 2.100 18.760 74.900 ;
    RECT 19.040 2.100 20.440 74.900 ;
    RECT 20.720 2.100 22.120 74.900 ;
    RECT 22.400 2.100 23.800 74.900 ;
    RECT 24.080 2.100 25.480 74.900 ;
    RECT 25.760 2.100 27.160 74.900 ;
    RECT 27.440 2.100 28.840 74.900 ;
    RECT 29.120 2.100 30.520 74.900 ;
    RECT 30.800 2.100 32.200 74.900 ;
    RECT 32.480 2.100 33.880 74.900 ;
    RECT 34.160 2.100 35.560 74.900 ;
    RECT 35.840 2.100 37.240 74.900 ;
    RECT 37.520 2.100 38.920 74.900 ;
    RECT 39.200 2.100 40.600 74.900 ;
    RECT 40.880 2.100 42.280 74.900 ;
    RECT 42.560 2.100 43.960 74.900 ;
    RECT 44.240 2.100 45.640 74.900 ;
    RECT 45.920 2.100 47.320 74.900 ;
    RECT 47.600 2.100 49.000 74.900 ;
    RECT 49.280 2.100 50.680 74.900 ;
    RECT 50.960 2.100 54.530 74.900 ;
    LAYER OVERLAP ;
    RECT 0 0 54.530 77.000 ;
  END
END fakeram45_64x96

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_64x64
  FOREIGN fakeram45_64x64 0 0 ;
  SYMMETRY X Y ;
  SIZE 56.050 BY 102.200 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.785 0.070 8.855 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.985 0.070 13.055 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.505 0.070 15.575 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.345 0.070 16.415 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.185 0.070 17.255 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.605 0.070 17.675 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.025 0.070 18.095 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.545 0.070 20.615 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.225 0.070 22.295 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.905 0.070 23.975 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.425 0.070 26.495 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.685 0.070 27.755 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.105 0.070 28.175 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END w_mask_in[63]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.885 0.070 31.955 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.305 0.070 32.375 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.145 0.070 33.215 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.985 0.070 34.055 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.825 0.070 34.895 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.505 0.070 36.575 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.185 0.070 38.255 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.325 0.070 45.395 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.745 0.070 45.815 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.585 0.070 46.655 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.265 0.070 48.335 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.945 0.070 50.015 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.785 0.070 50.855 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.205 0.070 51.275 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.625 0.070 51.695 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.045 0.070 52.115 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.305 0.070 53.375 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.145 0.070 54.215 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.985 0.070 55.055 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.825 0.070 55.895 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.665 0.070 56.735 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.085 0.070 57.155 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.505 0.070 57.575 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.345 0.070 58.415 ;
    END
  END rd_out[63]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.705 0.070 61.775 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.125 0.070 62.195 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.545 0.070 62.615 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.965 0.070 63.035 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.385 0.070 63.455 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.805 0.070 63.875 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.225 0.070 64.295 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.645 0.070 64.715 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.065 0.070 65.135 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.485 0.070 65.555 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.905 0.070 65.975 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.325 0.070 66.395 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.745 0.070 66.815 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.165 0.070 67.235 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.585 0.070 67.655 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.425 0.070 68.495 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.845 0.070 68.915 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.265 0.070 69.335 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.685 0.070 69.755 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.105 0.070 70.175 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.945 0.070 71.015 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.785 0.070 71.855 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.205 0.070 72.275 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.625 0.070 72.695 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.465 0.070 73.535 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.305 0.070 74.375 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.725 0.070 74.795 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.145 0.070 75.215 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.405 0.070 76.475 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.825 0.070 76.895 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.245 0.070 77.315 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.665 0.070 77.735 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.085 0.070 78.155 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.505 0.070 78.575 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.925 0.070 78.995 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.345 0.070 79.415 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.185 0.070 80.255 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.605 0.070 80.675 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.025 0.070 81.095 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.445 0.070 81.515 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.285 0.070 82.355 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.705 0.070 82.775 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.125 0.070 83.195 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.545 0.070 83.615 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.965 0.070 84.035 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.385 0.070 84.455 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.225 0.070 85.295 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.065 0.070 86.135 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.485 0.070 86.555 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.905 0.070 86.975 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.325 0.070 87.395 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.745 0.070 87.815 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.165 0.070 88.235 ;
    END
  END wd_in[63]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.525 0.070 91.595 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.945 0.070 92.015 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.365 0.070 92.435 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.785 0.070 92.855 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.205 0.070 93.275 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.625 0.070 93.695 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.985 0.070 97.055 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.405 0.070 97.475 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.825 0.070 97.895 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 100.100 ;
      RECT 5.320 2.100 5.600 100.100 ;
      RECT 8.680 2.100 8.960 100.100 ;
      RECT 12.040 2.100 12.320 100.100 ;
      RECT 15.400 2.100 15.680 100.100 ;
      RECT 18.760 2.100 19.040 100.100 ;
      RECT 22.120 2.100 22.400 100.100 ;
      RECT 25.480 2.100 25.760 100.100 ;
      RECT 28.840 2.100 29.120 100.100 ;
      RECT 32.200 2.100 32.480 100.100 ;
      RECT 35.560 2.100 35.840 100.100 ;
      RECT 38.920 2.100 39.200 100.100 ;
      RECT 42.280 2.100 42.560 100.100 ;
      RECT 45.640 2.100 45.920 100.100 ;
      RECT 49.000 2.100 49.280 100.100 ;
      RECT 52.360 2.100 52.640 100.100 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 100.100 ;
      RECT 7.000 2.100 7.280 100.100 ;
      RECT 10.360 2.100 10.640 100.100 ;
      RECT 13.720 2.100 14.000 100.100 ;
      RECT 17.080 2.100 17.360 100.100 ;
      RECT 20.440 2.100 20.720 100.100 ;
      RECT 23.800 2.100 24.080 100.100 ;
      RECT 27.160 2.100 27.440 100.100 ;
      RECT 30.520 2.100 30.800 100.100 ;
      RECT 33.880 2.100 34.160 100.100 ;
      RECT 37.240 2.100 37.520 100.100 ;
      RECT 40.600 2.100 40.880 100.100 ;
      RECT 43.960 2.100 44.240 100.100 ;
      RECT 47.320 2.100 47.600 100.100 ;
      RECT 50.680 2.100 50.960 100.100 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 56.050 102.200 ;
    LAYER metal2 ;
    RECT 0 0 56.050 102.200 ;
    LAYER metal3 ;
    RECT 0.070 0 56.050 102.200 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.485 ;
    RECT 0 2.555 0.070 2.905 ;
    RECT 0 2.975 0.070 3.325 ;
    RECT 0 3.395 0.070 3.745 ;
    RECT 0 3.815 0.070 4.165 ;
    RECT 0 4.235 0.070 4.585 ;
    RECT 0 4.655 0.070 5.005 ;
    RECT 0 5.075 0.070 5.425 ;
    RECT 0 5.495 0.070 5.845 ;
    RECT 0 5.915 0.070 6.265 ;
    RECT 0 6.335 0.070 6.685 ;
    RECT 0 6.755 0.070 7.105 ;
    RECT 0 7.175 0.070 7.525 ;
    RECT 0 7.595 0.070 7.945 ;
    RECT 0 8.015 0.070 8.365 ;
    RECT 0 8.435 0.070 8.785 ;
    RECT 0 8.855 0.070 9.205 ;
    RECT 0 9.275 0.070 9.625 ;
    RECT 0 9.695 0.070 10.045 ;
    RECT 0 10.115 0.070 10.465 ;
    RECT 0 10.535 0.070 10.885 ;
    RECT 0 10.955 0.070 11.305 ;
    RECT 0 11.375 0.070 11.725 ;
    RECT 0 11.795 0.070 12.145 ;
    RECT 0 12.215 0.070 12.565 ;
    RECT 0 12.635 0.070 12.985 ;
    RECT 0 13.055 0.070 13.405 ;
    RECT 0 13.475 0.070 13.825 ;
    RECT 0 13.895 0.070 14.245 ;
    RECT 0 14.315 0.070 14.665 ;
    RECT 0 14.735 0.070 15.085 ;
    RECT 0 15.155 0.070 15.505 ;
    RECT 0 15.575 0.070 15.925 ;
    RECT 0 15.995 0.070 16.345 ;
    RECT 0 16.415 0.070 16.765 ;
    RECT 0 16.835 0.070 17.185 ;
    RECT 0 17.255 0.070 17.605 ;
    RECT 0 17.675 0.070 18.025 ;
    RECT 0 18.095 0.070 18.445 ;
    RECT 0 18.515 0.070 18.865 ;
    RECT 0 18.935 0.070 19.285 ;
    RECT 0 19.355 0.070 19.705 ;
    RECT 0 19.775 0.070 20.125 ;
    RECT 0 20.195 0.070 20.545 ;
    RECT 0 20.615 0.070 20.965 ;
    RECT 0 21.035 0.070 21.385 ;
    RECT 0 21.455 0.070 21.805 ;
    RECT 0 21.875 0.070 22.225 ;
    RECT 0 22.295 0.070 22.645 ;
    RECT 0 22.715 0.070 23.065 ;
    RECT 0 23.135 0.070 23.485 ;
    RECT 0 23.555 0.070 23.905 ;
    RECT 0 23.975 0.070 24.325 ;
    RECT 0 24.395 0.070 24.745 ;
    RECT 0 24.815 0.070 25.165 ;
    RECT 0 25.235 0.070 25.585 ;
    RECT 0 25.655 0.070 26.005 ;
    RECT 0 26.075 0.070 26.425 ;
    RECT 0 26.495 0.070 26.845 ;
    RECT 0 26.915 0.070 27.265 ;
    RECT 0 27.335 0.070 27.685 ;
    RECT 0 27.755 0.070 28.105 ;
    RECT 0 28.175 0.070 28.525 ;
    RECT 0 28.595 0.070 31.885 ;
    RECT 0 31.955 0.070 32.305 ;
    RECT 0 32.375 0.070 32.725 ;
    RECT 0 32.795 0.070 33.145 ;
    RECT 0 33.215 0.070 33.565 ;
    RECT 0 33.635 0.070 33.985 ;
    RECT 0 34.055 0.070 34.405 ;
    RECT 0 34.475 0.070 34.825 ;
    RECT 0 34.895 0.070 35.245 ;
    RECT 0 35.315 0.070 35.665 ;
    RECT 0 35.735 0.070 36.085 ;
    RECT 0 36.155 0.070 36.505 ;
    RECT 0 36.575 0.070 36.925 ;
    RECT 0 36.995 0.070 37.345 ;
    RECT 0 37.415 0.070 37.765 ;
    RECT 0 37.835 0.070 38.185 ;
    RECT 0 38.255 0.070 38.605 ;
    RECT 0 38.675 0.070 39.025 ;
    RECT 0 39.095 0.070 39.445 ;
    RECT 0 39.515 0.070 39.865 ;
    RECT 0 39.935 0.070 40.285 ;
    RECT 0 40.355 0.070 40.705 ;
    RECT 0 40.775 0.070 41.125 ;
    RECT 0 41.195 0.070 41.545 ;
    RECT 0 41.615 0.070 41.965 ;
    RECT 0 42.035 0.070 42.385 ;
    RECT 0 42.455 0.070 42.805 ;
    RECT 0 42.875 0.070 43.225 ;
    RECT 0 43.295 0.070 43.645 ;
    RECT 0 43.715 0.070 44.065 ;
    RECT 0 44.135 0.070 44.485 ;
    RECT 0 44.555 0.070 44.905 ;
    RECT 0 44.975 0.070 45.325 ;
    RECT 0 45.395 0.070 45.745 ;
    RECT 0 45.815 0.070 46.165 ;
    RECT 0 46.235 0.070 46.585 ;
    RECT 0 46.655 0.070 47.005 ;
    RECT 0 47.075 0.070 47.425 ;
    RECT 0 47.495 0.070 47.845 ;
    RECT 0 47.915 0.070 48.265 ;
    RECT 0 48.335 0.070 48.685 ;
    RECT 0 48.755 0.070 49.105 ;
    RECT 0 49.175 0.070 49.525 ;
    RECT 0 49.595 0.070 49.945 ;
    RECT 0 50.015 0.070 50.365 ;
    RECT 0 50.435 0.070 50.785 ;
    RECT 0 50.855 0.070 51.205 ;
    RECT 0 51.275 0.070 51.625 ;
    RECT 0 51.695 0.070 52.045 ;
    RECT 0 52.115 0.070 52.465 ;
    RECT 0 52.535 0.070 52.885 ;
    RECT 0 52.955 0.070 53.305 ;
    RECT 0 53.375 0.070 53.725 ;
    RECT 0 53.795 0.070 54.145 ;
    RECT 0 54.215 0.070 54.565 ;
    RECT 0 54.635 0.070 54.985 ;
    RECT 0 55.055 0.070 55.405 ;
    RECT 0 55.475 0.070 55.825 ;
    RECT 0 55.895 0.070 56.245 ;
    RECT 0 56.315 0.070 56.665 ;
    RECT 0 56.735 0.070 57.085 ;
    RECT 0 57.155 0.070 57.505 ;
    RECT 0 57.575 0.070 57.925 ;
    RECT 0 57.995 0.070 58.345 ;
    RECT 0 58.415 0.070 61.705 ;
    RECT 0 61.775 0.070 62.125 ;
    RECT 0 62.195 0.070 62.545 ;
    RECT 0 62.615 0.070 62.965 ;
    RECT 0 63.035 0.070 63.385 ;
    RECT 0 63.455 0.070 63.805 ;
    RECT 0 63.875 0.070 64.225 ;
    RECT 0 64.295 0.070 64.645 ;
    RECT 0 64.715 0.070 65.065 ;
    RECT 0 65.135 0.070 65.485 ;
    RECT 0 65.555 0.070 65.905 ;
    RECT 0 65.975 0.070 66.325 ;
    RECT 0 66.395 0.070 66.745 ;
    RECT 0 66.815 0.070 67.165 ;
    RECT 0 67.235 0.070 67.585 ;
    RECT 0 67.655 0.070 68.005 ;
    RECT 0 68.075 0.070 68.425 ;
    RECT 0 68.495 0.070 68.845 ;
    RECT 0 68.915 0.070 69.265 ;
    RECT 0 69.335 0.070 69.685 ;
    RECT 0 69.755 0.070 70.105 ;
    RECT 0 70.175 0.070 70.525 ;
    RECT 0 70.595 0.070 70.945 ;
    RECT 0 71.015 0.070 71.365 ;
    RECT 0 71.435 0.070 71.785 ;
    RECT 0 71.855 0.070 72.205 ;
    RECT 0 72.275 0.070 72.625 ;
    RECT 0 72.695 0.070 73.045 ;
    RECT 0 73.115 0.070 73.465 ;
    RECT 0 73.535 0.070 73.885 ;
    RECT 0 73.955 0.070 74.305 ;
    RECT 0 74.375 0.070 74.725 ;
    RECT 0 74.795 0.070 75.145 ;
    RECT 0 75.215 0.070 75.565 ;
    RECT 0 75.635 0.070 75.985 ;
    RECT 0 76.055 0.070 76.405 ;
    RECT 0 76.475 0.070 76.825 ;
    RECT 0 76.895 0.070 77.245 ;
    RECT 0 77.315 0.070 77.665 ;
    RECT 0 77.735 0.070 78.085 ;
    RECT 0 78.155 0.070 78.505 ;
    RECT 0 78.575 0.070 78.925 ;
    RECT 0 78.995 0.070 79.345 ;
    RECT 0 79.415 0.070 79.765 ;
    RECT 0 79.835 0.070 80.185 ;
    RECT 0 80.255 0.070 80.605 ;
    RECT 0 80.675 0.070 81.025 ;
    RECT 0 81.095 0.070 81.445 ;
    RECT 0 81.515 0.070 81.865 ;
    RECT 0 81.935 0.070 82.285 ;
    RECT 0 82.355 0.070 82.705 ;
    RECT 0 82.775 0.070 83.125 ;
    RECT 0 83.195 0.070 83.545 ;
    RECT 0 83.615 0.070 83.965 ;
    RECT 0 84.035 0.070 84.385 ;
    RECT 0 84.455 0.070 84.805 ;
    RECT 0 84.875 0.070 85.225 ;
    RECT 0 85.295 0.070 85.645 ;
    RECT 0 85.715 0.070 86.065 ;
    RECT 0 86.135 0.070 86.485 ;
    RECT 0 86.555 0.070 86.905 ;
    RECT 0 86.975 0.070 87.325 ;
    RECT 0 87.395 0.070 87.745 ;
    RECT 0 87.815 0.070 88.165 ;
    RECT 0 88.235 0.070 91.525 ;
    RECT 0 91.595 0.070 91.945 ;
    RECT 0 92.015 0.070 92.365 ;
    RECT 0 92.435 0.070 92.785 ;
    RECT 0 92.855 0.070 93.205 ;
    RECT 0 93.275 0.070 93.625 ;
    RECT 0 93.695 0.070 96.985 ;
    RECT 0 97.055 0.070 97.405 ;
    RECT 0 97.475 0.070 97.825 ;
    RECT 0 97.895 0.070 102.200 ;
    LAYER metal4 ;
    RECT 0 0 56.050 2.100 ;
    RECT 0 100.100 56.050 102.200 ;
    RECT 0.000 2.100 1.960 100.100 ;
    RECT 2.240 2.100 3.640 100.100 ;
    RECT 3.920 2.100 5.320 100.100 ;
    RECT 5.600 2.100 7.000 100.100 ;
    RECT 7.280 2.100 8.680 100.100 ;
    RECT 8.960 2.100 10.360 100.100 ;
    RECT 10.640 2.100 12.040 100.100 ;
    RECT 12.320 2.100 13.720 100.100 ;
    RECT 14.000 2.100 15.400 100.100 ;
    RECT 15.680 2.100 17.080 100.100 ;
    RECT 17.360 2.100 18.760 100.100 ;
    RECT 19.040 2.100 20.440 100.100 ;
    RECT 20.720 2.100 22.120 100.100 ;
    RECT 22.400 2.100 23.800 100.100 ;
    RECT 24.080 2.100 25.480 100.100 ;
    RECT 25.760 2.100 27.160 100.100 ;
    RECT 27.440 2.100 28.840 100.100 ;
    RECT 29.120 2.100 30.520 100.100 ;
    RECT 30.800 2.100 32.200 100.100 ;
    RECT 32.480 2.100 33.880 100.100 ;
    RECT 34.160 2.100 35.560 100.100 ;
    RECT 35.840 2.100 37.240 100.100 ;
    RECT 37.520 2.100 38.920 100.100 ;
    RECT 39.200 2.100 40.600 100.100 ;
    RECT 40.880 2.100 42.280 100.100 ;
    RECT 42.560 2.100 43.960 100.100 ;
    RECT 44.240 2.100 45.640 100.100 ;
    RECT 45.920 2.100 47.320 100.100 ;
    RECT 47.600 2.100 49.000 100.100 ;
    RECT 49.280 2.100 50.680 100.100 ;
    RECT 50.960 2.100 52.360 100.100 ;
    RECT 52.640 2.100 56.050 100.100 ;
    LAYER OVERLAP ;
    RECT 0 0 56.050 102.200 ;
  END
END fakeram45_64x64

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_64x62
  FOREIGN fakeram45_64x62 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 56.050 BY 102.200 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.785 0.070 8.855 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.985 0.070 13.055 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.505 0.070 15.575 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.345 0.070 16.415 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.185 0.070 17.255 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.605 0.070 17.675 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.025 0.070 18.095 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.545 0.070 20.615 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.225 0.070 22.295 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.905 0.070 23.975 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.425 0.070 26.495 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.685 0.070 27.755 ;
    END
  END w_mask_in[61]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.675 0.070 31.745 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.095 0.070 32.165 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.515 0.070 32.585 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.935 0.070 33.005 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.355 0.070 33.425 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.775 0.070 33.845 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.195 0.070 34.265 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.615 0.070 34.685 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.035 0.070 35.105 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.455 0.070 35.525 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.875 0.070 35.945 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.295 0.070 36.365 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.715 0.070 36.785 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.135 0.070 37.205 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.555 0.070 37.625 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.975 0.070 38.045 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.395 0.070 38.465 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.815 0.070 38.885 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.235 0.070 39.305 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.655 0.070 39.725 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.075 0.070 40.145 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.495 0.070 40.565 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.915 0.070 40.985 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.335 0.070 41.405 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.755 0.070 41.825 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.175 0.070 42.245 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.595 0.070 42.665 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.015 0.070 43.085 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.435 0.070 43.505 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.855 0.070 43.925 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.275 0.070 44.345 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.695 0.070 44.765 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.115 0.070 45.185 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.535 0.070 45.605 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.955 0.070 46.025 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.375 0.070 46.445 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.795 0.070 46.865 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.215 0.070 47.285 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.635 0.070 47.705 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.055 0.070 48.125 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.475 0.070 48.545 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.895 0.070 48.965 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.315 0.070 49.385 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.735 0.070 49.805 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.155 0.070 50.225 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.575 0.070 50.645 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.995 0.070 51.065 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.415 0.070 51.485 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.835 0.070 51.905 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.255 0.070 52.325 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.675 0.070 52.745 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.095 0.070 53.165 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.515 0.070 53.585 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.935 0.070 54.005 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.355 0.070 54.425 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.775 0.070 54.845 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.195 0.070 55.265 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.615 0.070 55.685 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.035 0.070 56.105 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.455 0.070 56.525 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.875 0.070 56.945 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.295 0.070 57.365 ;
    END
  END rd_out[61]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.285 0.070 61.355 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.705 0.070 61.775 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.125 0.070 62.195 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.545 0.070 62.615 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.965 0.070 63.035 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.385 0.070 63.455 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 63.805 0.070 63.875 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.225 0.070 64.295 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.645 0.070 64.715 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.065 0.070 65.135 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.485 0.070 65.555 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.905 0.070 65.975 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.325 0.070 66.395 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.745 0.070 66.815 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.165 0.070 67.235 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.585 0.070 67.655 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.005 0.070 68.075 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.425 0.070 68.495 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.845 0.070 68.915 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.265 0.070 69.335 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.685 0.070 69.755 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.105 0.070 70.175 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.945 0.070 71.015 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.785 0.070 71.855 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.205 0.070 72.275 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.625 0.070 72.695 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.465 0.070 73.535 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.305 0.070 74.375 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.725 0.070 74.795 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.145 0.070 75.215 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.405 0.070 76.475 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.825 0.070 76.895 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.245 0.070 77.315 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.665 0.070 77.735 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.085 0.070 78.155 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.505 0.070 78.575 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.925 0.070 78.995 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.345 0.070 79.415 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.185 0.070 80.255 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.605 0.070 80.675 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.025 0.070 81.095 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.445 0.070 81.515 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.285 0.070 82.355 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.705 0.070 82.775 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.125 0.070 83.195 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.545 0.070 83.615 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.965 0.070 84.035 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.385 0.070 84.455 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.225 0.070 85.295 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.065 0.070 86.135 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.485 0.070 86.555 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.905 0.070 86.975 ;
    END
  END wd_in[61]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.895 0.070 90.965 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.315 0.070 91.385 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.735 0.070 91.805 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.155 0.070 92.225 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.575 0.070 92.645 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.995 0.070 93.065 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.985 0.070 97.055 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.405 0.070 97.475 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 97.825 0.070 97.895 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 100.100 ;
      RECT 5.320 2.100 5.600 100.100 ;
      RECT 8.680 2.100 8.960 100.100 ;
      RECT 12.040 2.100 12.320 100.100 ;
      RECT 15.400 2.100 15.680 100.100 ;
      RECT 18.760 2.100 19.040 100.100 ;
      RECT 22.120 2.100 22.400 100.100 ;
      RECT 25.480 2.100 25.760 100.100 ;
      RECT 28.840 2.100 29.120 100.100 ;
      RECT 32.200 2.100 32.480 100.100 ;
      RECT 35.560 2.100 35.840 100.100 ;
      RECT 38.920 2.100 39.200 100.100 ;
      RECT 42.280 2.100 42.560 100.100 ;
      RECT 45.640 2.100 45.920 100.100 ;
      RECT 49.000 2.100 49.280 100.100 ;
      RECT 52.360 2.100 52.640 100.100 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 100.100 ;
      RECT 7.000 2.100 7.280 100.100 ;
      RECT 10.360 2.100 10.640 100.100 ;
      RECT 13.720 2.100 14.000 100.100 ;
      RECT 17.080 2.100 17.360 100.100 ;
      RECT 20.440 2.100 20.720 100.100 ;
      RECT 23.800 2.100 24.080 100.100 ;
      RECT 27.160 2.100 27.440 100.100 ;
      RECT 30.520 2.100 30.800 100.100 ;
      RECT 33.880 2.100 34.160 100.100 ;
      RECT 37.240 2.100 37.520 100.100 ;
      RECT 40.600 2.100 40.880 100.100 ;
      RECT 43.960 2.100 44.240 100.100 ;
      RECT 47.320 2.100 47.600 100.100 ;
      RECT 50.680 2.100 50.960 100.100 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 56.050 102.200 ;
    LAYER metal2 ;
    RECT 0 0 56.050 102.200 ;
    LAYER metal3 ;
    RECT 0.070 0 56.050 102.200 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.485 ;
    RECT 0 2.555 0.070 2.905 ;
    RECT 0 2.975 0.070 3.325 ;
    RECT 0 3.395 0.070 3.745 ;
    RECT 0 3.815 0.070 4.165 ;
    RECT 0 4.235 0.070 4.585 ;
    RECT 0 4.655 0.070 5.005 ;
    RECT 0 5.075 0.070 5.425 ;
    RECT 0 5.495 0.070 5.845 ;
    RECT 0 5.915 0.070 6.265 ;
    RECT 0 6.335 0.070 6.685 ;
    RECT 0 6.755 0.070 7.105 ;
    RECT 0 7.175 0.070 7.525 ;
    RECT 0 7.595 0.070 7.945 ;
    RECT 0 8.015 0.070 8.365 ;
    RECT 0 8.435 0.070 8.785 ;
    RECT 0 8.855 0.070 9.205 ;
    RECT 0 9.275 0.070 9.625 ;
    RECT 0 9.695 0.070 10.045 ;
    RECT 0 10.115 0.070 10.465 ;
    RECT 0 10.535 0.070 10.885 ;
    RECT 0 10.955 0.070 11.305 ;
    RECT 0 11.375 0.070 11.725 ;
    RECT 0 11.795 0.070 12.145 ;
    RECT 0 12.215 0.070 12.565 ;
    RECT 0 12.635 0.070 12.985 ;
    RECT 0 13.055 0.070 13.405 ;
    RECT 0 13.475 0.070 13.825 ;
    RECT 0 13.895 0.070 14.245 ;
    RECT 0 14.315 0.070 14.665 ;
    RECT 0 14.735 0.070 15.085 ;
    RECT 0 15.155 0.070 15.505 ;
    RECT 0 15.575 0.070 15.925 ;
    RECT 0 15.995 0.070 16.345 ;
    RECT 0 16.415 0.070 16.765 ;
    RECT 0 16.835 0.070 17.185 ;
    RECT 0 17.255 0.070 17.605 ;
    RECT 0 17.675 0.070 18.025 ;
    RECT 0 18.095 0.070 18.445 ;
    RECT 0 18.515 0.070 18.865 ;
    RECT 0 18.935 0.070 19.285 ;
    RECT 0 19.355 0.070 19.705 ;
    RECT 0 19.775 0.070 20.125 ;
    RECT 0 20.195 0.070 20.545 ;
    RECT 0 20.615 0.070 20.965 ;
    RECT 0 21.035 0.070 21.385 ;
    RECT 0 21.455 0.070 21.805 ;
    RECT 0 21.875 0.070 22.225 ;
    RECT 0 22.295 0.070 22.645 ;
    RECT 0 22.715 0.070 23.065 ;
    RECT 0 23.135 0.070 23.485 ;
    RECT 0 23.555 0.070 23.905 ;
    RECT 0 23.975 0.070 24.325 ;
    RECT 0 24.395 0.070 24.745 ;
    RECT 0 24.815 0.070 25.165 ;
    RECT 0 25.235 0.070 25.585 ;
    RECT 0 25.655 0.070 26.005 ;
    RECT 0 26.075 0.070 26.425 ;
    RECT 0 26.495 0.070 26.845 ;
    RECT 0 26.915 0.070 27.265 ;
    RECT 0 27.335 0.070 27.685 ;
    RECT 0 27.755 0.070 31.675 ;
    RECT 0 31.745 0.070 32.095 ;
    RECT 0 32.165 0.070 32.515 ;
    RECT 0 32.585 0.070 32.935 ;
    RECT 0 33.005 0.070 33.355 ;
    RECT 0 33.425 0.070 33.775 ;
    RECT 0 33.845 0.070 34.195 ;
    RECT 0 34.265 0.070 34.615 ;
    RECT 0 34.685 0.070 35.035 ;
    RECT 0 35.105 0.070 35.455 ;
    RECT 0 35.525 0.070 35.875 ;
    RECT 0 35.945 0.070 36.295 ;
    RECT 0 36.365 0.070 36.715 ;
    RECT 0 36.785 0.070 37.135 ;
    RECT 0 37.205 0.070 37.555 ;
    RECT 0 37.625 0.070 37.975 ;
    RECT 0 38.045 0.070 38.395 ;
    RECT 0 38.465 0.070 38.815 ;
    RECT 0 38.885 0.070 39.235 ;
    RECT 0 39.305 0.070 39.655 ;
    RECT 0 39.725 0.070 40.075 ;
    RECT 0 40.145 0.070 40.495 ;
    RECT 0 40.565 0.070 40.915 ;
    RECT 0 40.985 0.070 41.335 ;
    RECT 0 41.405 0.070 41.755 ;
    RECT 0 41.825 0.070 42.175 ;
    RECT 0 42.245 0.070 42.595 ;
    RECT 0 42.665 0.070 43.015 ;
    RECT 0 43.085 0.070 43.435 ;
    RECT 0 43.505 0.070 43.855 ;
    RECT 0 43.925 0.070 44.275 ;
    RECT 0 44.345 0.070 44.695 ;
    RECT 0 44.765 0.070 45.115 ;
    RECT 0 45.185 0.070 45.535 ;
    RECT 0 45.605 0.070 45.955 ;
    RECT 0 46.025 0.070 46.375 ;
    RECT 0 46.445 0.070 46.795 ;
    RECT 0 46.865 0.070 47.215 ;
    RECT 0 47.285 0.070 47.635 ;
    RECT 0 47.705 0.070 48.055 ;
    RECT 0 48.125 0.070 48.475 ;
    RECT 0 48.545 0.070 48.895 ;
    RECT 0 48.965 0.070 49.315 ;
    RECT 0 49.385 0.070 49.735 ;
    RECT 0 49.805 0.070 50.155 ;
    RECT 0 50.225 0.070 50.575 ;
    RECT 0 50.645 0.070 50.995 ;
    RECT 0 51.065 0.070 51.415 ;
    RECT 0 51.485 0.070 51.835 ;
    RECT 0 51.905 0.070 52.255 ;
    RECT 0 52.325 0.070 52.675 ;
    RECT 0 52.745 0.070 53.095 ;
    RECT 0 53.165 0.070 53.515 ;
    RECT 0 53.585 0.070 53.935 ;
    RECT 0 54.005 0.070 54.355 ;
    RECT 0 54.425 0.070 54.775 ;
    RECT 0 54.845 0.070 55.195 ;
    RECT 0 55.265 0.070 55.615 ;
    RECT 0 55.685 0.070 56.035 ;
    RECT 0 56.105 0.070 56.455 ;
    RECT 0 56.525 0.070 56.875 ;
    RECT 0 56.945 0.070 57.295 ;
    RECT 0 57.365 0.070 61.285 ;
    RECT 0 61.355 0.070 61.705 ;
    RECT 0 61.775 0.070 62.125 ;
    RECT 0 62.195 0.070 62.545 ;
    RECT 0 62.615 0.070 62.965 ;
    RECT 0 63.035 0.070 63.385 ;
    RECT 0 63.455 0.070 63.805 ;
    RECT 0 63.875 0.070 64.225 ;
    RECT 0 64.295 0.070 64.645 ;
    RECT 0 64.715 0.070 65.065 ;
    RECT 0 65.135 0.070 65.485 ;
    RECT 0 65.555 0.070 65.905 ;
    RECT 0 65.975 0.070 66.325 ;
    RECT 0 66.395 0.070 66.745 ;
    RECT 0 66.815 0.070 67.165 ;
    RECT 0 67.235 0.070 67.585 ;
    RECT 0 67.655 0.070 68.005 ;
    RECT 0 68.075 0.070 68.425 ;
    RECT 0 68.495 0.070 68.845 ;
    RECT 0 68.915 0.070 69.265 ;
    RECT 0 69.335 0.070 69.685 ;
    RECT 0 69.755 0.070 70.105 ;
    RECT 0 70.175 0.070 70.525 ;
    RECT 0 70.595 0.070 70.945 ;
    RECT 0 71.015 0.070 71.365 ;
    RECT 0 71.435 0.070 71.785 ;
    RECT 0 71.855 0.070 72.205 ;
    RECT 0 72.275 0.070 72.625 ;
    RECT 0 72.695 0.070 73.045 ;
    RECT 0 73.115 0.070 73.465 ;
    RECT 0 73.535 0.070 73.885 ;
    RECT 0 73.955 0.070 74.305 ;
    RECT 0 74.375 0.070 74.725 ;
    RECT 0 74.795 0.070 75.145 ;
    RECT 0 75.215 0.070 75.565 ;
    RECT 0 75.635 0.070 75.985 ;
    RECT 0 76.055 0.070 76.405 ;
    RECT 0 76.475 0.070 76.825 ;
    RECT 0 76.895 0.070 77.245 ;
    RECT 0 77.315 0.070 77.665 ;
    RECT 0 77.735 0.070 78.085 ;
    RECT 0 78.155 0.070 78.505 ;
    RECT 0 78.575 0.070 78.925 ;
    RECT 0 78.995 0.070 79.345 ;
    RECT 0 79.415 0.070 79.765 ;
    RECT 0 79.835 0.070 80.185 ;
    RECT 0 80.255 0.070 80.605 ;
    RECT 0 80.675 0.070 81.025 ;
    RECT 0 81.095 0.070 81.445 ;
    RECT 0 81.515 0.070 81.865 ;
    RECT 0 81.935 0.070 82.285 ;
    RECT 0 82.355 0.070 82.705 ;
    RECT 0 82.775 0.070 83.125 ;
    RECT 0 83.195 0.070 83.545 ;
    RECT 0 83.615 0.070 83.965 ;
    RECT 0 84.035 0.070 84.385 ;
    RECT 0 84.455 0.070 84.805 ;
    RECT 0 84.875 0.070 85.225 ;
    RECT 0 85.295 0.070 85.645 ;
    RECT 0 85.715 0.070 86.065 ;
    RECT 0 86.135 0.070 86.485 ;
    RECT 0 86.555 0.070 86.905 ;
    RECT 0 86.975 0.070 90.895 ;
    RECT 0 90.965 0.070 91.315 ;
    RECT 0 91.385 0.070 91.735 ;
    RECT 0 91.805 0.070 92.155 ;
    RECT 0 92.225 0.070 92.575 ;
    RECT 0 92.645 0.070 92.995 ;
    RECT 0 93.065 0.070 96.985 ;
    RECT 0 97.055 0.070 97.405 ;
    RECT 0 97.475 0.070 97.825 ;
    RECT 0 97.895 0.070 102.200 ;
    LAYER metal4 ;
    RECT 0 0 56.050 2.100 ;
    RECT 0 100.100 56.050 102.200 ;
    RECT 0.000 2.100 1.960 100.100 ;
    RECT 2.240 2.100 3.640 100.100 ;
    RECT 3.920 2.100 5.320 100.100 ;
    RECT 5.600 2.100 7.000 100.100 ;
    RECT 7.280 2.100 8.680 100.100 ;
    RECT 8.960 2.100 10.360 100.100 ;
    RECT 10.640 2.100 12.040 100.100 ;
    RECT 12.320 2.100 13.720 100.100 ;
    RECT 14.000 2.100 15.400 100.100 ;
    RECT 15.680 2.100 17.080 100.100 ;
    RECT 17.360 2.100 18.760 100.100 ;
    RECT 19.040 2.100 20.440 100.100 ;
    RECT 20.720 2.100 22.120 100.100 ;
    RECT 22.400 2.100 23.800 100.100 ;
    RECT 24.080 2.100 25.480 100.100 ;
    RECT 25.760 2.100 27.160 100.100 ;
    RECT 27.440 2.100 28.840 100.100 ;
    RECT 29.120 2.100 30.520 100.100 ;
    RECT 30.800 2.100 32.200 100.100 ;
    RECT 32.480 2.100 33.880 100.100 ;
    RECT 34.160 2.100 35.560 100.100 ;
    RECT 35.840 2.100 37.240 100.100 ;
    RECT 37.520 2.100 38.920 100.100 ;
    RECT 39.200 2.100 40.600 100.100 ;
    RECT 40.880 2.100 42.280 100.100 ;
    RECT 42.560 2.100 43.960 100.100 ;
    RECT 44.240 2.100 45.640 100.100 ;
    RECT 45.920 2.100 47.320 100.100 ;
    RECT 47.600 2.100 49.000 100.100 ;
    RECT 49.280 2.100 50.680 100.100 ;
    RECT 50.960 2.100 52.360 100.100 ;
    RECT 52.640 2.100 56.050 100.100 ;
    LAYER OVERLAP ;
    RECT 0 0 56.050 102.200 ;
  END
END fakeram45_64x62

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_64x32
  FOREIGN fakeram45_64x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 20.140 BY 61.600 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.785 0.070 8.855 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.985 0.070 13.055 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.235 0.070 18.305 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.655 0.070 18.725 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.075 0.070 19.145 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.495 0.070 19.565 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.915 0.070 19.985 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.335 0.070 20.405 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.755 0.070 20.825 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.175 0.070 21.245 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.595 0.070 21.665 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.015 0.070 22.085 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.435 0.070 22.505 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.855 0.070 22.925 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.275 0.070 23.345 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.695 0.070 23.765 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.115 0.070 24.185 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.535 0.070 24.605 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.955 0.070 25.025 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.375 0.070 25.445 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.795 0.070 25.865 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.215 0.070 26.285 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.635 0.070 26.705 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.055 0.070 27.125 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.475 0.070 27.545 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.895 0.070 27.965 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.315 0.070 28.385 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.735 0.070 28.805 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.155 0.070 29.225 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.575 0.070 29.645 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.995 0.070 30.065 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.415 0.070 30.485 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.835 0.070 30.905 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.255 0.070 31.325 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.825 0.070 34.895 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.505 0.070 36.575 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.185 0.070 38.255 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.325 0.070 45.395 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.745 0.070 45.815 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.585 0.070 46.655 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.575 0.070 50.645 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.995 0.070 51.065 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.415 0.070 51.485 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.835 0.070 51.905 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.255 0.070 52.325 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.675 0.070 52.745 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.825 0.070 55.895 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.665 0.070 56.735 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 59.500 ;
      RECT 5.320 2.100 5.600 59.500 ;
      RECT 8.680 2.100 8.960 59.500 ;
      RECT 12.040 2.100 12.320 59.500 ;
      RECT 15.400 2.100 15.680 59.500 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 59.500 ;
      RECT 7.000 2.100 7.280 59.500 ;
      RECT 10.360 2.100 10.640 59.500 ;
      RECT 13.720 2.100 14.000 59.500 ;
      RECT 17.080 2.100 17.360 59.500 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 20.140 61.600 ;
    LAYER metal2 ;
    RECT 0 0 20.140 61.600 ;
    LAYER metal3 ;
    RECT 0.070 0 20.140 61.600 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.485 ;
    RECT 0 2.555 0.070 2.905 ;
    RECT 0 2.975 0.070 3.325 ;
    RECT 0 3.395 0.070 3.745 ;
    RECT 0 3.815 0.070 4.165 ;
    RECT 0 4.235 0.070 4.585 ;
    RECT 0 4.655 0.070 5.005 ;
    RECT 0 5.075 0.070 5.425 ;
    RECT 0 5.495 0.070 5.845 ;
    RECT 0 5.915 0.070 6.265 ;
    RECT 0 6.335 0.070 6.685 ;
    RECT 0 6.755 0.070 7.105 ;
    RECT 0 7.175 0.070 7.525 ;
    RECT 0 7.595 0.070 7.945 ;
    RECT 0 8.015 0.070 8.365 ;
    RECT 0 8.435 0.070 8.785 ;
    RECT 0 8.855 0.070 9.205 ;
    RECT 0 9.275 0.070 9.625 ;
    RECT 0 9.695 0.070 10.045 ;
    RECT 0 10.115 0.070 10.465 ;
    RECT 0 10.535 0.070 10.885 ;
    RECT 0 10.955 0.070 11.305 ;
    RECT 0 11.375 0.070 11.725 ;
    RECT 0 11.795 0.070 12.145 ;
    RECT 0 12.215 0.070 12.565 ;
    RECT 0 12.635 0.070 12.985 ;
    RECT 0 13.055 0.070 13.405 ;
    RECT 0 13.475 0.070 13.825 ;
    RECT 0 13.895 0.070 14.245 ;
    RECT 0 14.315 0.070 14.665 ;
    RECT 0 14.735 0.070 15.085 ;
    RECT 0 15.155 0.070 18.235 ;
    RECT 0 18.305 0.070 18.655 ;
    RECT 0 18.725 0.070 19.075 ;
    RECT 0 19.145 0.070 19.495 ;
    RECT 0 19.565 0.070 19.915 ;
    RECT 0 19.985 0.070 20.335 ;
    RECT 0 20.405 0.070 20.755 ;
    RECT 0 20.825 0.070 21.175 ;
    RECT 0 21.245 0.070 21.595 ;
    RECT 0 21.665 0.070 22.015 ;
    RECT 0 22.085 0.070 22.435 ;
    RECT 0 22.505 0.070 22.855 ;
    RECT 0 22.925 0.070 23.275 ;
    RECT 0 23.345 0.070 23.695 ;
    RECT 0 23.765 0.070 24.115 ;
    RECT 0 24.185 0.070 24.535 ;
    RECT 0 24.605 0.070 24.955 ;
    RECT 0 25.025 0.070 25.375 ;
    RECT 0 25.445 0.070 25.795 ;
    RECT 0 25.865 0.070 26.215 ;
    RECT 0 26.285 0.070 26.635 ;
    RECT 0 26.705 0.070 27.055 ;
    RECT 0 27.125 0.070 27.475 ;
    RECT 0 27.545 0.070 27.895 ;
    RECT 0 27.965 0.070 28.315 ;
    RECT 0 28.385 0.070 28.735 ;
    RECT 0 28.805 0.070 29.155 ;
    RECT 0 29.225 0.070 29.575 ;
    RECT 0 29.645 0.070 29.995 ;
    RECT 0 30.065 0.070 30.415 ;
    RECT 0 30.485 0.070 30.835 ;
    RECT 0 30.905 0.070 31.255 ;
    RECT 0 31.325 0.070 34.405 ;
    RECT 0 34.475 0.070 34.825 ;
    RECT 0 34.895 0.070 35.245 ;
    RECT 0 35.315 0.070 35.665 ;
    RECT 0 35.735 0.070 36.085 ;
    RECT 0 36.155 0.070 36.505 ;
    RECT 0 36.575 0.070 36.925 ;
    RECT 0 36.995 0.070 37.345 ;
    RECT 0 37.415 0.070 37.765 ;
    RECT 0 37.835 0.070 38.185 ;
    RECT 0 38.255 0.070 38.605 ;
    RECT 0 38.675 0.070 39.025 ;
    RECT 0 39.095 0.070 39.445 ;
    RECT 0 39.515 0.070 39.865 ;
    RECT 0 39.935 0.070 40.285 ;
    RECT 0 40.355 0.070 40.705 ;
    RECT 0 40.775 0.070 41.125 ;
    RECT 0 41.195 0.070 41.545 ;
    RECT 0 41.615 0.070 41.965 ;
    RECT 0 42.035 0.070 42.385 ;
    RECT 0 42.455 0.070 42.805 ;
    RECT 0 42.875 0.070 43.225 ;
    RECT 0 43.295 0.070 43.645 ;
    RECT 0 43.715 0.070 44.065 ;
    RECT 0 44.135 0.070 44.485 ;
    RECT 0 44.555 0.070 44.905 ;
    RECT 0 44.975 0.070 45.325 ;
    RECT 0 45.395 0.070 45.745 ;
    RECT 0 45.815 0.070 46.165 ;
    RECT 0 46.235 0.070 46.585 ;
    RECT 0 46.655 0.070 47.005 ;
    RECT 0 47.075 0.070 47.425 ;
    RECT 0 47.495 0.070 50.575 ;
    RECT 0 50.645 0.070 50.995 ;
    RECT 0 51.065 0.070 51.415 ;
    RECT 0 51.485 0.070 51.835 ;
    RECT 0 51.905 0.070 52.255 ;
    RECT 0 52.325 0.070 52.675 ;
    RECT 0 52.745 0.070 55.825 ;
    RECT 0 55.895 0.070 56.245 ;
    RECT 0 56.315 0.070 56.665 ;
    RECT 0 56.735 0.070 61.600 ;
    LAYER metal4 ;
    RECT 0 0 20.140 2.100 ;
    RECT 0 59.500 20.140 61.600 ;
    RECT 0.000 2.100 1.960 59.500 ;
    RECT 2.240 2.100 3.640 59.500 ;
    RECT 3.920 2.100 5.320 59.500 ;
    RECT 5.600 2.100 7.000 59.500 ;
    RECT 7.280 2.100 8.680 59.500 ;
    RECT 8.960 2.100 10.360 59.500 ;
    RECT 10.640 2.100 12.040 59.500 ;
    RECT 12.320 2.100 13.720 59.500 ;
    RECT 14.000 2.100 15.400 59.500 ;
    RECT 15.680 2.100 17.080 59.500 ;
    RECT 17.360 2.100 20.140 59.500 ;
    LAYER OVERLAP ;
    RECT 0 0 20.140 61.600 ;
  END
END fakeram45_64x32

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_64x21
  FOREIGN fakeram45_64x21 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 15.770 BY 60.200 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.695 0.070 2.765 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.955 0.070 4.025 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.215 0.070 5.285 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.475 0.070 6.545 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.735 0.070 7.805 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.995 0.070 9.065 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.255 0.070 10.325 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.515 0.070 11.585 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.775 0.070 12.845 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.035 0.070 14.105 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[20]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.185 0.070 17.255 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.815 0.070 17.885 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.075 0.070 19.145 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.335 0.070 20.405 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.595 0.070 21.665 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.225 0.070 22.295 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.855 0.070 22.925 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.115 0.070 24.185 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.375 0.070 25.445 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.635 0.070 26.705 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.895 0.070 27.965 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.155 0.070 29.225 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.785 0.070 29.855 ;
    END
  END rd_out[20]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.305 0.070 32.375 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.935 0.070 33.005 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.195 0.070 34.265 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.825 0.070 34.895 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.455 0.070 35.525 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.715 0.070 36.785 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.975 0.070 38.045 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.235 0.070 39.305 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.495 0.070 40.565 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.755 0.070 41.825 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.015 0.070 43.085 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.275 0.070 44.345 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END wd_in[20]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.055 0.070 48.125 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.315 0.070 49.385 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.945 0.070 50.015 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.575 0.070 50.645 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.095 0.070 53.165 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.355 0.070 54.425 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 58.100 ;
      RECT 5.320 2.100 5.600 58.100 ;
      RECT 8.680 2.100 8.960 58.100 ;
      RECT 12.040 2.100 12.320 58.100 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 58.100 ;
      RECT 7.000 2.100 7.280 58.100 ;
      RECT 10.360 2.100 10.640 58.100 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 15.770 60.200 ;
    LAYER metal2 ;
    RECT 0 0 15.770 60.200 ;
    LAYER metal3 ;
    RECT 0.070 0 15.770 60.200 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.695 ;
    RECT 0 2.765 0.070 3.325 ;
    RECT 0 3.395 0.070 3.955 ;
    RECT 0 4.025 0.070 4.585 ;
    RECT 0 4.655 0.070 5.215 ;
    RECT 0 5.285 0.070 5.845 ;
    RECT 0 5.915 0.070 6.475 ;
    RECT 0 6.545 0.070 7.105 ;
    RECT 0 7.175 0.070 7.735 ;
    RECT 0 7.805 0.070 8.365 ;
    RECT 0 8.435 0.070 8.995 ;
    RECT 0 9.065 0.070 9.625 ;
    RECT 0 9.695 0.070 10.255 ;
    RECT 0 10.325 0.070 10.885 ;
    RECT 0 10.955 0.070 11.515 ;
    RECT 0 11.585 0.070 12.145 ;
    RECT 0 12.215 0.070 12.775 ;
    RECT 0 12.845 0.070 13.405 ;
    RECT 0 13.475 0.070 14.035 ;
    RECT 0 14.105 0.070 14.665 ;
    RECT 0 14.735 0.070 17.185 ;
    RECT 0 17.255 0.070 17.815 ;
    RECT 0 17.885 0.070 18.445 ;
    RECT 0 18.515 0.070 19.075 ;
    RECT 0 19.145 0.070 19.705 ;
    RECT 0 19.775 0.070 20.335 ;
    RECT 0 20.405 0.070 20.965 ;
    RECT 0 21.035 0.070 21.595 ;
    RECT 0 21.665 0.070 22.225 ;
    RECT 0 22.295 0.070 22.855 ;
    RECT 0 22.925 0.070 23.485 ;
    RECT 0 23.555 0.070 24.115 ;
    RECT 0 24.185 0.070 24.745 ;
    RECT 0 24.815 0.070 25.375 ;
    RECT 0 25.445 0.070 26.005 ;
    RECT 0 26.075 0.070 26.635 ;
    RECT 0 26.705 0.070 27.265 ;
    RECT 0 27.335 0.070 27.895 ;
    RECT 0 27.965 0.070 28.525 ;
    RECT 0 28.595 0.070 29.155 ;
    RECT 0 29.225 0.070 29.785 ;
    RECT 0 29.855 0.070 32.305 ;
    RECT 0 32.375 0.070 32.935 ;
    RECT 0 33.005 0.070 33.565 ;
    RECT 0 33.635 0.070 34.195 ;
    RECT 0 34.265 0.070 34.825 ;
    RECT 0 34.895 0.070 35.455 ;
    RECT 0 35.525 0.070 36.085 ;
    RECT 0 36.155 0.070 36.715 ;
    RECT 0 36.785 0.070 37.345 ;
    RECT 0 37.415 0.070 37.975 ;
    RECT 0 38.045 0.070 38.605 ;
    RECT 0 38.675 0.070 39.235 ;
    RECT 0 39.305 0.070 39.865 ;
    RECT 0 39.935 0.070 40.495 ;
    RECT 0 40.565 0.070 41.125 ;
    RECT 0 41.195 0.070 41.755 ;
    RECT 0 41.825 0.070 42.385 ;
    RECT 0 42.455 0.070 43.015 ;
    RECT 0 43.085 0.070 43.645 ;
    RECT 0 43.715 0.070 44.275 ;
    RECT 0 44.345 0.070 44.905 ;
    RECT 0 44.975 0.070 47.425 ;
    RECT 0 47.495 0.070 48.055 ;
    RECT 0 48.125 0.070 48.685 ;
    RECT 0 48.755 0.070 49.315 ;
    RECT 0 49.385 0.070 49.945 ;
    RECT 0 50.015 0.070 50.575 ;
    RECT 0 50.645 0.070 53.095 ;
    RECT 0 53.165 0.070 53.725 ;
    RECT 0 53.795 0.070 54.355 ;
    RECT 0 54.425 0.070 60.200 ;
    LAYER metal4 ;
    RECT 0 0 15.770 2.100 ;
    RECT 0 58.100 15.770 60.200 ;
    RECT 0.000 2.100 1.960 58.100 ;
    RECT 2.240 2.100 3.640 58.100 ;
    RECT 3.920 2.100 5.320 58.100 ;
    RECT 5.600 2.100 7.000 58.100 ;
    RECT 7.280 2.100 8.680 58.100 ;
    RECT 8.960 2.100 10.360 58.100 ;
    RECT 10.640 2.100 12.040 58.100 ;
    RECT 12.320 2.100 15.770 58.100 ;
    LAYER OVERLAP ;
    RECT 0 0 15.770 60.200 ;
  END
END fakeram45_64x21

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_64x15
  FOREIGN fakeram45_64x15 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 11.210 BY 58.800 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.785 0.070 8.855 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.985 0.070 13.055 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[14]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.135 0.070 16.205 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.975 0.070 17.045 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.815 0.070 17.885 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.655 0.070 18.725 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.495 0.070 19.565 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.335 0.070 20.405 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.175 0.070 21.245 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.015 0.070 22.085 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.855 0.070 22.925 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.695 0.070 23.765 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.535 0.070 24.605 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.375 0.070 25.445 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.215 0.070 26.285 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.055 0.070 27.125 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.895 0.070 27.965 ;
    END
  END rd_out[14]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.205 0.070 30.275 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.045 0.070 31.115 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.885 0.070 31.955 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END wd_in[14]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.275 0.070 44.345 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.115 0.070 45.185 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.955 0.070 46.025 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.795 0.070 46.865 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.635 0.070 47.705 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.475 0.070 48.545 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.785 0.070 50.855 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.625 0.070 51.695 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 56.700 ;
      RECT 5.320 2.100 5.600 56.700 ;
      RECT 8.680 2.100 8.960 56.700 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 56.700 ;
      RECT 7.000 2.100 7.280 56.700 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 11.210 58.800 ;
    LAYER metal2 ;
    RECT 0 0 11.210 58.800 ;
    LAYER metal3 ;
    RECT 0.070 0 11.210 58.800 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.905 ;
    RECT 0 2.975 0.070 3.745 ;
    RECT 0 3.815 0.070 4.585 ;
    RECT 0 4.655 0.070 5.425 ;
    RECT 0 5.495 0.070 6.265 ;
    RECT 0 6.335 0.070 7.105 ;
    RECT 0 7.175 0.070 7.945 ;
    RECT 0 8.015 0.070 8.785 ;
    RECT 0 8.855 0.070 9.625 ;
    RECT 0 9.695 0.070 10.465 ;
    RECT 0 10.535 0.070 11.305 ;
    RECT 0 11.375 0.070 12.145 ;
    RECT 0 12.215 0.070 12.985 ;
    RECT 0 13.055 0.070 13.825 ;
    RECT 0 13.895 0.070 16.135 ;
    RECT 0 16.205 0.070 16.975 ;
    RECT 0 17.045 0.070 17.815 ;
    RECT 0 17.885 0.070 18.655 ;
    RECT 0 18.725 0.070 19.495 ;
    RECT 0 19.565 0.070 20.335 ;
    RECT 0 20.405 0.070 21.175 ;
    RECT 0 21.245 0.070 22.015 ;
    RECT 0 22.085 0.070 22.855 ;
    RECT 0 22.925 0.070 23.695 ;
    RECT 0 23.765 0.070 24.535 ;
    RECT 0 24.605 0.070 25.375 ;
    RECT 0 25.445 0.070 26.215 ;
    RECT 0 26.285 0.070 27.055 ;
    RECT 0 27.125 0.070 27.895 ;
    RECT 0 27.965 0.070 30.205 ;
    RECT 0 30.275 0.070 31.045 ;
    RECT 0 31.115 0.070 31.885 ;
    RECT 0 31.955 0.070 32.725 ;
    RECT 0 32.795 0.070 33.565 ;
    RECT 0 33.635 0.070 34.405 ;
    RECT 0 34.475 0.070 35.245 ;
    RECT 0 35.315 0.070 36.085 ;
    RECT 0 36.155 0.070 36.925 ;
    RECT 0 36.995 0.070 37.765 ;
    RECT 0 37.835 0.070 38.605 ;
    RECT 0 38.675 0.070 39.445 ;
    RECT 0 39.515 0.070 40.285 ;
    RECT 0 40.355 0.070 41.125 ;
    RECT 0 41.195 0.070 41.965 ;
    RECT 0 42.035 0.070 44.275 ;
    RECT 0 44.345 0.070 45.115 ;
    RECT 0 45.185 0.070 45.955 ;
    RECT 0 46.025 0.070 46.795 ;
    RECT 0 46.865 0.070 47.635 ;
    RECT 0 47.705 0.070 48.475 ;
    RECT 0 48.545 0.070 50.785 ;
    RECT 0 50.855 0.070 51.625 ;
    RECT 0 51.695 0.070 52.465 ;
    RECT 0 52.535 0.070 58.800 ;
    LAYER metal4 ;
    RECT 0 0 11.210 2.100 ;
    RECT 0 56.700 11.210 58.800 ;
    RECT 0.000 2.100 1.960 56.700 ;
    RECT 2.240 2.100 3.640 56.700 ;
    RECT 3.920 2.100 5.320 56.700 ;
    RECT 5.600 2.100 7.000 56.700 ;
    RECT 7.280 2.100 8.680 56.700 ;
    RECT 8.960 2.100 11.210 56.700 ;
    LAYER OVERLAP ;
    RECT 0 0 11.210 58.800 ;
  END
END fakeram45_64x15

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_64x7
  FOREIGN fakeram45_64x7 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 10.640 BY 36.400 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.115 0.070 3.185 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.215 0.070 5.285 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.315 0.070 7.385 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[6]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.575 0.070 8.645 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.675 0.070 10.745 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.775 0.070 12.845 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.875 0.070 14.945 ;
    END
  END rd_out[6]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.135 0.070 16.205 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.185 0.070 17.255 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.235 0.070 18.305 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.335 0.070 20.405 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END wd_in[6]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.595 0.070 21.665 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.695 0.070 23.765 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.795 0.070 25.865 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.055 0.070 27.125 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.105 0.070 28.175 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.155 0.070 29.225 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 34.300 ;
      RECT 5.320 2.100 5.600 34.300 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 34.300 ;
      RECT 7.000 2.100 7.280 34.300 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 10.640 36.400 ;
    LAYER metal2 ;
    RECT 0 0 10.640 36.400 ;
    LAYER metal3 ;
    RECT 0.070 0 10.640 36.400 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 3.115 ;
    RECT 0 3.185 0.070 4.165 ;
    RECT 0 4.235 0.070 5.215 ;
    RECT 0 5.285 0.070 6.265 ;
    RECT 0 6.335 0.070 7.315 ;
    RECT 0 7.385 0.070 8.365 ;
    RECT 0 8.435 0.070 8.575 ;
    RECT 0 8.645 0.070 9.625 ;
    RECT 0 9.695 0.070 10.675 ;
    RECT 0 10.745 0.070 11.725 ;
    RECT 0 11.795 0.070 12.775 ;
    RECT 0 12.845 0.070 13.825 ;
    RECT 0 13.895 0.070 14.875 ;
    RECT 0 14.945 0.070 15.085 ;
    RECT 0 15.155 0.070 16.135 ;
    RECT 0 16.205 0.070 17.185 ;
    RECT 0 17.255 0.070 18.235 ;
    RECT 0 18.305 0.070 19.285 ;
    RECT 0 19.355 0.070 20.335 ;
    RECT 0 20.405 0.070 21.385 ;
    RECT 0 21.455 0.070 21.595 ;
    RECT 0 21.665 0.070 22.645 ;
    RECT 0 22.715 0.070 23.695 ;
    RECT 0 23.765 0.070 24.745 ;
    RECT 0 24.815 0.070 25.795 ;
    RECT 0 25.865 0.070 26.845 ;
    RECT 0 26.915 0.070 27.055 ;
    RECT 0 27.125 0.070 28.105 ;
    RECT 0 28.175 0.070 29.155 ;
    RECT 0 29.225 0.070 36.400 ;
    LAYER metal4 ;
    RECT 0 0 10.640 2.100 ;
    RECT 0 34.300 10.640 36.400 ;
    RECT 0.000 2.100 1.960 34.300 ;
    RECT 2.240 2.100 3.640 34.300 ;
    RECT 3.920 2.100 5.320 34.300 ;
    RECT 5.600 2.100 7.000 34.300 ;
    RECT 7.280 2.100 10.640 34.300 ;
    LAYER OVERLAP ;
    RECT 0 0 10.640 36.400 ;
  END
END fakeram45_64x7

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_32x64
  FOREIGN fakeram45_32x64 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 36.860 BY 47.600 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.275 0.070 2.345 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.695 0.070 2.765 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.115 0.070 3.185 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.535 0.070 3.605 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.955 0.070 4.025 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.375 0.070 4.445 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.795 0.070 4.865 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.215 0.070 5.285 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.635 0.070 5.705 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.055 0.070 6.125 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.475 0.070 6.545 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.895 0.070 6.965 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.315 0.070 7.385 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.735 0.070 7.805 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.155 0.070 8.225 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.575 0.070 8.645 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.785 0.070 8.855 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.995 0.070 9.065 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.415 0.070 9.485 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.625 0.070 9.695 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.835 0.070 9.905 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.255 0.070 10.325 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.675 0.070 10.745 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.095 0.070 11.165 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.515 0.070 11.585 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.935 0.070 12.005 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.355 0.070 12.425 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.775 0.070 12.845 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.985 0.070 13.055 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.195 0.070 13.265 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.615 0.070 13.685 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.035 0.070 14.105 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.455 0.070 14.525 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.875 0.070 14.945 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.295 0.070 15.365 ;
    END
  END w_mask_in[63]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.505 0.070 15.575 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.715 0.070 15.785 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.135 0.070 16.205 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.345 0.070 16.415 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.555 0.070 16.625 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.975 0.070 17.045 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.185 0.070 17.255 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.395 0.070 17.465 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.605 0.070 17.675 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.815 0.070 17.885 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.025 0.070 18.095 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.235 0.070 18.305 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.655 0.070 18.725 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.075 0.070 19.145 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.495 0.070 19.565 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.915 0.070 19.985 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.335 0.070 20.405 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.545 0.070 20.615 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.755 0.070 20.825 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.175 0.070 21.245 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.595 0.070 21.665 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.015 0.070 22.085 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.225 0.070 22.295 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.435 0.070 22.505 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.855 0.070 22.925 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.275 0.070 23.345 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.695 0.070 23.765 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.905 0.070 23.975 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.115 0.070 24.185 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.535 0.070 24.605 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.955 0.070 25.025 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.375 0.070 25.445 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.795 0.070 25.865 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.215 0.070 26.285 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.425 0.070 26.495 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.635 0.070 26.705 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.055 0.070 27.125 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.475 0.070 27.545 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.685 0.070 27.755 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.895 0.070 27.965 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.105 0.070 28.175 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.315 0.070 28.385 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.735 0.070 28.805 ;
    END
  END rd_out[63]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.945 0.070 29.015 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.155 0.070 29.225 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.365 0.070 29.435 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.575 0.070 29.645 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.785 0.070 29.855 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.995 0.070 30.065 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.205 0.070 30.275 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.415 0.070 30.485 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.625 0.070 30.695 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.835 0.070 30.905 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.045 0.070 31.115 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.255 0.070 31.325 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.465 0.070 31.535 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.675 0.070 31.745 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.885 0.070 31.955 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.095 0.070 32.165 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.305 0.070 32.375 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.515 0.070 32.585 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.725 0.070 32.795 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.935 0.070 33.005 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.145 0.070 33.215 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.355 0.070 33.425 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.565 0.070 33.635 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.775 0.070 33.845 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.985 0.070 34.055 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.195 0.070 34.265 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.615 0.070 34.685 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.825 0.070 34.895 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.035 0.070 35.105 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.455 0.070 35.525 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.875 0.070 35.945 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.295 0.070 36.365 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.505 0.070 36.575 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.715 0.070 36.785 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.135 0.070 37.205 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.555 0.070 37.625 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.975 0.070 38.045 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.185 0.070 38.255 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.395 0.070 38.465 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.815 0.070 38.885 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.235 0.070 39.305 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.655 0.070 39.725 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.075 0.070 40.145 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.495 0.070 40.565 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.915 0.070 40.985 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.335 0.070 41.405 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.755 0.070 41.825 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.175 0.070 42.245 ;
    END
  END wd_in[63]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.595 0.070 42.665 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.015 0.070 43.085 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END addr_in[4]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.435 0.070 43.505 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.855 0.070 43.925 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 45.500 ;
      RECT 5.320 2.100 5.600 45.500 ;
      RECT 8.680 2.100 8.960 45.500 ;
      RECT 12.040 2.100 12.320 45.500 ;
      RECT 15.400 2.100 15.680 45.500 ;
      RECT 18.760 2.100 19.040 45.500 ;
      RECT 22.120 2.100 22.400 45.500 ;
      RECT 25.480 2.100 25.760 45.500 ;
      RECT 28.840 2.100 29.120 45.500 ;
      RECT 32.200 2.100 32.480 45.500 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 45.500 ;
      RECT 7.000 2.100 7.280 45.500 ;
      RECT 10.360 2.100 10.640 45.500 ;
      RECT 13.720 2.100 14.000 45.500 ;
      RECT 17.080 2.100 17.360 45.500 ;
      RECT 20.440 2.100 20.720 45.500 ;
      RECT 23.800 2.100 24.080 45.500 ;
      RECT 27.160 2.100 27.440 45.500 ;
      RECT 30.520 2.100 30.800 45.500 ;
      RECT 33.880 2.100 34.160 45.500 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 36.860 47.600 ;
    LAYER metal2 ;
    RECT 0 0 36.860 47.600 ;
    LAYER metal3 ;
    RECT 0.070 0 36.860 47.600 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.275 ;
    RECT 0 2.345 0.070 2.485 ;
    RECT 0 2.555 0.070 2.695 ;
    RECT 0 2.765 0.070 2.905 ;
    RECT 0 2.975 0.070 3.115 ;
    RECT 0 3.185 0.070 3.325 ;
    RECT 0 3.395 0.070 3.535 ;
    RECT 0 3.605 0.070 3.745 ;
    RECT 0 3.815 0.070 3.955 ;
    RECT 0 4.025 0.070 4.165 ;
    RECT 0 4.235 0.070 4.375 ;
    RECT 0 4.445 0.070 4.585 ;
    RECT 0 4.655 0.070 4.795 ;
    RECT 0 4.865 0.070 5.005 ;
    RECT 0 5.075 0.070 5.215 ;
    RECT 0 5.285 0.070 5.425 ;
    RECT 0 5.495 0.070 5.635 ;
    RECT 0 5.705 0.070 5.845 ;
    RECT 0 5.915 0.070 6.055 ;
    RECT 0 6.125 0.070 6.265 ;
    RECT 0 6.335 0.070 6.475 ;
    RECT 0 6.545 0.070 6.685 ;
    RECT 0 6.755 0.070 6.895 ;
    RECT 0 6.965 0.070 7.105 ;
    RECT 0 7.175 0.070 7.315 ;
    RECT 0 7.385 0.070 7.525 ;
    RECT 0 7.595 0.070 7.735 ;
    RECT 0 7.805 0.070 7.945 ;
    RECT 0 8.015 0.070 8.155 ;
    RECT 0 8.225 0.070 8.365 ;
    RECT 0 8.435 0.070 8.575 ;
    RECT 0 8.645 0.070 8.785 ;
    RECT 0 8.855 0.070 8.995 ;
    RECT 0 9.065 0.070 9.205 ;
    RECT 0 9.275 0.070 9.415 ;
    RECT 0 9.485 0.070 9.625 ;
    RECT 0 9.695 0.070 9.835 ;
    RECT 0 9.905 0.070 10.045 ;
    RECT 0 10.115 0.070 10.255 ;
    RECT 0 10.325 0.070 10.465 ;
    RECT 0 10.535 0.070 10.675 ;
    RECT 0 10.745 0.070 10.885 ;
    RECT 0 10.955 0.070 11.095 ;
    RECT 0 11.165 0.070 11.305 ;
    RECT 0 11.375 0.070 11.515 ;
    RECT 0 11.585 0.070 11.725 ;
    RECT 0 11.795 0.070 11.935 ;
    RECT 0 12.005 0.070 12.145 ;
    RECT 0 12.215 0.070 12.355 ;
    RECT 0 12.425 0.070 12.565 ;
    RECT 0 12.635 0.070 12.775 ;
    RECT 0 12.845 0.070 12.985 ;
    RECT 0 13.055 0.070 13.195 ;
    RECT 0 13.265 0.070 13.405 ;
    RECT 0 13.475 0.070 13.615 ;
    RECT 0 13.685 0.070 13.825 ;
    RECT 0 13.895 0.070 14.035 ;
    RECT 0 14.105 0.070 14.245 ;
    RECT 0 14.315 0.070 14.455 ;
    RECT 0 14.525 0.070 14.665 ;
    RECT 0 14.735 0.070 14.875 ;
    RECT 0 14.945 0.070 15.085 ;
    RECT 0 15.155 0.070 15.295 ;
    RECT 0 15.365 0.070 15.505 ;
    RECT 0 15.575 0.070 15.715 ;
    RECT 0 15.785 0.070 15.925 ;
    RECT 0 15.995 0.070 16.135 ;
    RECT 0 16.205 0.070 16.345 ;
    RECT 0 16.415 0.070 16.555 ;
    RECT 0 16.625 0.070 16.765 ;
    RECT 0 16.835 0.070 16.975 ;
    RECT 0 17.045 0.070 17.185 ;
    RECT 0 17.255 0.070 17.395 ;
    RECT 0 17.465 0.070 17.605 ;
    RECT 0 17.675 0.070 17.815 ;
    RECT 0 17.885 0.070 18.025 ;
    RECT 0 18.095 0.070 18.235 ;
    RECT 0 18.305 0.070 18.445 ;
    RECT 0 18.515 0.070 18.655 ;
    RECT 0 18.725 0.070 18.865 ;
    RECT 0 18.935 0.070 19.075 ;
    RECT 0 19.145 0.070 19.285 ;
    RECT 0 19.355 0.070 19.495 ;
    RECT 0 19.565 0.070 19.705 ;
    RECT 0 19.775 0.070 19.915 ;
    RECT 0 19.985 0.070 20.125 ;
    RECT 0 20.195 0.070 20.335 ;
    RECT 0 20.405 0.070 20.545 ;
    RECT 0 20.615 0.070 20.755 ;
    RECT 0 20.825 0.070 20.965 ;
    RECT 0 21.035 0.070 21.175 ;
    RECT 0 21.245 0.070 21.385 ;
    RECT 0 21.455 0.070 21.595 ;
    RECT 0 21.665 0.070 21.805 ;
    RECT 0 21.875 0.070 22.015 ;
    RECT 0 22.085 0.070 22.225 ;
    RECT 0 22.295 0.070 22.435 ;
    RECT 0 22.505 0.070 22.645 ;
    RECT 0 22.715 0.070 22.855 ;
    RECT 0 22.925 0.070 23.065 ;
    RECT 0 23.135 0.070 23.275 ;
    RECT 0 23.345 0.070 23.485 ;
    RECT 0 23.555 0.070 23.695 ;
    RECT 0 23.765 0.070 23.905 ;
    RECT 0 23.975 0.070 24.115 ;
    RECT 0 24.185 0.070 24.325 ;
    RECT 0 24.395 0.070 24.535 ;
    RECT 0 24.605 0.070 24.745 ;
    RECT 0 24.815 0.070 24.955 ;
    RECT 0 25.025 0.070 25.165 ;
    RECT 0 25.235 0.070 25.375 ;
    RECT 0 25.445 0.070 25.585 ;
    RECT 0 25.655 0.070 25.795 ;
    RECT 0 25.865 0.070 26.005 ;
    RECT 0 26.075 0.070 26.215 ;
    RECT 0 26.285 0.070 26.425 ;
    RECT 0 26.495 0.070 26.635 ;
    RECT 0 26.705 0.070 26.845 ;
    RECT 0 26.915 0.070 27.055 ;
    RECT 0 27.125 0.070 27.265 ;
    RECT 0 27.335 0.070 27.475 ;
    RECT 0 27.545 0.070 27.685 ;
    RECT 0 27.755 0.070 27.895 ;
    RECT 0 27.965 0.070 28.105 ;
    RECT 0 28.175 0.070 28.315 ;
    RECT 0 28.385 0.070 28.525 ;
    RECT 0 28.595 0.070 28.735 ;
    RECT 0 28.805 0.070 28.945 ;
    RECT 0 29.015 0.070 29.155 ;
    RECT 0 29.225 0.070 29.365 ;
    RECT 0 29.435 0.070 29.575 ;
    RECT 0 29.645 0.070 29.785 ;
    RECT 0 29.855 0.070 29.995 ;
    RECT 0 30.065 0.070 30.205 ;
    RECT 0 30.275 0.070 30.415 ;
    RECT 0 30.485 0.070 30.625 ;
    RECT 0 30.695 0.070 30.835 ;
    RECT 0 30.905 0.070 31.045 ;
    RECT 0 31.115 0.070 31.255 ;
    RECT 0 31.325 0.070 31.465 ;
    RECT 0 31.535 0.070 31.675 ;
    RECT 0 31.745 0.070 31.885 ;
    RECT 0 31.955 0.070 32.095 ;
    RECT 0 32.165 0.070 32.305 ;
    RECT 0 32.375 0.070 32.515 ;
    RECT 0 32.585 0.070 32.725 ;
    RECT 0 32.795 0.070 32.935 ;
    RECT 0 33.005 0.070 33.145 ;
    RECT 0 33.215 0.070 33.355 ;
    RECT 0 33.425 0.070 33.565 ;
    RECT 0 33.635 0.070 33.775 ;
    RECT 0 33.845 0.070 33.985 ;
    RECT 0 34.055 0.070 34.195 ;
    RECT 0 34.265 0.070 34.405 ;
    RECT 0 34.475 0.070 34.615 ;
    RECT 0 34.685 0.070 34.825 ;
    RECT 0 34.895 0.070 35.035 ;
    RECT 0 35.105 0.070 35.245 ;
    RECT 0 35.315 0.070 35.455 ;
    RECT 0 35.525 0.070 35.665 ;
    RECT 0 35.735 0.070 35.875 ;
    RECT 0 35.945 0.070 36.085 ;
    RECT 0 36.155 0.070 36.295 ;
    RECT 0 36.365 0.070 36.505 ;
    RECT 0 36.575 0.070 36.715 ;
    RECT 0 36.785 0.070 36.925 ;
    RECT 0 36.995 0.070 37.135 ;
    RECT 0 37.205 0.070 37.345 ;
    RECT 0 37.415 0.070 37.555 ;
    RECT 0 37.625 0.070 37.765 ;
    RECT 0 37.835 0.070 37.975 ;
    RECT 0 38.045 0.070 38.185 ;
    RECT 0 38.255 0.070 38.395 ;
    RECT 0 38.465 0.070 38.605 ;
    RECT 0 38.675 0.070 38.815 ;
    RECT 0 38.885 0.070 39.025 ;
    RECT 0 39.095 0.070 39.235 ;
    RECT 0 39.305 0.070 39.445 ;
    RECT 0 39.515 0.070 39.655 ;
    RECT 0 39.725 0.070 39.865 ;
    RECT 0 39.935 0.070 40.075 ;
    RECT 0 40.145 0.070 40.285 ;
    RECT 0 40.355 0.070 40.495 ;
    RECT 0 40.565 0.070 40.705 ;
    RECT 0 40.775 0.070 40.915 ;
    RECT 0 40.985 0.070 41.125 ;
    RECT 0 41.195 0.070 41.335 ;
    RECT 0 41.405 0.070 41.545 ;
    RECT 0 41.615 0.070 41.755 ;
    RECT 0 41.825 0.070 41.965 ;
    RECT 0 42.035 0.070 42.175 ;
    RECT 0 42.245 0.070 42.385 ;
    RECT 0 42.455 0.070 42.595 ;
    RECT 0 42.665 0.070 42.805 ;
    RECT 0 42.875 0.070 43.015 ;
    RECT 0 43.085 0.070 43.225 ;
    RECT 0 43.295 0.070 43.435 ;
    RECT 0 43.505 0.070 43.645 ;
    RECT 0 43.715 0.070 43.855 ;
    RECT 0 43.925 0.070 47.600 ;
    LAYER metal4 ;
    RECT 0 0 36.860 2.100 ;
    RECT 0 45.500 36.860 47.600 ;
    RECT 0.000 2.100 1.960 45.500 ;
    RECT 2.240 2.100 3.640 45.500 ;
    RECT 3.920 2.100 5.320 45.500 ;
    RECT 5.600 2.100 7.000 45.500 ;
    RECT 7.280 2.100 8.680 45.500 ;
    RECT 8.960 2.100 10.360 45.500 ;
    RECT 10.640 2.100 12.040 45.500 ;
    RECT 12.320 2.100 13.720 45.500 ;
    RECT 14.000 2.100 15.400 45.500 ;
    RECT 15.680 2.100 17.080 45.500 ;
    RECT 17.360 2.100 18.760 45.500 ;
    RECT 19.040 2.100 20.440 45.500 ;
    RECT 20.720 2.100 22.120 45.500 ;
    RECT 22.400 2.100 23.800 45.500 ;
    RECT 24.080 2.100 25.480 45.500 ;
    RECT 25.760 2.100 27.160 45.500 ;
    RECT 27.440 2.100 28.840 45.500 ;
    RECT 29.120 2.100 30.520 45.500 ;
    RECT 30.800 2.100 32.200 45.500 ;
    RECT 32.480 2.100 33.880 45.500 ;
    RECT 34.160 2.100 36.860 45.500 ;
    LAYER OVERLAP ;
    RECT 0 0 36.860 47.600 ;
  END
END fakeram45_32x64

# END LIBRARY
#VERSION 5.7 ;
#BUSBITCHARS "[]" ;
MACRO fakeram45_32x32
  FOREIGN fakeram45_32x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 55.100 BY 33.600 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.275 0.070 2.345 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.695 0.070 2.765 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.905 0.070 2.975 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.115 0.070 3.185 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.535 0.070 3.605 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.745 0.070 3.815 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.955 0.070 4.025 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.375 0.070 4.445 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.585 0.070 4.655 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.795 0.070 4.865 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.215 0.070 5.285 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.425 0.070 5.495 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.635 0.070 5.705 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.055 0.070 6.125 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.475 0.070 6.545 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.895 0.070 6.965 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.105 0.070 7.175 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.315 0.070 7.385 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.735 0.070 7.805 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.155 0.070 8.225 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.575 0.070 8.645 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.675 0.070 10.745 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.095 0.070 11.165 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.305 0.070 11.375 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.515 0.070 11.585 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.935 0.070 12.005 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.145 0.070 12.215 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.355 0.070 12.425 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.775 0.070 12.845 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.985 0.070 13.055 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.195 0.070 13.265 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.615 0.070 13.685 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.035 0.070 14.105 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.455 0.070 14.525 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.875 0.070 14.945 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.295 0.070 15.365 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.505 0.070 15.575 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.715 0.070 15.785 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.135 0.070 16.205 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.345 0.070 16.415 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.555 0.070 16.625 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.975 0.070 17.045 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.075 0.070 19.145 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.495 0.070 19.565 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.915 0.070 19.985 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.335 0.070 20.405 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.545 0.070 20.615 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.755 0.070 20.825 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.175 0.070 21.245 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.385 0.070 21.455 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.595 0.070 21.665 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.015 0.070 22.085 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.225 0.070 22.295 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.435 0.070 22.505 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.855 0.070 22.925 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.275 0.070 23.345 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.695 0.070 23.765 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.905 0.070 23.975 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.115 0.070 24.185 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.535 0.070 24.605 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.745 0.070 24.815 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.955 0.070 25.025 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.375 0.070 25.445 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.475 0.070 27.545 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.685 0.070 27.755 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.895 0.070 27.965 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.105 0.070 28.175 ;
    END
  END addr_in[4]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.995 0.070 30.065 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.205 0.070 30.275 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.415 0.070 30.485 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 31.500 ;
      RECT 5.320 2.100 5.600 31.500 ;
      RECT 8.680 2.100 8.960 31.500 ;
      RECT 12.040 2.100 12.320 31.500 ;
      RECT 15.400 2.100 15.680 31.500 ;
      RECT 18.760 2.100 19.040 31.500 ;
      RECT 22.120 2.100 22.400 31.500 ;
      RECT 25.480 2.100 25.760 31.500 ;
      RECT 28.840 2.100 29.120 31.500 ;
      RECT 32.200 2.100 32.480 31.500 ;
      RECT 35.560 2.100 35.840 31.500 ;
      RECT 38.920 2.100 39.200 31.500 ;
      RECT 42.280 2.100 42.560 31.500 ;
      RECT 45.640 2.100 45.920 31.500 ;
      RECT 49.000 2.100 49.280 31.500 ;
      RECT 52.360 2.100 52.640 31.500 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 31.500 ;
      RECT 7.000 2.100 7.280 31.500 ;
      RECT 10.360 2.100 10.640 31.500 ;
      RECT 13.720 2.100 14.000 31.500 ;
      RECT 17.080 2.100 17.360 31.500 ;
      RECT 20.440 2.100 20.720 31.500 ;
      RECT 23.800 2.100 24.080 31.500 ;
      RECT 27.160 2.100 27.440 31.500 ;
      RECT 30.520 2.100 30.800 31.500 ;
      RECT 33.880 2.100 34.160 31.500 ;
      RECT 37.240 2.100 37.520 31.500 ;
      RECT 40.600 2.100 40.880 31.500 ;
      RECT 43.960 2.100 44.240 31.500 ;
      RECT 47.320 2.100 47.600 31.500 ;
      RECT 50.680 2.100 50.960 31.500 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 55.100 33.600 ;
    LAYER metal2 ;
    RECT 0 0 55.100 33.600 ;
    LAYER metal3 ;
    RECT 0.070 0 55.100 33.600 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 2.275 ;
    RECT 0 2.345 0.070 2.485 ;
    RECT 0 2.555 0.070 2.695 ;
    RECT 0 2.765 0.070 2.905 ;
    RECT 0 2.975 0.070 3.115 ;
    RECT 0 3.185 0.070 3.325 ;
    RECT 0 3.395 0.070 3.535 ;
    RECT 0 3.605 0.070 3.745 ;
    RECT 0 3.815 0.070 3.955 ;
    RECT 0 4.025 0.070 4.165 ;
    RECT 0 4.235 0.070 4.375 ;
    RECT 0 4.445 0.070 4.585 ;
    RECT 0 4.655 0.070 4.795 ;
    RECT 0 4.865 0.070 5.005 ;
    RECT 0 5.075 0.070 5.215 ;
    RECT 0 5.285 0.070 5.425 ;
    RECT 0 5.495 0.070 5.635 ;
    RECT 0 5.705 0.070 5.845 ;
    RECT 0 5.915 0.070 6.055 ;
    RECT 0 6.125 0.070 6.265 ;
    RECT 0 6.335 0.070 6.475 ;
    RECT 0 6.545 0.070 6.685 ;
    RECT 0 6.755 0.070 6.895 ;
    RECT 0 6.965 0.070 7.105 ;
    RECT 0 7.175 0.070 7.315 ;
    RECT 0 7.385 0.070 7.525 ;
    RECT 0 7.595 0.070 7.735 ;
    RECT 0 7.805 0.070 7.945 ;
    RECT 0 8.015 0.070 8.155 ;
    RECT 0 8.225 0.070 8.365 ;
    RECT 0 8.435 0.070 8.575 ;
    RECT 0 8.645 0.070 10.465 ;
    RECT 0 10.535 0.070 10.675 ;
    RECT 0 10.745 0.070 10.885 ;
    RECT 0 10.955 0.070 11.095 ;
    RECT 0 11.165 0.070 11.305 ;
    RECT 0 11.375 0.070 11.515 ;
    RECT 0 11.585 0.070 11.725 ;
    RECT 0 11.795 0.070 11.935 ;
    RECT 0 12.005 0.070 12.145 ;
    RECT 0 12.215 0.070 12.355 ;
    RECT 0 12.425 0.070 12.565 ;
    RECT 0 12.635 0.070 12.775 ;
    RECT 0 12.845 0.070 12.985 ;
    RECT 0 13.055 0.070 13.195 ;
    RECT 0 13.265 0.070 13.405 ;
    RECT 0 13.475 0.070 13.615 ;
    RECT 0 13.685 0.070 13.825 ;
    RECT 0 13.895 0.070 14.035 ;
    RECT 0 14.105 0.070 14.245 ;
    RECT 0 14.315 0.070 14.455 ;
    RECT 0 14.525 0.070 14.665 ;
    RECT 0 14.735 0.070 14.875 ;
    RECT 0 14.945 0.070 15.085 ;
    RECT 0 15.155 0.070 15.295 ;
    RECT 0 15.365 0.070 15.505 ;
    RECT 0 15.575 0.070 15.715 ;
    RECT 0 15.785 0.070 15.925 ;
    RECT 0 15.995 0.070 16.135 ;
    RECT 0 16.205 0.070 16.345 ;
    RECT 0 16.415 0.070 16.555 ;
    RECT 0 16.625 0.070 16.765 ;
    RECT 0 16.835 0.070 16.975 ;
    RECT 0 17.045 0.070 18.865 ;
    RECT 0 18.935 0.070 19.075 ;
    RECT 0 19.145 0.070 19.285 ;
    RECT 0 19.355 0.070 19.495 ;
    RECT 0 19.565 0.070 19.705 ;
    RECT 0 19.775 0.070 19.915 ;
    RECT 0 19.985 0.070 20.125 ;
    RECT 0 20.195 0.070 20.335 ;
    RECT 0 20.405 0.070 20.545 ;
    RECT 0 20.615 0.070 20.755 ;
    RECT 0 20.825 0.070 20.965 ;
    RECT 0 21.035 0.070 21.175 ;
    RECT 0 21.245 0.070 21.385 ;
    RECT 0 21.455 0.070 21.595 ;
    RECT 0 21.665 0.070 21.805 ;
    RECT 0 21.875 0.070 22.015 ;
    RECT 0 22.085 0.070 22.225 ;
    RECT 0 22.295 0.070 22.435 ;
    RECT 0 22.505 0.070 22.645 ;
    RECT 0 22.715 0.070 22.855 ;
    RECT 0 22.925 0.070 23.065 ;
    RECT 0 23.135 0.070 23.275 ;
    RECT 0 23.345 0.070 23.485 ;
    RECT 0 23.555 0.070 23.695 ;
    RECT 0 23.765 0.070 23.905 ;
    RECT 0 23.975 0.070 24.115 ;
    RECT 0 24.185 0.070 24.325 ;
    RECT 0 24.395 0.070 24.535 ;
    RECT 0 24.605 0.070 24.745 ;
    RECT 0 24.815 0.070 24.955 ;
    RECT 0 25.025 0.070 25.165 ;
    RECT 0 25.235 0.070 25.375 ;
    RECT 0 25.445 0.070 27.265 ;
    RECT 0 27.335 0.070 27.475 ;
    RECT 0 27.545 0.070 27.685 ;
    RECT 0 27.755 0.070 27.895 ;
    RECT 0 27.965 0.070 28.105 ;
    RECT 0 28.175 0.070 29.995 ;
    RECT 0 30.065 0.070 30.205 ;
    RECT 0 30.275 0.070 30.415 ;
    RECT 0 30.485 0.070 33.600 ;
    LAYER metal4 ;
    RECT 0 0 55.100 2.100 ;
    RECT 0 31.500 55.100 33.600 ;
    RECT 0.000 2.100 1.960 31.500 ;
    RECT 2.240 2.100 3.640 31.500 ;
    RECT 3.920 2.100 5.320 31.500 ;
    RECT 5.600 2.100 7.000 31.500 ;
    RECT 7.280 2.100 8.680 31.500 ;
    RECT 8.960 2.100 10.360 31.500 ;
    RECT 10.640 2.100 12.040 31.500 ;
    RECT 12.320 2.100 13.720 31.500 ;
    RECT 14.000 2.100 15.400 31.500 ;
    RECT 15.680 2.100 17.080 31.500 ;
    RECT 17.360 2.100 18.760 31.500 ;
    RECT 19.040 2.100 20.440 31.500 ;
    RECT 20.720 2.100 22.120 31.500 ;
    RECT 22.400 2.100 23.800 31.500 ;
    RECT 24.080 2.100 25.480 31.500 ;
    RECT 25.760 2.100 27.160 31.500 ;
    RECT 27.440 2.100 28.840 31.500 ;
    RECT 29.120 2.100 30.520 31.500 ;
    RECT 30.800 2.100 32.200 31.500 ;
    RECT 32.480 2.100 33.880 31.500 ;
    RECT 34.160 2.100 35.560 31.500 ;
    RECT 35.840 2.100 37.240 31.500 ;
    RECT 37.520 2.100 38.920 31.500 ;
    RECT 39.200 2.100 40.600 31.500 ;
    RECT 40.880 2.100 42.280 31.500 ;
    RECT 42.560 2.100 43.960 31.500 ;
    RECT 44.240 2.100 45.640 31.500 ;
    RECT 45.920 2.100 47.320 31.500 ;
    RECT 47.600 2.100 49.000 31.500 ;
    RECT 49.280 2.100 50.680 31.500 ;
    RECT 50.960 2.100 52.360 31.500 ;
    RECT 52.640 2.100 55.100 31.500 ;
    LAYER OVERLAP ;
    RECT 0 0 55.100 33.600 ;
  END
END fakeram45_32x32

END LIBRARY
