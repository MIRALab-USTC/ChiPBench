VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MACRO macro_9x3
  FOREIGN macro_9x3 0 0 ;
  CLASS BLOCK ;
  SIZE 43.935 BY 169.73 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 166.515 42.75 166.685 ;
        RECT  1.14 163.715 42.75 163.885 ;
        RECT  1.14 160.915 42.75 161.085 ;
        RECT  1.14 158.115 42.75 158.285 ;
        RECT  1.14 155.315 42.75 155.485 ;
        RECT  1.14 152.515 42.75 152.685 ;
        RECT  1.14 149.715 42.75 149.885 ;
        RECT  1.14 146.915 42.75 147.085 ;
        RECT  1.14 144.115 42.75 144.285 ;
        RECT  1.14 141.315 42.75 141.485 ;
        RECT  1.14 138.515 42.75 138.685 ;
        RECT  1.14 135.715 42.75 135.885 ;
        RECT  1.14 132.915 42.75 133.085 ;
        RECT  1.14 130.115 42.75 130.285 ;
        RECT  1.14 127.315 42.75 127.485 ;
        RECT  1.14 124.515 42.75 124.685 ;
        RECT  1.14 121.715 42.75 121.885 ;
        RECT  1.14 118.915 42.75 119.085 ;
        RECT  1.14 116.115 42.75 116.285 ;
        RECT  1.14 113.315 42.75 113.485 ;
        RECT  1.14 110.515 42.75 110.685 ;
        RECT  1.14 107.715 42.75 107.885 ;
        RECT  1.14 104.915 42.75 105.085 ;
        RECT  1.14 102.115 42.75 102.285 ;
        RECT  1.14 99.315 42.75 99.485 ;
        RECT  1.14 96.515 42.75 96.685 ;
        RECT  1.14 93.715 42.75 93.885 ;
        RECT  1.14 90.915 42.75 91.085 ;
        RECT  1.14 88.115 42.75 88.285 ;
        RECT  1.14 85.315 42.75 85.485 ;
        RECT  1.14 82.515 42.75 82.685 ;
        RECT  1.14 79.715 42.75 79.885 ;
        RECT  1.14 76.915 42.75 77.085 ;
        RECT  1.14 74.115 42.75 74.285 ;
        RECT  1.14 71.315 42.75 71.485 ;
        RECT  1.14 68.515 42.75 68.685 ;
        RECT  1.14 65.715 42.75 65.885 ;
        RECT  1.14 62.915 42.75 63.085 ;
        RECT  1.14 60.115 42.75 60.285 ;
        RECT  1.14 57.315 42.75 57.485 ;
        RECT  1.14 54.515 42.75 54.685 ;
        RECT  1.14 51.715 42.75 51.885 ;
        RECT  1.14 48.915 42.75 49.085 ;
        RECT  1.14 46.115 42.75 46.285 ;
        RECT  1.14 43.315 42.75 43.485 ;
        RECT  1.14 40.515 42.75 40.685 ;
        RECT  1.14 37.715 42.75 37.885 ;
        RECT  1.14 34.915 42.75 35.085 ;
        RECT  1.14 32.115 42.75 32.285 ;
        RECT  1.14 29.315 42.75 29.485 ;
        RECT  1.14 26.515 42.75 26.685 ;
        RECT  1.14 23.715 42.75 23.885 ;
        RECT  1.14 20.915 42.75 21.085 ;
        RECT  1.14 18.115 42.75 18.285 ;
        RECT  1.14 15.315 42.75 15.485 ;
        RECT  1.14 12.515 42.75 12.685 ;
        RECT  1.14 9.715 42.75 9.885 ;
        RECT  1.14 6.915 42.75 7.085 ;
        RECT  1.14 4.115 42.75 4.285 ;
        RECT  1.14 1.315 42.75 1.485 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 167.915 42.75 168.085 ;
        RECT  1.14 165.115 42.75 165.285 ;
        RECT  1.14 162.315 42.75 162.485 ;
        RECT  1.14 159.515 42.75 159.685 ;
        RECT  1.14 156.715 42.75 156.885 ;
        RECT  1.14 153.915 42.75 154.085 ;
        RECT  1.14 151.115 42.75 151.285 ;
        RECT  1.14 148.315 42.75 148.485 ;
        RECT  1.14 145.515 42.75 145.685 ;
        RECT  1.14 142.715 42.75 142.885 ;
        RECT  1.14 139.915 42.75 140.085 ;
        RECT  1.14 137.115 42.75 137.285 ;
        RECT  1.14 134.315 42.75 134.485 ;
        RECT  1.14 131.515 42.75 131.685 ;
        RECT  1.14 128.715 42.75 128.885 ;
        RECT  1.14 125.915 42.75 126.085 ;
        RECT  1.14 123.115 42.75 123.285 ;
        RECT  1.14 120.315 42.75 120.485 ;
        RECT  1.14 117.515 42.75 117.685 ;
        RECT  1.14 114.715 42.75 114.885 ;
        RECT  1.14 111.915 42.75 112.085 ;
        RECT  1.14 109.115 42.75 109.285 ;
        RECT  1.14 106.315 42.75 106.485 ;
        RECT  1.14 103.515 42.75 103.685 ;
        RECT  1.14 100.715 42.75 100.885 ;
        RECT  1.14 97.915 42.75 98.085 ;
        RECT  1.14 95.115 42.75 95.285 ;
        RECT  1.14 92.315 42.75 92.485 ;
        RECT  1.14 89.515 42.75 89.685 ;
        RECT  1.14 86.715 42.75 86.885 ;
        RECT  1.14 83.915 42.75 84.085 ;
        RECT  1.14 81.115 42.75 81.285 ;
        RECT  1.14 78.315 42.75 78.485 ;
        RECT  1.14 75.515 42.75 75.685 ;
        RECT  1.14 72.715 42.75 72.885 ;
        RECT  1.14 69.915 42.75 70.085 ;
        RECT  1.14 67.115 42.75 67.285 ;
        RECT  1.14 64.315 42.75 64.485 ;
        RECT  1.14 61.515 42.75 61.685 ;
        RECT  1.14 58.715 42.75 58.885 ;
        RECT  1.14 55.915 42.75 56.085 ;
        RECT  1.14 53.115 42.75 53.285 ;
        RECT  1.14 50.315 42.75 50.485 ;
        RECT  1.14 47.515 42.75 47.685 ;
        RECT  1.14 44.715 42.75 44.885 ;
        RECT  1.14 41.915 42.75 42.085 ;
        RECT  1.14 39.115 42.75 39.285 ;
        RECT  1.14 36.315 42.75 36.485 ;
        RECT  1.14 33.515 42.75 33.685 ;
        RECT  1.14 30.715 42.75 30.885 ;
        RECT  1.14 27.915 42.75 28.085 ;
        RECT  1.14 25.115 42.75 25.285 ;
        RECT  1.14 22.315 42.75 22.485 ;
        RECT  1.14 19.515 42.75 19.685 ;
        RECT  1.14 16.715 42.75 16.885 ;
        RECT  1.14 13.915 42.75 14.085 ;
        RECT  1.14 11.115 42.75 11.285 ;
        RECT  1.14 8.315 42.75 8.485 ;
        RECT  1.14 5.515 42.75 5.685 ;
        RECT  1.14 2.715 42.75 2.885 ;
    END
  END VDD
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.865 84.595 43.935 84.665 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.865 147.595 43.935 147.665 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 148.155 0.07 148.225 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.865 42.315 43.935 42.385 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 84.875 0.07 84.945 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 127.155 0.07 127.225 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  43.145 169.59 43.285 169.73 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.865 63.315 43.935 63.385 ;
    END
  END addr[8]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  42.585 0 42.725 0.14 ;
    END
  END clk
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.875 0.07 21.945 ;
    END
  END cs
  PIN di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.865 126.595 43.935 126.665 ;
    END
  END di[0]
  PIN di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 42.875 0.07 42.945 ;
    END
  END di[1]
  PIN di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  1.145 169.59 1.285 169.73 ;
    END
  END di[2]
  PIN doq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.865 21.315 43.935 21.385 ;
    END
  END doq[0]
  PIN doq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 63.875 0.07 63.945 ;
    END
  END doq[1]
  PIN doq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 106.155 0.07 106.225 ;
    END
  END doq[2]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  43.865 105.595 43.935 105.665 ;
    END
  END we
  OBS
    LAYER metal1 ;
     RECT  0 -0.085 3.23 169.73 ;
     RECT  3.23 0 43.935 169.73 ;
    LAYER metal2 ;
     RECT  0 0 43.935 169.73 ;
    LAYER metal3 ;
     RECT  0 0 43.935 169.73 ;
    LAYER metal4 ;
     RECT  0 0 43.935 169.73 ;
  END
END macro_9x3
END LIBRARY
