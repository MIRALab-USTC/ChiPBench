VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MACRO fifo_v3_1
  FOREIGN fifo_v3_1 0 0 ;
  CLASS BLOCK ;
  SIZE 35.905 BY 42.685 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 40.515 34.77 40.685 ;
        RECT  1.14 37.715 34.77 37.885 ;
        RECT  1.14 34.915 34.77 35.085 ;
        RECT  1.14 32.115 34.77 32.285 ;
        RECT  1.14 29.315 34.77 29.485 ;
        RECT  1.14 26.515 34.77 26.685 ;
        RECT  1.14 23.715 34.77 23.885 ;
        RECT  1.14 20.915 34.77 21.085 ;
        RECT  1.14 18.115 34.77 18.285 ;
        RECT  1.14 15.315 34.77 15.485 ;
        RECT  1.14 12.515 34.77 12.685 ;
        RECT  1.14 9.715 34.77 9.885 ;
        RECT  1.14 6.915 34.77 7.085 ;
        RECT  1.14 4.115 34.77 4.285 ;
        RECT  1.14 1.315 34.77 1.485 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal4 ;
        RECT  1.14 39.115 34.77 39.285 ;
        RECT  1.14 36.315 34.77 36.485 ;
        RECT  1.14 33.515 34.77 33.685 ;
        RECT  1.14 30.715 34.77 30.885 ;
        RECT  1.14 27.915 34.77 28.085 ;
        RECT  1.14 25.115 34.77 25.285 ;
        RECT  1.14 22.315 34.77 22.485 ;
        RECT  1.14 19.515 34.77 19.685 ;
        RECT  1.14 16.715 34.77 16.885 ;
        RECT  1.14 13.915 34.77 14.085 ;
        RECT  1.14 11.115 34.77 11.285 ;
        RECT  1.14 8.315 34.77 8.485 ;
        RECT  1.14 5.515 34.77 5.685 ;
        RECT  1.14 2.715 34.77 2.885 ;
    END
  END VDD
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  5.065 42.545 5.205 42.685 ;
    END
  END clk_i
  PIN data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 35.035 0.07 35.105 ;
    END
  END data_i[0]
  PIN data_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 21.315 35.905 21.385 ;
    END
  END data_i[100]
  PIN data_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 42.545 0.725 42.685 ;
    END
  END data_i[101]
  PIN data_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 6.475 35.905 6.545 ;
    END
  END data_i[102]
  PIN data_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 15.995 35.905 16.065 ;
    END
  END data_i[103]
  PIN data_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 8.715 35.905 8.785 ;
    END
  END data_i[104]
  PIN data_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 28.875 35.905 28.945 ;
    END
  END data_i[105]
  PIN data_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  33.065 42.545 33.205 42.685 ;
    END
  END data_i[106]
  PIN data_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.315 0.07 21.385 ;
    END
  END data_i[107]
  PIN data_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 10.395 35.905 10.465 ;
    END
  END data_i[108]
  PIN data_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 5.355 35.905 5.425 ;
    END
  END data_i[109]
  PIN data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 26.635 0.07 26.705 ;
    END
  END data_i[10]
  PIN data_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 2.555 0.07 2.625 ;
    END
  END data_i[110]
  PIN data_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 30.275 0.07 30.345 ;
    END
  END data_i[111]
  PIN data_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.945 42.545 18.085 42.685 ;
    END
  END data_i[112]
  PIN data_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 29.715 35.905 29.785 ;
    END
  END data_i[113]
  PIN data_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  22.985 0 23.125 0.14 ;
    END
  END data_i[114]
  PIN data_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 34.195 35.905 34.265 ;
    END
  END data_i[115]
  PIN data_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  25.785 0 25.925 0.14 ;
    END
  END data_i[116]
  PIN data_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 37.835 35.905 37.905 ;
    END
  END data_i[117]
  PIN data_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.105 42.545 10.245 42.685 ;
    END
  END data_i[118]
  PIN data_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 32.515 0.07 32.585 ;
    END
  END data_i[119]
  PIN data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 40.075 0.07 40.145 ;
    END
  END data_i[11]
  PIN data_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 15.155 0.07 15.225 ;
    END
  END data_i[120]
  PIN data_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 39.235 35.905 39.305 ;
    END
  END data_i[121]
  PIN data_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 17.675 0.07 17.745 ;
    END
  END data_i[122]
  PIN data_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  15.705 0 15.845 0.14 ;
    END
  END data_i[123]
  PIN data_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 36.715 0.07 36.785 ;
    END
  END data_i[124]
  PIN data_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 19.635 35.905 19.705 ;
    END
  END data_i[125]
  PIN data_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 23.555 0.07 23.625 ;
    END
  END data_i[126]
  PIN data_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 31.955 35.905 32.025 ;
    END
  END data_i[127]
  PIN data_i[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 30.275 35.905 30.345 ;
    END
  END data_i[128]
  PIN data_i[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 24.395 35.905 24.465 ;
    END
  END data_i[129]
  PIN data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 17.115 0.07 17.185 ;
    END
  END data_i[12]
  PIN data_i[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 41.755 35.905 41.825 ;
    END
  END data_i[130]
  PIN data_i[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  24.665 0 24.805 0.14 ;
    END
  END data_i[131]
  PIN data_i[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 1.155 0.07 1.225 ;
    END
  END data_i[132]
  PIN data_i[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 10.395 0.07 10.465 ;
    END
  END data_i[133]
  PIN data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 14.315 35.905 14.385 ;
    END
  END data_i[13]
  PIN data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 36.155 0.07 36.225 ;
    END
  END data_i[14]
  PIN data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.585 0 14.725 0.14 ;
    END
  END data_i[15]
  PIN data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.905 42.545 13.045 42.685 ;
    END
  END data_i[16]
  PIN data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 18.515 0.07 18.585 ;
    END
  END data_i[17]
  PIN data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  23.545 42.545 23.685 42.685 ;
    END
  END data_i[18]
  PIN data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  21.305 42.545 21.445 42.685 ;
    END
  END data_i[19]
  PIN data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.945 42.545 32.085 42.685 ;
    END
  END data_i[1]
  PIN data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  2.265 42.545 2.405 42.685 ;
    END
  END data_i[20]
  PIN data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  6.745 42.545 6.885 42.685 ;
    END
  END data_i[21]
  PIN data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  13.465 42.545 13.605 42.685 ;
    END
  END data_i[22]
  PIN data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  3.945 42.545 4.085 42.685 ;
    END
  END data_i[23]
  PIN data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 18.795 0.07 18.865 ;
    END
  END data_i[24]
  PIN data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 3.955 35.905 4.025 ;
    END
  END data_i[25]
  PIN data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 39.235 0.07 39.305 ;
    END
  END data_i[26]
  PIN data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 35.315 0.07 35.385 ;
    END
  END data_i[27]
  PIN data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  32.505 0 32.645 0.14 ;
    END
  END data_i[28]
  PIN data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 15.435 0.07 15.505 ;
    END
  END data_i[29]
  PIN data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 10.115 35.905 10.185 ;
    END
  END data_i[2]
  PIN data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  3.945 0 4.085 0.14 ;
    END
  END data_i[30]
  PIN data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 36.155 35.905 36.225 ;
    END
  END data_i[31]
  PIN data_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 33.355 35.905 33.425 ;
    END
  END data_i[32]
  PIN data_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.665 0 10.805 0.14 ;
    END
  END data_i[33]
  PIN data_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 37.835 0.07 37.905 ;
    END
  END data_i[34]
  PIN data_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 24.955 0.07 25.025 ;
    END
  END data_i[35]
  PIN data_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 40.075 35.905 40.145 ;
    END
  END data_i[36]
  PIN data_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  8.985 42.545 9.125 42.685 ;
    END
  END data_i[37]
  PIN data_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.025 0 14.165 0.14 ;
    END
  END data_i[38]
  PIN data_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 17.675 35.905 17.745 ;
    END
  END data_i[39]
  PIN data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.675 0.07 31.745 ;
    END
  END data_i[3]
  PIN data_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 38.395 0.07 38.465 ;
    END
  END data_i[40]
  PIN data_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 27.475 0.07 27.545 ;
    END
  END data_i[41]
  PIN data_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 29.435 35.905 29.505 ;
    END
  END data_i[42]
  PIN data_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 34.195 0.07 34.265 ;
    END
  END data_i[43]
  PIN data_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 40.915 0.07 40.985 ;
    END
  END data_i[44]
  PIN data_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 3.115 35.905 3.185 ;
    END
  END data_i[45]
  PIN data_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 20.475 35.905 20.545 ;
    END
  END data_i[46]
  PIN data_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 17.115 35.905 17.185 ;
    END
  END data_i[47]
  PIN data_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 6.195 0.07 6.265 ;
    END
  END data_i[48]
  PIN data_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.305 0 7.445 0.14 ;
    END
  END data_i[49]
  PIN data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 17.955 35.905 18.025 ;
    END
  END data_i[4]
  PIN data_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 20.195 0.07 20.265 ;
    END
  END data_i[50]
  PIN data_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 30.835 0.07 30.905 ;
    END
  END data_i[51]
  PIN data_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  29.705 0 29.845 0.14 ;
    END
  END data_i[52]
  PIN data_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 8.435 35.905 8.505 ;
    END
  END data_i[53]
  PIN data_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 22.995 0.07 23.065 ;
    END
  END data_i[54]
  PIN data_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.955 0.07 32.025 ;
    END
  END data_i[55]
  PIN data_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.385 42.545 31.525 42.685 ;
    END
  END data_i[56]
  PIN data_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  19.065 0 19.205 0.14 ;
    END
  END data_i[57]
  PIN data_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 19.635 0.07 19.705 ;
    END
  END data_i[58]
  PIN data_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.945 0 18.085 0.14 ;
    END
  END data_i[59]
  PIN data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 6.755 0.07 6.825 ;
    END
  END data_i[5]
  PIN data_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 11.235 35.905 11.305 ;
    END
  END data_i[60]
  PIN data_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 40.915 35.905 40.985 ;
    END
  END data_i[61]
  PIN data_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 26.915 0.07 26.985 ;
    END
  END data_i[62]
  PIN data_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  3.385 42.545 3.525 42.685 ;
    END
  END data_i[63]
  PIN data_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  14.585 42.545 14.725 42.685 ;
    END
  END data_i[64]
  PIN data_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  9.545 0 9.685 0.14 ;
    END
  END data_i[65]
  PIN data_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 30.835 35.905 30.905 ;
    END
  END data_i[66]
  PIN data_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 29.995 0.07 30.065 ;
    END
  END data_i[67]
  PIN data_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 7.035 35.905 7.105 ;
    END
  END data_i[68]
  PIN data_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  28.025 42.545 28.165 42.685 ;
    END
  END data_i[69]
  PIN data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  24.105 0 24.245 0.14 ;
    END
  END data_i[6]
  PIN data_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 10.955 35.905 11.025 ;
    END
  END data_i[70]
  PIN data_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.875 0.07 7.945 ;
    END
  END data_i[71]
  PIN data_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 15.435 35.905 15.505 ;
    END
  END data_i[72]
  PIN data_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 12.915 35.905 12.985 ;
    END
  END data_i[73]
  PIN data_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 26.075 0.07 26.145 ;
    END
  END data_i[74]
  PIN data_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 13.755 35.905 13.825 ;
    END
  END data_i[75]
  PIN data_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 22.155 0.07 22.225 ;
    END
  END data_i[76]
  PIN data_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 11.795 0.07 11.865 ;
    END
  END data_i[77]
  PIN data_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  16.825 42.545 16.965 42.685 ;
    END
  END data_i[78]
  PIN data_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 39.515 0.07 39.585 ;
    END
  END data_i[79]
  PIN data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 41.195 0.07 41.265 ;
    END
  END data_i[7]
  PIN data_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  18.505 42.545 18.645 42.685 ;
    END
  END data_i[80]
  PIN data_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 13.475 35.905 13.545 ;
    END
  END data_i[81]
  PIN data_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 41.755 0.07 41.825 ;
    END
  END data_i[82]
  PIN data_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 25.515 35.905 25.585 ;
    END
  END data_i[83]
  PIN data_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 28.595 35.905 28.665 ;
    END
  END data_i[84]
  PIN data_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 3.395 0.07 3.465 ;
    END
  END data_i[85]
  PIN data_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 37.555 0.07 37.625 ;
    END
  END data_i[86]
  PIN data_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 1.435 35.905 1.505 ;
    END
  END data_i[87]
  PIN data_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 31.115 35.905 31.185 ;
    END
  END data_i[88]
  PIN data_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.865 0 8.005 0.14 ;
    END
  END data_i[89]
  PIN data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 15.155 35.905 15.225 ;
    END
  END data_i[8]
  PIN data_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 35.875 0.07 35.945 ;
    END
  END data_i[90]
  PIN data_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 25.235 35.905 25.305 ;
    END
  END data_i[91]
  PIN data_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 22.155 35.905 22.225 ;
    END
  END data_i[92]
  PIN data_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 37.555 35.905 37.625 ;
    END
  END data_i[93]
  PIN data_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 21.875 35.905 21.945 ;
    END
  END data_i[94]
  PIN data_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  21.305 0 21.445 0.14 ;
    END
  END data_i[95]
  PIN data_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 28.035 35.905 28.105 ;
    END
  END data_i[96]
  PIN data_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 15.995 0.07 16.065 ;
    END
  END data_i[97]
  PIN data_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.635 0.07 12.705 ;
    END
  END data_i[98]
  PIN data_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  33.065 0 33.205 0.14 ;
    END
  END data_i[99]
  PIN data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 5.915 0.07 5.985 ;
    END
  END data_i[9]
  PIN data_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  25.225 42.545 25.365 42.685 ;
    END
  END data_o[0]
  PIN data_o[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 27.755 35.905 27.825 ;
    END
  END data_o[100]
  PIN data_o[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 7.875 35.905 7.945 ;
    END
  END data_o[101]
  PIN data_o[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 11.235 0.07 11.305 ;
    END
  END data_o[102]
  PIN data_o[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 28.595 0.07 28.665 ;
    END
  END data_o[103]
  PIN data_o[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 24.395 0.07 24.465 ;
    END
  END data_o[104]
  PIN data_o[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  19.625 0 19.765 0.14 ;
    END
  END data_o[105]
  PIN data_o[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 23.835 0.07 23.905 ;
    END
  END data_o[106]
  PIN data_o[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  21.865 42.545 22.005 42.685 ;
    END
  END data_o[107]
  PIN data_o[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.035 0.07 7.105 ;
    END
  END data_o[108]
  PIN data_o[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.185 0 34.325 0.14 ;
    END
  END data_o[109]
  PIN data_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 31.115 0.07 31.185 ;
    END
  END data_o[10]
  PIN data_o[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 14.315 0.07 14.385 ;
    END
  END data_o[110]
  PIN data_o[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 5.355 0.07 5.425 ;
    END
  END data_o[111]
  PIN data_o[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  30.265 42.545 30.405 42.685 ;
    END
  END data_o[112]
  PIN data_o[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.035 0.07 21.105 ;
    END
  END data_o[113]
  PIN data_o[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 21.035 35.905 21.105 ;
    END
  END data_o[114]
  PIN data_o[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 36.715 35.905 36.785 ;
    END
  END data_o[115]
  PIN data_o[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 18.515 35.905 18.585 ;
    END
  END data_o[116]
  PIN data_o[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 1.155 35.905 1.225 ;
    END
  END data_o[117]
  PIN data_o[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 32.515 35.905 32.585 ;
    END
  END data_o[118]
  PIN data_o[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 9.275 35.905 9.345 ;
    END
  END data_o[119]
  PIN data_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 39.515 35.905 39.585 ;
    END
  END data_o[11]
  PIN data_o[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 4.795 35.905 4.865 ;
    END
  END data_o[120]
  PIN data_o[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  11.785 42.545 11.925 42.685 ;
    END
  END data_o[121]
  PIN data_o[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  6.185 0 6.325 0.14 ;
    END
  END data_o[122]
  PIN data_o[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 20.475 0.07 20.545 ;
    END
  END data_o[123]
  PIN data_o[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  26.345 0 26.485 0.14 ;
    END
  END data_o[124]
  PIN data_o[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 22.715 35.905 22.785 ;
    END
  END data_o[125]
  PIN data_o[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 10.115 0.07 10.185 ;
    END
  END data_o[126]
  PIN data_o[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 6.195 35.905 6.265 ;
    END
  END data_o[127]
  PIN data_o[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  8.425 42.545 8.565 42.685 ;
    END
  END data_o[128]
  PIN data_o[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 35.035 35.905 35.105 ;
    END
  END data_o[129]
  PIN data_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 26.075 35.905 26.145 ;
    END
  END data_o[12]
  PIN data_o[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  19.625 42.545 19.765 42.685 ;
    END
  END data_o[130]
  PIN data_o[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  22.985 42.545 23.125 42.685 ;
    END
  END data_o[131]
  PIN data_o[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 11.795 35.905 11.865 ;
    END
  END data_o[132]
  PIN data_o[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 3.675 0.07 3.745 ;
    END
  END data_o[133]
  PIN data_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 10.955 0.07 11.025 ;
    END
  END data_o[13]
  PIN data_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 29.435 0.07 29.505 ;
    END
  END data_o[14]
  PIN data_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  26.905 42.545 27.045 42.685 ;
    END
  END data_o[15]
  PIN data_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  7.305 42.545 7.445 42.685 ;
    END
  END data_o[16]
  PIN data_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 16.835 0.07 16.905 ;
    END
  END data_o[17]
  PIN data_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 36.995 0.07 37.065 ;
    END
  END data_o[18]
  PIN data_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 1.715 0.07 1.785 ;
    END
  END data_o[19]
  PIN data_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 24.675 35.905 24.745 ;
    END
  END data_o[1]
  PIN data_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 8.435 0.07 8.505 ;
    END
  END data_o[20]
  PIN data_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 23.555 35.905 23.625 ;
    END
  END data_o[21]
  PIN data_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 16.275 35.905 16.345 ;
    END
  END data_o[22]
  PIN data_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 7.595 35.905 7.665 ;
    END
  END data_o[23]
  PIN data_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  33.625 42.545 33.765 42.685 ;
    END
  END data_o[24]
  PIN data_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 35.315 35.905 35.385 ;
    END
  END data_o[25]
  PIN data_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  29.145 0 29.285 0.14 ;
    END
  END data_o[26]
  PIN data_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 2.835 0.07 2.905 ;
    END
  END data_o[27]
  PIN data_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 14.595 0.07 14.665 ;
    END
  END data_o[28]
  PIN data_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  5.625 42.545 5.765 42.685 ;
    END
  END data_o[29]
  PIN data_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  28.025 0 28.165 0.14 ;
    END
  END data_o[2]
  PIN data_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  5.625 0 5.765 0.14 ;
    END
  END data_o[30]
  PIN data_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 4.235 0.07 4.305 ;
    END
  END data_o[31]
  PIN data_o[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 27.755 0.07 27.825 ;
    END
  END data_o[32]
  PIN data_o[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 5.075 0.07 5.145 ;
    END
  END data_o[33]
  PIN data_o[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  20.745 0 20.885 0.14 ;
    END
  END data_o[34]
  PIN data_o[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 40.355 35.905 40.425 ;
    END
  END data_o[35]
  PIN data_o[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 1.995 0.07 2.065 ;
    END
  END data_o[36]
  PIN data_o[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 3.675 35.905 3.745 ;
    END
  END data_o[37]
  PIN data_o[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 41.195 35.905 41.265 ;
    END
  END data_o[38]
  PIN data_o[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 2.835 35.905 2.905 ;
    END
  END data_o[39]
  PIN data_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  16.265 0 16.405 0.14 ;
    END
  END data_o[3]
  PIN data_o[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  2.825 0 2.965 0.14 ;
    END
  END data_o[40]
  PIN data_o[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 9.555 35.905 9.625 ;
    END
  END data_o[41]
  PIN data_o[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 16.835 35.905 16.905 ;
    END
  END data_o[42]
  PIN data_o[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 9.275 0.07 9.345 ;
    END
  END data_o[43]
  PIN data_o[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 32.795 35.905 32.865 ;
    END
  END data_o[44]
  PIN data_o[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 32.795 0.07 32.865 ;
    END
  END data_o[45]
  PIN data_o[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 34.475 0.07 34.545 ;
    END
  END data_o[46]
  PIN data_o[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 33.355 0.07 33.425 ;
    END
  END data_o[47]
  PIN data_o[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  2.265 0 2.405 0.14 ;
    END
  END data_o[48]
  PIN data_o[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  11.225 0 11.365 0.14 ;
    END
  END data_o[49]
  PIN data_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 23.835 35.905 23.905 ;
    END
  END data_o[4]
  PIN data_o[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  30.825 0 30.965 0.14 ;
    END
  END data_o[50]
  PIN data_o[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  28.585 42.545 28.725 42.685 ;
    END
  END data_o[51]
  PIN data_o[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 38.675 35.905 38.745 ;
    END
  END data_o[52]
  PIN data_o[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 38.675 0.07 38.745 ;
    END
  END data_o[53]
  PIN data_o[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 19.355 0.07 19.425 ;
    END
  END data_o[54]
  PIN data_o[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 26.355 35.905 26.425 ;
    END
  END data_o[55]
  PIN data_o[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 38.395 35.905 38.465 ;
    END
  END data_o[56]
  PIN data_o[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 25.795 0.07 25.865 ;
    END
  END data_o[57]
  PIN data_o[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 31.675 35.905 31.745 ;
    END
  END data_o[58]
  PIN data_o[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 19.355 35.905 19.425 ;
    END
  END data_o[59]
  PIN data_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 1.995 35.905 2.065 ;
    END
  END data_o[5]
  PIN data_o[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.745 42.545 34.885 42.685 ;
    END
  END data_o[60]
  PIN data_o[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  1.705 42.545 1.845 42.685 ;
    END
  END data_o[61]
  PIN data_o[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  17.385 0 17.525 0.14 ;
    END
  END data_o[62]
  PIN data_o[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 16.275 0.07 16.345 ;
    END
  END data_o[63]
  PIN data_o[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.075 0.07 12.145 ;
    END
  END data_o[64]
  PIN data_o[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 18.795 35.905 18.865 ;
    END
  END data_o[65]
  PIN data_o[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 22.715 0.07 22.785 ;
    END
  END data_o[66]
  PIN data_o[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 12.075 35.905 12.145 ;
    END
  END data_o[67]
  PIN data_o[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  8.985 0 9.125 0.14 ;
    END
  END data_o[68]
  PIN data_o[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  27.465 0 27.605 0.14 ;
    END
  END data_o[69]
  PIN data_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 22.995 35.905 23.065 ;
    END
  END data_o[6]
  PIN data_o[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  29.705 42.545 29.845 42.685 ;
    END
  END data_o[70]
  PIN data_o[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 35.875 35.905 35.945 ;
    END
  END data_o[71]
  PIN data_o[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 12.635 35.905 12.705 ;
    END
  END data_o[72]
  PIN data_o[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 9.555 0.07 9.625 ;
    END
  END data_o[73]
  PIN data_o[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 27.195 35.905 27.265 ;
    END
  END data_o[74]
  PIN data_o[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  1.145 0 1.285 0.14 ;
    END
  END data_o[75]
  PIN data_o[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 36.995 35.905 37.065 ;
    END
  END data_o[76]
  PIN data_o[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  26.345 42.545 26.485 42.685 ;
    END
  END data_o[77]
  PIN data_o[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 14.595 35.905 14.665 ;
    END
  END data_o[78]
  PIN data_o[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  24.665 42.545 24.805 42.685 ;
    END
  END data_o[79]
  PIN data_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 12.915 0.07 12.985 ;
    END
  END data_o[7]
  PIN data_o[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 13.755 0.07 13.825 ;
    END
  END data_o[80]
  PIN data_o[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 2.275 35.905 2.345 ;
    END
  END data_o[81]
  PIN data_o[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END data_o[82]
  PIN data_o[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 5.635 35.905 5.705 ;
    END
  END data_o[83]
  PIN data_o[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 17.955 0.07 18.025 ;
    END
  END data_o[84]
  PIN data_o[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 29.155 0.07 29.225 ;
    END
  END data_o[85]
  PIN data_o[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 8.715 0.07 8.785 ;
    END
  END data_o[86]
  PIN data_o[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 13.475 0.07 13.545 ;
    END
  END data_o[87]
  PIN data_o[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.345 0 12.485 0.14 ;
    END
  END data_o[88]
  PIN data_o[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  4.505 0 4.645 0.14 ;
    END
  END data_o[89]
  PIN data_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  10.665 42.545 10.805 42.685 ;
    END
  END data_o[8]
  PIN data_o[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 40.355 0.07 40.425 ;
    END
  END data_o[90]
  PIN data_o[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  31.385 0 31.525 0.14 ;
    END
  END data_o[91]
  PIN data_o[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  20.185 42.545 20.325 42.685 ;
    END
  END data_o[92]
  PIN data_o[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 20.195 35.905 20.265 ;
    END
  END data_o[93]
  PIN data_o[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 21.875 0.07 21.945 ;
    END
  END data_o[94]
  PIN data_o[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 34.475 35.905 34.545 ;
    END
  END data_o[95]
  PIN data_o[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  12.905 0 13.045 0.14 ;
    END
  END data_o[96]
  PIN data_o[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  22.425 0 22.565 0.14 ;
    END
  END data_o[97]
  PIN data_o[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 4.515 0.07 4.585 ;
    END
  END data_o[98]
  PIN data_o[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 33.635 35.905 33.705 ;
    END
  END data_o[99]
  PIN data_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  34.745 0 34.885 0.14 ;
    END
  END data_o[9]
  PIN empty_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  16.265 42.545 16.405 42.685 ;
    END
  END empty_o
  PIN flush_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT  15.145 42.545 15.285 42.685 ;
    END
  END flush_i
  PIN full_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 28.315 0.07 28.385 ;
    END
  END full_o
  PIN pop_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 33.635 0.07 33.705 ;
    END
  END pop_i
  PIN push_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 4.515 35.905 4.585 ;
    END
  END push_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 7.595 0.07 7.665 ;
    END
  END rst_ni
  PIN testmode_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  0 25.235 0.07 25.305 ;
    END
  END testmode_i
  PIN usage_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT  35.835 26.915 35.905 26.985 ;
    END
  END usage_o
  OBS
    LAYER metal1 ;
     RECT  0 -0.085 3.8 42.685 ;
     RECT  3.8 0 35.905 42.685 ;
    LAYER metal2 ;
     RECT  0 0 35.905 42.685 ;
    LAYER metal3 ;
     RECT  0 0 35.905 42.685 ;
    LAYER metal4 ;
     RECT  0 0 35.905 42.685 ;
  END
END fifo_v3_1
END LIBRARY
